
# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0
#
# Autogenerated by https://www.asicsforthemasses.com
#

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;


MACRO sky130_fd_io__corner_bus_overlay
  CLASS PAD ;
  ORIGIN  0.000000  0.000000 ;
  FOREIGN sky130_fd_io__corner_bus_overlay  0.000000  0.000000 ;
  SIZE 200 BY  203.6650 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT  0.000000 56.790000  0.500000 59.770000 ;
        RECT 53.125000  0.000000 56.105000  0.500000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT  0.000000 52.030000  0.575000 55.010000 ;
        RECT 48.365000  0.000000 51.345000  0.575000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.550000 1.270000 17.200000 ;
      LAYER met4 ;
        RECT 8.885000 0.000000 13.535000 1.270000 ;
      LAYER met5 ;
        RECT 0.000000 12.650000 1.270000 17.100000 ;
      LAYER met5 ;
        RECT 8.985000 0.000000 13.435000 1.270000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 5.700000 1.270000 11.150000 ;
      LAYER met4 ;
        RECT 2.035000 0.000000 7.485000 1.270000 ;
      LAYER met5 ;
        RECT 0.000000 5.800000 1.270000 11.050000 ;
      LAYER met5 ;
        RECT 2.135000 0.000000 7.385000 1.270000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 18.600000 1.255000 22.050000 ;
      LAYER met4 ;
        RECT 14.935000 0.000000 18.385000 1.255000 ;
      LAYER met5 ;
        RECT 0.000000 18.700000 1.255000 21.950000 ;
      LAYER met5 ;
        RECT 15.035000 0.000000 18.285000 1.255000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 23.450000 1.270000 28.100000 ;
      LAYER met4 ;
        RECT 0.000000 73.705000 1.270000 98.665000 ;
      LAYER met4 ;
        RECT 19.785000 0.000000 24.435000 1.270000 ;
        RECT 70.040000 0.000000 95.000000 1.270000 ;
      LAYER met5 ;
        RECT 0.000000 23.550000 1.270000 28.000000 ;
        RECT 0.000000 73.700000 1.270000 98.650000 ;
      LAYER met5 ;
        RECT 19.885000 0.000000 24.335000 1.270000 ;
        RECT 70.035000 0.000000 94.985000 1.270000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 67.750000 1.270000 72.200000 ;
      LAYER met4 ;
        RECT 64.085000 0.000000 68.535000 1.270000 ;
      LAYER met5 ;
        RECT  0.000000 67.850000  1.270000 72.100000 ;
        RECT 64.185000  0.000000 68.435000  1.270000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 40.400000 1.270000 43.850000 ;
      LAYER met4 ;
        RECT 0.000000 51.400000 1.270000 51.730000 ;
        RECT 0.000000 55.310000 1.270000 56.490000 ;
        RECT 0.000000 60.070000 1.270000 60.400000 ;
      LAYER met4 ;
        RECT 36.735000 0.000000 40.185000 1.270000 ;
        RECT 47.735000 0.000000 48.065000 1.270000 ;
        RECT 51.645000 0.000000 52.825000 1.270000 ;
        RECT 56.405000 0.000000 56.735000 1.270000 ;
      LAYER met5 ;
        RECT 0.000000 40.505000 1.270000 43.750000 ;
      LAYER met5 ;
        RECT 0.000000 51.400000 1.270000 60.400000 ;
      LAYER met5 ;
        RECT 36.840000 0.000000 40.085000 1.270000 ;
        RECT 47.735000 0.000000 56.735000 1.270000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 45.250000 1.270000 49.900000 ;
      LAYER met4 ;
        RECT 41.585000 0.000000 46.235000 1.270000 ;
      LAYER met5 ;
        RECT  0.000000 45.350000  1.270000 49.800000 ;
        RECT 41.685000  0.000000 46.135000  1.270000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT  25.835000 0.000000  30.485000 1.270000 ;
        RECT 175.785000 0.000000 200.000000 1.270000 ;
      LAYER met4 ;
        RECT 0.000000 179.450000 1.270000 203.665000 ;
      LAYER met4 ;
        RECT 0.000000 29.500000 1.270000 34.150000 ;
      LAYER met5 ;
        RECT  25.935000 0.000000  30.385000 1.270000 ;
        RECT 175.785000 0.000000 200.000000 1.270000 ;
      LAYER met5 ;
        RECT 0.000000  29.600000 1.270000  34.050000 ;
        RECT 0.000000 179.450000 1.270000 203.665000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 61.900000 1.270000 66.350000 ;
      LAYER met4 ;
        RECT 58.235000 0.000000 62.685000 1.270000 ;
      LAYER met5 ;
        RECT  0.000000 62.000000  1.270000 66.250000 ;
        RECT 58.335000  0.000000 62.585000  1.270000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 35.550000 1.270000 39.000000 ;
      LAYER met4 ;
        RECT 31.885000 0.000000 35.335000 1.270000 ;
      LAYER met5 ;
        RECT 0.000000 35.650000 1.270000 38.900000 ;
      LAYER met5 ;
        RECT 31.985000 0.000000 35.235000 1.270000 ;
    END
  END VSWITCH
END sky130_fd_io__corner_bus_overlay


MACRO sky130_fd_io__top_ground_lvc_wpad
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN G_PAD
    ANTENNAPARTIALMETALSIDEAREA  243.2170 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 31.695000 162.765000 52.340000 167.120000 ;
    END
  END G_PAD
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 17.630000 5.115000 53.535000 9.540000 ;
        RECT 17.635000 5.110000 53.535000 5.115000 ;
        RECT 17.705000 5.040000 53.535000 5.110000 ;
        RECT 17.775000 4.970000 53.535000 5.040000 ;
        RECT 17.845000 4.900000 53.535000 4.970000 ;
        RECT 17.915000 4.830000 53.535000 4.900000 ;
        RECT 17.985000 4.760000 53.535000 4.830000 ;
        RECT 18.055000 4.690000 53.535000 4.760000 ;
        RECT 18.125000 4.620000 53.535000 4.690000 ;
        RECT 18.195000 4.550000 53.535000 4.620000 ;
        RECT 18.265000 4.480000 53.535000 4.550000 ;
        RECT 18.335000 4.410000 53.535000 4.480000 ;
        RECT 18.405000 4.340000 53.535000 4.410000 ;
        RECT 18.475000 4.270000 53.535000 4.340000 ;
        RECT 18.545000 4.200000 53.535000 4.270000 ;
        RECT 18.615000 4.130000 53.535000 4.200000 ;
        RECT 18.685000 4.060000 53.535000 4.130000 ;
        RECT 18.755000 3.990000 53.535000 4.060000 ;
        RECT 18.825000 3.920000 53.535000 3.990000 ;
        RECT 18.895000 3.850000 53.535000 3.920000 ;
        RECT 18.965000 3.780000 53.535000 3.850000 ;
        RECT 19.035000 3.710000 53.535000 3.780000 ;
        RECT 19.105000 3.640000 53.535000 3.710000 ;
        RECT 19.175000 3.570000 53.535000 3.640000 ;
        RECT 19.245000 3.500000 53.535000 3.570000 ;
        RECT 19.315000 3.430000 53.535000 3.500000 ;
        RECT 19.385000 3.360000 53.535000 3.430000 ;
        RECT 19.455000 3.290000 53.535000 3.360000 ;
        RECT 19.525000 3.220000 53.535000 3.290000 ;
        RECT 19.595000 3.150000 53.535000 3.220000 ;
        RECT 19.665000 3.080000 53.535000 3.150000 ;
        RECT 19.735000 3.010000 53.535000 3.080000 ;
        RECT 19.805000 2.940000 53.535000 3.010000 ;
        RECT 19.875000 2.870000 53.535000 2.940000 ;
        RECT 19.945000 2.800000 53.535000 2.870000 ;
        RECT 20.015000 2.730000 53.535000 2.800000 ;
        RECT 20.085000 2.660000 53.535000 2.730000 ;
        RECT 20.155000 2.590000 53.535000 2.660000 ;
        RECT 20.225000 2.520000 53.535000 2.590000 ;
        RECT 20.295000 2.450000 53.535000 2.520000 ;
        RECT 20.365000 2.380000 53.535000 2.450000 ;
        RECT 20.435000 2.310000 53.535000 2.380000 ;
        RECT 20.505000 2.240000 53.535000 2.310000 ;
        RECT 20.575000 2.170000 53.535000 2.240000 ;
        RECT 20.645000 2.100000 53.535000 2.170000 ;
        RECT 20.715000 2.030000 53.535000 2.100000 ;
        RECT 20.785000 1.960000 53.535000 2.030000 ;
        RECT 20.855000 1.890000 53.535000 1.960000 ;
        RECT 20.925000 0.000000 53.535000 1.820000 ;
        RECT 20.925000 1.820000 53.535000 1.890000 ;
    END
  END BDY2_B2B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 15.605000  94.310000 23.935000  94.460000 ;
        RECT 15.605000  94.460000 23.785000  94.610000 ;
        RECT 15.605000  94.610000 23.635000  94.760000 ;
        RECT 15.605000  94.760000 23.485000  94.910000 ;
        RECT 15.605000  94.910000 23.335000  95.060000 ;
        RECT 15.605000  95.060000 23.185000  95.210000 ;
        RECT 15.605000  95.210000 23.035000  95.360000 ;
        RECT 15.605000  95.360000 22.885000  95.510000 ;
        RECT 15.605000  95.510000 22.735000  95.660000 ;
        RECT 15.605000  95.660000 22.585000  95.810000 ;
        RECT 15.605000  95.810000 22.435000  95.960000 ;
        RECT 15.605000  95.960000 22.285000  96.110000 ;
        RECT 15.605000  96.110000 22.135000  96.260000 ;
        RECT 15.605000  96.260000 21.985000  96.410000 ;
        RECT 15.605000  96.410000 21.835000  96.560000 ;
        RECT 15.605000  96.560000 21.685000  96.710000 ;
        RECT 15.605000  96.710000 21.605000  96.790000 ;
        RECT 15.605000  96.790000 21.605000 167.100000 ;
        RECT 15.605000 167.100000 21.605000 167.250000 ;
        RECT 15.605000 167.250000 21.755000 167.400000 ;
        RECT 15.605000 167.400000 21.905000 167.550000 ;
        RECT 15.605000 167.550000 22.055000 167.700000 ;
        RECT 15.605000 167.700000 22.205000 167.850000 ;
        RECT 15.605000 167.850000 22.355000 168.000000 ;
        RECT 15.605000 168.000000 22.505000 168.150000 ;
        RECT 15.605000 168.150000 22.655000 168.300000 ;
        RECT 15.605000 168.300000 22.805000 168.450000 ;
        RECT 15.605000 168.450000 22.955000 168.600000 ;
        RECT 15.605000 168.600000 23.105000 168.750000 ;
        RECT 15.605000 168.750000 23.255000 168.900000 ;
        RECT 15.605000 168.900000 23.405000 169.050000 ;
        RECT 15.605000 169.050000 23.555000 169.200000 ;
        RECT 15.605000 169.200000 23.705000 169.350000 ;
        RECT 15.605000 169.350000 23.855000 169.500000 ;
        RECT 15.605000 169.500000 24.005000 169.650000 ;
        RECT 15.605000 169.650000 24.155000 169.800000 ;
        RECT 15.605000 169.800000 24.305000 169.950000 ;
        RECT 15.605000 169.950000 24.455000 170.100000 ;
        RECT 15.605000 170.100000 24.605000 170.250000 ;
        RECT 15.605000 170.250000 24.755000 170.400000 ;
        RECT 15.605000 170.400000 24.905000 170.550000 ;
        RECT 15.605000 170.550000 25.055000 170.610000 ;
        RECT 15.605000 170.610000 25.115000 189.515000 ;
        RECT 15.715000  94.200000 24.085000  94.310000 ;
        RECT 15.865000  94.050000 24.195000  94.200000 ;
        RECT 16.015000  93.900000 24.345000  94.050000 ;
        RECT 16.165000  93.750000 24.495000  93.900000 ;
        RECT 16.315000  93.600000 24.645000  93.750000 ;
        RECT 16.465000  93.450000 24.795000  93.600000 ;
        RECT 16.615000  93.300000 24.945000  93.450000 ;
        RECT 16.765000  93.150000 25.095000  93.300000 ;
        RECT 16.915000  93.000000 25.245000  93.150000 ;
        RECT 17.065000  92.850000 25.395000  93.000000 ;
        RECT 17.215000  92.700000 25.545000  92.850000 ;
        RECT 17.365000  92.550000 25.695000  92.700000 ;
        RECT 17.515000  92.400000 25.845000  92.550000 ;
        RECT 17.665000  92.250000 25.995000  92.400000 ;
        RECT 17.815000  92.100000 26.145000  92.250000 ;
        RECT 17.965000  91.950000 26.295000  92.100000 ;
        RECT 18.115000  91.800000 26.445000  91.950000 ;
        RECT 18.265000  91.650000 26.595000  91.800000 ;
        RECT 18.415000  91.500000 26.745000  91.650000 ;
        RECT 18.565000  91.350000 26.895000  91.500000 ;
        RECT 18.715000  91.200000 27.045000  91.350000 ;
        RECT 18.865000  91.050000 27.195000  91.200000 ;
        RECT 19.015000  90.900000 27.345000  91.050000 ;
        RECT 19.165000  90.750000 27.495000  90.900000 ;
        RECT 19.315000  90.600000 27.645000  90.750000 ;
        RECT 19.465000  90.450000 27.795000  90.600000 ;
        RECT 19.615000  90.300000 27.945000  90.450000 ;
        RECT 19.765000  90.150000 28.095000  90.300000 ;
        RECT 19.915000  90.000000 28.245000  90.150000 ;
        RECT 20.065000  89.850000 28.395000  90.000000 ;
        RECT 20.215000  89.700000 28.545000  89.850000 ;
        RECT 20.365000  89.550000 28.695000  89.700000 ;
        RECT 20.515000  89.400000 28.845000  89.550000 ;
        RECT 20.665000  89.250000 28.995000  89.400000 ;
        RECT 20.815000  89.100000 29.145000  89.250000 ;
        RECT 20.965000  88.950000 29.295000  89.100000 ;
        RECT 21.115000  88.800000 29.445000  88.950000 ;
        RECT 21.265000  88.650000 29.595000  88.800000 ;
        RECT 21.415000  88.500000 29.745000  88.650000 ;
        RECT 21.565000  88.350000 29.895000  88.500000 ;
        RECT 21.715000  88.200000 30.045000  88.350000 ;
        RECT 21.865000  88.050000 30.195000  88.200000 ;
        RECT 22.015000  87.900000 30.345000  88.050000 ;
        RECT 22.165000  87.750000 30.495000  87.900000 ;
        RECT 22.315000  87.600000 30.645000  87.750000 ;
        RECT 22.465000  87.450000 30.795000  87.600000 ;
        RECT 22.615000  87.300000 30.945000  87.450000 ;
        RECT 22.765000  87.150000 31.095000  87.300000 ;
        RECT 22.915000  87.000000 31.245000  87.150000 ;
        RECT 23.065000  86.850000 31.395000  87.000000 ;
        RECT 23.215000  86.700000 31.545000  86.850000 ;
        RECT 23.365000  86.550000 31.695000  86.700000 ;
        RECT 23.515000  86.400000 31.845000  86.550000 ;
        RECT 23.665000  86.250000 31.995000  86.400000 ;
        RECT 23.670000  86.245000 32.145000  86.250000 ;
        RECT 23.760000  86.155000 32.145000  86.245000 ;
        RECT 23.850000  84.650000 32.165000  84.670000 ;
        RECT 23.850000  84.670000 32.145000  84.690000 ;
        RECT 23.850000  84.690000 32.145000  86.065000 ;
        RECT 23.850000  86.065000 32.145000  86.155000 ;
        RECT 23.920000  84.580000 32.185000  84.650000 ;
        RECT 24.070000  84.430000 32.255000  84.580000 ;
        RECT 24.220000  84.280000 32.405000  84.430000 ;
        RECT 24.370000  84.130000 32.555000  84.280000 ;
        RECT 24.520000  83.980000 32.705000  84.130000 ;
        RECT 24.650000  83.850000 48.870000  83.980000 ;
        RECT 24.800000  83.700000 48.870000  83.850000 ;
        RECT 24.950000  83.550000 48.870000  83.700000 ;
        RECT 25.100000  83.400000 48.870000  83.550000 ;
        RECT 25.250000  83.250000 48.870000  83.400000 ;
        RECT 25.400000  83.100000 48.870000  83.250000 ;
        RECT 25.550000  82.950000 48.870000  83.100000 ;
        RECT 25.700000  82.800000 48.870000  82.950000 ;
        RECT 25.850000  82.650000 48.870000  82.800000 ;
        RECT 26.000000   0.000000 36.880000  71.105000 ;
        RECT 26.000000  71.105000 36.880000  71.255000 ;
        RECT 26.000000  71.255000 37.030000  71.405000 ;
        RECT 26.000000  71.405000 37.180000  71.555000 ;
        RECT 26.000000  71.555000 37.330000  71.705000 ;
        RECT 26.000000  71.705000 37.480000  71.855000 ;
        RECT 26.000000  71.855000 37.630000  72.005000 ;
        RECT 26.000000  72.005000 37.780000  72.155000 ;
        RECT 26.000000  72.155000 37.930000  72.305000 ;
        RECT 26.000000  72.305000 38.080000  72.455000 ;
        RECT 26.000000  72.455000 38.230000  72.605000 ;
        RECT 26.000000  72.605000 38.380000  72.755000 ;
        RECT 26.000000  72.755000 38.530000  72.905000 ;
        RECT 26.000000  72.905000 38.680000  73.055000 ;
        RECT 26.000000  73.055000 38.830000  73.205000 ;
        RECT 26.000000  73.205000 38.980000  73.355000 ;
        RECT 26.000000  73.355000 39.130000  73.505000 ;
        RECT 26.000000  73.505000 39.280000  73.655000 ;
        RECT 26.000000  73.655000 39.430000  73.805000 ;
        RECT 26.000000  73.805000 39.580000  73.955000 ;
        RECT 26.000000  73.955000 39.730000  74.105000 ;
        RECT 26.000000  74.105000 39.880000  74.255000 ;
        RECT 26.000000  74.255000 40.030000  74.405000 ;
        RECT 26.000000  74.405000 40.180000  74.555000 ;
        RECT 26.000000  74.555000 40.330000  74.705000 ;
        RECT 26.000000  74.705000 40.480000  74.740000 ;
        RECT 26.000000  74.740000 46.795000  74.890000 ;
        RECT 26.000000  74.890000 46.945000  75.040000 ;
        RECT 26.000000  75.040000 47.095000  75.190000 ;
        RECT 26.000000  75.190000 47.245000  75.340000 ;
        RECT 26.000000  75.340000 47.395000  75.490000 ;
        RECT 26.000000  75.490000 47.545000  75.640000 ;
        RECT 26.000000  75.640000 47.695000  75.790000 ;
        RECT 26.000000  75.790000 47.845000  75.940000 ;
        RECT 26.000000  75.940000 47.995000  76.090000 ;
        RECT 26.000000  76.090000 48.145000  76.240000 ;
        RECT 26.000000  76.240000 48.295000  76.390000 ;
        RECT 26.000000  76.390000 48.445000  76.540000 ;
        RECT 26.000000  76.540000 48.595000  76.690000 ;
        RECT 26.000000  76.690000 48.745000  76.815000 ;
        RECT 26.000000  76.815000 48.870000  82.500000 ;
        RECT 26.000000  82.500000 48.870000  82.650000 ;
        RECT 26.035000  94.500000 32.035000 162.570000 ;
        RECT 26.035000 162.570000 32.035000 162.720000 ;
        RECT 26.035000 162.720000 32.185000 162.870000 ;
        RECT 26.035000 162.870000 32.335000 163.020000 ;
        RECT 26.035000 163.020000 32.485000 163.170000 ;
        RECT 26.035000 163.170000 32.635000 163.320000 ;
        RECT 26.035000 163.320000 32.785000 163.470000 ;
        RECT 26.035000 163.470000 32.935000 163.620000 ;
        RECT 26.035000 163.620000 33.085000 163.770000 ;
        RECT 26.035000 163.770000 33.235000 163.920000 ;
        RECT 26.035000 163.920000 33.385000 164.070000 ;
        RECT 26.035000 164.070000 33.535000 164.220000 ;
        RECT 26.035000 164.220000 33.685000 164.370000 ;
        RECT 26.035000 164.370000 33.835000 164.520000 ;
        RECT 26.035000 164.520000 33.985000 164.670000 ;
        RECT 26.035000 164.670000 34.135000 164.820000 ;
        RECT 26.035000 164.820000 34.285000 164.970000 ;
        RECT 26.035000 164.970000 34.435000 165.120000 ;
        RECT 26.035000 165.120000 34.585000 165.270000 ;
        RECT 26.035000 165.270000 34.735000 165.420000 ;
        RECT 26.035000 165.420000 34.885000 165.570000 ;
        RECT 26.035000 165.570000 35.035000 165.720000 ;
        RECT 26.035000 165.720000 35.185000 165.870000 ;
        RECT 26.035000 165.870000 35.335000 166.020000 ;
        RECT 26.035000 166.020000 35.485000 166.170000 ;
        RECT 26.035000 166.170000 35.635000 166.320000 ;
        RECT 26.035000 166.320000 35.785000 166.470000 ;
        RECT 26.035000 166.470000 35.935000 166.620000 ;
        RECT 26.035000 166.620000 36.085000 166.770000 ;
        RECT 26.035000 166.770000 36.235000 166.920000 ;
        RECT 26.035000 166.920000 36.385000 167.070000 ;
        RECT 26.035000 167.070000 36.535000 167.220000 ;
        RECT 26.035000 167.220000 36.685000 167.370000 ;
        RECT 26.035000 167.370000 36.835000 167.460000 ;
        RECT 26.035000 167.460000 36.925000 189.515000 ;
        RECT 26.095000  94.440000 32.035000  94.500000 ;
        RECT 26.245000  94.290000 32.035000  94.440000 ;
        RECT 26.395000  94.140000 32.035000  94.290000 ;
        RECT 26.545000  93.990000 32.035000  94.140000 ;
        RECT 26.695000  93.840000 32.035000  93.990000 ;
        RECT 26.845000  93.690000 32.035000  93.840000 ;
        RECT 26.995000  93.540000 32.035000  93.690000 ;
        RECT 27.145000  93.390000 32.035000  93.540000 ;
        RECT 27.160000  93.375000 32.035000  93.390000 ;
        RECT 27.310000  93.225000 32.050000  93.375000 ;
        RECT 27.460000  93.075000 32.200000  93.225000 ;
        RECT 27.610000  92.925000 32.350000  93.075000 ;
        RECT 27.760000  92.775000 32.500000  92.925000 ;
        RECT 27.910000  92.625000 32.650000  92.775000 ;
        RECT 28.060000  92.475000 32.800000  92.625000 ;
        RECT 28.210000  92.325000 32.950000  92.475000 ;
        RECT 28.360000  92.175000 33.100000  92.325000 ;
        RECT 28.510000  92.025000 33.250000  92.175000 ;
        RECT 28.660000  91.875000 33.400000  92.025000 ;
        RECT 28.810000  91.725000 33.550000  91.875000 ;
        RECT 28.960000  91.575000 33.700000  91.725000 ;
        RECT 29.110000  91.425000 33.850000  91.575000 ;
        RECT 29.260000  91.275000 34.000000  91.425000 ;
        RECT 29.410000  91.125000 34.150000  91.275000 ;
        RECT 29.560000  90.975000 34.300000  91.125000 ;
        RECT 29.710000  90.825000 34.450000  90.975000 ;
        RECT 29.860000  90.675000 34.600000  90.825000 ;
        RECT 30.010000  90.525000 34.750000  90.675000 ;
        RECT 30.160000  90.375000 34.900000  90.525000 ;
        RECT 30.175000  90.360000 42.385000  90.375000 ;
        RECT 30.325000  90.210000 42.235000  90.360000 ;
        RECT 30.475000  90.060000 42.085000  90.210000 ;
        RECT 30.625000  89.910000 41.935000  90.060000 ;
        RECT 30.775000  89.760000 41.785000  89.910000 ;
        RECT 30.925000  89.610000 41.635000  89.760000 ;
        RECT 31.075000  89.460000 41.485000  89.610000 ;
        RECT 31.225000  89.310000 41.335000  89.460000 ;
        RECT 31.375000  89.160000 41.185000  89.310000 ;
        RECT 31.525000  89.010000 41.035000  89.160000 ;
        RECT 31.675000  88.860000 40.885000  89.010000 ;
        RECT 31.825000  88.710000 40.735000  88.860000 ;
        RECT 31.975000  88.560000 40.585000  88.710000 ;
        RECT 32.125000  88.410000 40.435000  88.560000 ;
        RECT 32.275000  88.260000 40.285000  88.410000 ;
        RECT 32.425000  88.110000 40.135000  88.260000 ;
        RECT 32.575000  87.960000 39.985000  88.110000 ;
        RECT 32.725000  87.810000 39.835000  87.960000 ;
        RECT 32.875000  87.660000 39.685000  87.810000 ;
        RECT 33.025000  87.510000 39.535000  87.660000 ;
        RECT 33.175000  87.360000 39.385000  87.510000 ;
        RECT 33.305000  87.230000 39.385000  87.360000 ;
        RECT 33.455000  87.080000 39.385000  87.230000 ;
        RECT 33.605000  86.930000 39.385000  87.080000 ;
        RECT 33.755000  86.780000 39.385000  86.930000 ;
        RECT 33.905000  86.630000 39.385000  86.780000 ;
        RECT 33.945000  83.980000 39.945000  84.130000 ;
        RECT 34.055000  86.480000 39.385000  86.630000 ;
        RECT 34.095000  84.130000 39.795000  84.280000 ;
        RECT 34.205000  86.330000 39.385000  86.480000 ;
        RECT 34.245000  84.280000 39.645000  84.430000 ;
        RECT 34.355000  86.180000 39.385000  86.330000 ;
        RECT 34.395000  84.430000 39.495000  84.580000 ;
        RECT 34.505000  84.580000 39.385000  84.690000 ;
        RECT 34.505000  84.690000 39.385000  86.030000 ;
        RECT 34.505000  86.030000 39.385000  86.180000 ;
        RECT 37.945000  90.375000 42.400000  90.525000 ;
        RECT 37.945000 169.025000 48.835000 189.515000 ;
        RECT 38.035000 168.935000 48.835000 169.025000 ;
        RECT 38.095000  90.525000 42.550000  90.675000 ;
        RECT 38.185000 168.785000 48.835000 168.935000 ;
        RECT 38.245000  90.675000 42.700000  90.825000 ;
        RECT 38.335000 168.635000 48.835000 168.785000 ;
        RECT 38.395000  90.825000 42.850000  90.975000 ;
        RECT 38.485000 168.485000 48.835000 168.635000 ;
        RECT 38.545000  90.975000 43.000000  91.125000 ;
        RECT 38.635000 168.335000 48.835000 168.485000 ;
        RECT 38.695000  91.125000 43.150000  91.275000 ;
        RECT 38.785000 168.185000 48.835000 168.335000 ;
        RECT 38.845000  91.275000 43.300000  91.425000 ;
        RECT 38.935000 168.035000 48.835000 168.185000 ;
        RECT 38.995000  91.425000 43.450000  91.575000 ;
        RECT 39.085000 167.885000 48.835000 168.035000 ;
        RECT 39.145000  91.575000 43.600000  91.725000 ;
        RECT 39.235000 167.735000 48.835000 167.885000 ;
        RECT 39.295000  91.725000 43.750000  91.875000 ;
        RECT 39.385000 167.585000 48.835000 167.735000 ;
        RECT 39.445000  91.875000 43.900000  92.025000 ;
        RECT 39.535000 167.435000 48.835000 167.585000 ;
        RECT 39.595000  92.025000 44.050000  92.175000 ;
        RECT 39.685000 167.285000 48.835000 167.435000 ;
        RECT 39.745000  92.175000 44.200000  92.325000 ;
        RECT 39.835000 167.135000 48.835000 167.285000 ;
        RECT 39.895000  92.325000 44.350000  92.475000 ;
        RECT 39.985000 166.985000 48.835000 167.135000 ;
        RECT 40.045000  92.475000 44.500000  92.625000 ;
        RECT 40.135000 166.835000 48.835000 166.985000 ;
        RECT 40.195000  92.625000 44.650000  92.775000 ;
        RECT 40.285000 166.685000 48.835000 166.835000 ;
        RECT 40.345000  92.775000 44.800000  92.925000 ;
        RECT 40.435000 166.535000 48.835000 166.685000 ;
        RECT 40.495000  92.925000 44.950000  93.075000 ;
        RECT 40.585000 166.385000 48.835000 166.535000 ;
        RECT 40.645000  93.075000 45.100000  93.225000 ;
        RECT 40.735000 166.235000 48.835000 166.385000 ;
        RECT 40.795000  93.225000 45.250000  93.375000 ;
        RECT 40.885000 166.085000 48.835000 166.235000 ;
        RECT 40.945000  93.375000 45.400000  93.525000 ;
        RECT 41.035000 165.935000 48.835000 166.085000 ;
        RECT 41.050000  83.980000 48.870000  84.130000 ;
        RECT 41.095000  93.525000 45.550000  93.675000 ;
        RECT 41.185000 165.785000 48.835000 165.935000 ;
        RECT 41.200000  84.130000 48.870000  84.280000 ;
        RECT 41.245000  93.675000 45.700000  93.825000 ;
        RECT 41.335000 165.635000 48.835000 165.785000 ;
        RECT 41.350000  84.280000 48.870000  84.430000 ;
        RECT 41.395000  93.825000 45.850000  93.975000 ;
        RECT 41.485000 165.485000 48.835000 165.635000 ;
        RECT 41.500000  84.430000 48.870000  84.580000 ;
        RECT 41.545000  93.975000 46.000000  94.125000 ;
        RECT 41.610000  84.580000 48.870000  84.690000 ;
        RECT 41.610000  84.690000 48.870000  84.810000 ;
        RECT 41.610000  84.810000 48.870000  84.960000 ;
        RECT 41.610000  84.960000 49.020000  85.110000 ;
        RECT 41.610000  85.110000 49.170000  85.260000 ;
        RECT 41.610000  85.260000 49.320000  85.410000 ;
        RECT 41.610000  85.410000 49.470000  85.560000 ;
        RECT 41.610000  85.560000 49.620000  85.710000 ;
        RECT 41.610000  85.710000 49.770000  85.860000 ;
        RECT 41.610000  85.860000 49.920000  86.010000 ;
        RECT 41.610000  86.010000 50.070000  86.160000 ;
        RECT 41.610000  86.160000 50.220000  86.310000 ;
        RECT 41.610000  86.310000 50.370000  86.460000 ;
        RECT 41.610000  86.460000 50.520000  86.610000 ;
        RECT 41.610000  86.610000 50.670000  86.760000 ;
        RECT 41.610000  86.760000 50.820000  86.910000 ;
        RECT 41.610000  86.910000 50.970000  86.960000 ;
        RECT 41.610000  86.960000 51.020000  87.445000 ;
        RECT 41.635000 165.335000 48.835000 165.485000 ;
        RECT 41.695000  94.125000 46.150000  94.275000 ;
        RECT 41.760000  87.445000 51.020000  87.595000 ;
        RECT 41.785000 165.185000 48.835000 165.335000 ;
        RECT 41.845000  94.275000 46.300000  94.425000 ;
        RECT 41.910000  87.595000 51.020000  87.745000 ;
        RECT 41.935000 165.035000 48.835000 165.185000 ;
        RECT 41.995000  94.425000 46.450000  94.575000 ;
        RECT 42.060000  87.745000 51.020000  87.895000 ;
        RECT 42.085000 164.885000 48.835000 165.035000 ;
        RECT 42.145000  94.575000 46.600000  94.725000 ;
        RECT 42.210000  87.895000 51.020000  88.045000 ;
        RECT 42.235000 164.735000 48.835000 164.885000 ;
        RECT 42.295000  94.725000 46.750000  94.875000 ;
        RECT 42.360000  88.045000 51.020000  88.195000 ;
        RECT 42.385000 164.585000 48.835000 164.735000 ;
        RECT 42.445000  94.875000 46.900000  95.025000 ;
        RECT 42.510000  88.195000 51.020000  88.345000 ;
        RECT 42.535000 164.435000 48.835000 164.585000 ;
        RECT 42.540000  88.345000 51.020000  88.375000 ;
        RECT 42.595000  95.025000 47.050000  95.175000 ;
        RECT 42.685000 164.285000 48.835000 164.435000 ;
        RECT 42.690000  88.375000 51.020000  88.525000 ;
        RECT 42.745000  95.175000 47.200000  95.325000 ;
        RECT 42.835000  95.325000 47.350000  95.415000 ;
        RECT 42.835000  95.415000 47.440000  95.565000 ;
        RECT 42.835000  95.565000 47.590000  95.715000 ;
        RECT 42.835000  95.715000 47.740000  95.865000 ;
        RECT 42.835000  95.865000 47.890000  96.015000 ;
        RECT 42.835000  96.015000 48.040000  96.165000 ;
        RECT 42.835000  96.165000 48.190000  96.315000 ;
        RECT 42.835000  96.315000 48.340000  96.465000 ;
        RECT 42.835000  96.465000 48.490000  96.615000 ;
        RECT 42.835000  96.615000 48.640000  96.765000 ;
        RECT 42.835000  96.765000 48.790000  96.810000 ;
        RECT 42.835000  96.810000 48.835000 164.135000 ;
        RECT 42.835000 164.135000 48.835000 164.285000 ;
        RECT 42.840000  88.525000 51.170000  88.675000 ;
        RECT 42.990000  88.675000 51.320000  88.825000 ;
        RECT 43.140000  88.825000 51.470000  88.975000 ;
        RECT 43.290000  88.975000 51.620000  89.125000 ;
        RECT 43.440000  89.125000 51.770000  89.275000 ;
        RECT 43.590000  89.275000 51.920000  89.425000 ;
        RECT 43.740000  89.425000 52.070000  89.575000 ;
        RECT 43.890000  89.575000 52.220000  89.725000 ;
        RECT 44.040000  89.725000 52.370000  89.875000 ;
        RECT 44.190000  89.875000 52.520000  90.025000 ;
        RECT 44.340000  90.025000 52.670000  90.175000 ;
        RECT 44.490000  90.175000 52.820000  90.325000 ;
        RECT 44.640000  90.325000 52.970000  90.475000 ;
        RECT 44.790000  90.475000 53.120000  90.625000 ;
        RECT 44.940000  90.625000 53.270000  90.775000 ;
        RECT 45.090000  90.775000 53.420000  90.925000 ;
        RECT 45.240000  90.925000 53.570000  91.075000 ;
        RECT 45.390000  91.075000 53.720000  91.225000 ;
        RECT 45.540000  91.225000 53.870000  91.375000 ;
        RECT 45.690000  91.375000 54.020000  91.525000 ;
        RECT 45.840000  91.525000 54.170000  91.675000 ;
        RECT 45.990000  91.675000 54.320000  91.825000 ;
        RECT 46.140000  91.825000 54.470000  91.975000 ;
        RECT 46.290000  91.975000 54.620000  92.125000 ;
        RECT 46.440000  92.125000 54.770000  92.275000 ;
        RECT 46.590000  92.275000 54.920000  92.425000 ;
        RECT 46.740000  92.425000 55.070000  92.575000 ;
        RECT 46.890000  92.575000 55.220000  92.725000 ;
        RECT 47.040000  92.725000 55.370000  92.875000 ;
        RECT 47.190000  92.875000 55.520000  93.025000 ;
        RECT 47.340000  93.025000 55.670000  93.175000 ;
        RECT 47.490000  93.175000 55.820000  93.325000 ;
        RECT 47.640000  93.325000 55.970000  93.475000 ;
        RECT 47.790000  93.475000 56.120000  93.625000 ;
        RECT 47.940000  93.625000 56.270000  93.775000 ;
        RECT 48.090000  93.775000 56.420000  93.925000 ;
        RECT 48.240000  93.925000 56.570000  94.075000 ;
        RECT 48.390000  94.075000 56.720000  94.225000 ;
        RECT 48.540000  94.225000 56.870000  94.375000 ;
        RECT 48.690000  94.375000 57.020000  94.525000 ;
        RECT 48.840000  94.525000 57.170000  94.675000 ;
        RECT 48.990000  94.675000 57.320000  94.825000 ;
        RECT 49.140000  94.825000 57.470000  94.975000 ;
        RECT 49.290000  94.975000 57.620000  95.125000 ;
        RECT 49.440000  95.125000 57.770000  95.275000 ;
        RECT 49.590000  95.275000 57.920000  95.425000 ;
        RECT 49.740000  95.425000 58.070000  95.575000 ;
        RECT 49.870000 168.920000 60.330000 189.515000 ;
        RECT 49.890000  95.575000 58.220000  95.725000 ;
        RECT 49.980000 168.810000 60.330000 168.920000 ;
        RECT 50.040000  95.725000 58.370000  95.875000 ;
        RECT 50.130000 168.660000 60.330000 168.810000 ;
        RECT 50.190000  95.875000 58.520000  96.025000 ;
        RECT 50.280000 168.510000 60.330000 168.660000 ;
        RECT 50.340000  96.025000 58.670000  96.175000 ;
        RECT 50.430000 168.360000 60.330000 168.510000 ;
        RECT 50.490000  96.175000 58.820000  96.325000 ;
        RECT 50.580000 168.210000 60.330000 168.360000 ;
        RECT 50.640000  96.325000 58.970000  96.475000 ;
        RECT 50.730000 168.060000 60.330000 168.210000 ;
        RECT 50.790000  96.475000 59.120000  96.625000 ;
        RECT 50.880000 167.910000 60.330000 168.060000 ;
        RECT 50.940000  96.625000 59.270000  96.775000 ;
        RECT 51.030000 167.760000 60.330000 167.910000 ;
        RECT 51.090000  96.775000 59.420000  96.925000 ;
        RECT 51.180000 167.610000 60.330000 167.760000 ;
        RECT 51.240000  96.925000 59.570000  97.075000 ;
        RECT 51.330000 167.460000 60.330000 167.610000 ;
        RECT 51.390000  97.075000 59.720000  97.225000 ;
        RECT 51.480000 167.310000 60.330000 167.460000 ;
        RECT 51.540000  97.225000 59.870000  97.375000 ;
        RECT 51.630000 167.160000 60.330000 167.310000 ;
        RECT 51.690000  97.375000 60.020000  97.525000 ;
        RECT 51.780000 167.010000 60.330000 167.160000 ;
        RECT 51.840000  97.525000 60.170000  97.675000 ;
        RECT 51.850000  97.675000 60.320000  97.685000 ;
        RECT 51.930000 166.860000 60.330000 167.010000 ;
        RECT 52.000000  97.685000 60.330000  97.835000 ;
        RECT 52.080000 166.710000 60.330000 166.860000 ;
        RECT 52.150000  97.835000 60.330000  97.985000 ;
        RECT 52.230000 166.560000 60.330000 166.710000 ;
        RECT 52.300000  97.985000 60.330000  98.135000 ;
        RECT 52.380000 166.410000 60.330000 166.560000 ;
        RECT 52.450000  98.135000 60.330000  98.285000 ;
        RECT 52.530000 166.260000 60.330000 166.410000 ;
        RECT 52.600000  98.285000 60.330000  98.435000 ;
        RECT 52.680000 166.110000 60.330000 166.260000 ;
        RECT 52.750000  98.435000 60.330000  98.585000 ;
        RECT 52.830000 165.960000 60.330000 166.110000 ;
        RECT 52.900000  98.585000 60.330000  98.735000 ;
        RECT 52.980000 165.810000 60.330000 165.960000 ;
        RECT 53.050000  98.735000 60.330000  98.885000 ;
        RECT 53.130000 165.660000 60.330000 165.810000 ;
        RECT 53.200000  98.885000 60.330000  99.035000 ;
        RECT 53.280000 165.510000 60.330000 165.660000 ;
        RECT 53.350000  99.035000 60.330000  99.185000 ;
        RECT 53.430000 165.360000 60.330000 165.510000 ;
        RECT 53.500000  99.185000 60.330000  99.335000 ;
        RECT 53.580000 165.210000 60.330000 165.360000 ;
        RECT 53.650000  99.335000 60.330000  99.485000 ;
        RECT 53.730000 165.060000 60.330000 165.210000 ;
        RECT 53.800000  99.485000 60.330000  99.635000 ;
        RECT 53.880000 164.910000 60.330000 165.060000 ;
        RECT 53.950000  99.635000 60.330000  99.785000 ;
        RECT 54.030000 164.760000 60.330000 164.910000 ;
        RECT 54.100000  99.785000 60.330000  99.935000 ;
        RECT 54.180000 164.610000 60.330000 164.760000 ;
        RECT 54.250000  99.935000 60.330000 100.085000 ;
        RECT 54.330000 100.085000 60.330000 100.165000 ;
        RECT 54.330000 100.165000 60.330000 164.460000 ;
        RECT 54.330000 164.460000 60.330000 164.610000 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380000 0.000000 49.255000 69.490000 ;
    END
  END DRN_LVC2
  PIN G_CORE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.500000  0.000000 24.500000  82.660000 ;
        RECT 0.500000 82.660000 24.350000  82.810000 ;
        RECT 0.500000 82.810000 24.200000  82.960000 ;
        RECT 0.500000 82.960000 24.050000  83.110000 ;
        RECT 0.500000 83.110000 23.900000  83.260000 ;
        RECT 0.500000 83.260000 23.750000  83.410000 ;
        RECT 0.500000 83.410000 23.600000  83.560000 ;
        RECT 0.500000 83.560000 23.450000  83.710000 ;
        RECT 0.500000 83.710000 23.300000  83.860000 ;
        RECT 0.500000 83.860000 23.150000  84.010000 ;
        RECT 0.500000 84.010000 23.000000  84.160000 ;
        RECT 0.500000 84.160000 22.850000  84.310000 ;
        RECT 0.500000 84.310000 22.700000  84.460000 ;
        RECT 0.500000 84.460000 22.550000  84.610000 ;
        RECT 0.500000 84.610000 22.400000  84.760000 ;
        RECT 0.500000 84.760000 22.250000  84.910000 ;
        RECT 0.500000 84.910000 22.100000  85.060000 ;
        RECT 0.500000 85.060000 21.950000  85.210000 ;
        RECT 0.500000 85.210000 21.800000  85.360000 ;
        RECT 0.500000 85.360000 21.650000  85.510000 ;
        RECT 0.500000 85.510000 21.500000  85.660000 ;
        RECT 0.500000 85.660000 21.350000  85.810000 ;
        RECT 0.500000 85.810000 21.200000  85.960000 ;
        RECT 0.500000 85.960000 21.050000  86.110000 ;
        RECT 0.500000 86.110000 20.900000  86.260000 ;
        RECT 0.500000 86.260000 20.750000  86.410000 ;
        RECT 0.500000 86.410000 20.600000  86.560000 ;
        RECT 0.500000 86.560000 20.450000  86.710000 ;
        RECT 0.500000 86.710000 20.300000  86.860000 ;
        RECT 0.500000 86.860000 20.150000  87.010000 ;
        RECT 0.500000 87.010000 20.000000  87.160000 ;
        RECT 0.500000 87.160000 19.850000  87.310000 ;
        RECT 0.500000 87.310000 19.700000  87.460000 ;
        RECT 0.500000 87.460000 19.550000  87.610000 ;
        RECT 0.500000 87.610000 19.400000  87.760000 ;
        RECT 0.500000 87.760000 19.250000  87.910000 ;
        RECT 0.500000 87.910000 19.100000  88.060000 ;
        RECT 0.500000 88.060000 18.950000  88.210000 ;
        RECT 0.500000 88.210000 18.800000  88.360000 ;
        RECT 0.500000 88.360000 18.650000  88.510000 ;
        RECT 0.500000 88.510000 18.500000  88.660000 ;
        RECT 0.500000 88.660000 18.350000  88.810000 ;
        RECT 0.500000 88.810000 18.200000  88.960000 ;
        RECT 0.500000 88.960000 18.050000  89.110000 ;
        RECT 0.500000 89.110000 17.900000  89.260000 ;
        RECT 0.500000 89.260000 17.750000  89.410000 ;
        RECT 0.500000 89.410000 17.600000  89.560000 ;
        RECT 0.500000 89.560000 17.450000  89.710000 ;
        RECT 0.500000 89.710000 17.300000  89.860000 ;
        RECT 0.500000 89.860000 17.150000  90.010000 ;
        RECT 0.500000 90.010000 17.000000  90.160000 ;
        RECT 0.500000 90.160000 16.850000  90.310000 ;
        RECT 0.500000 90.310000 16.700000  90.460000 ;
        RECT 0.500000 90.460000 16.550000  90.610000 ;
        RECT 0.500000 90.610000 16.400000  90.760000 ;
        RECT 0.500000 90.760000 16.250000  90.910000 ;
        RECT 0.500000 90.910000 16.100000  91.060000 ;
        RECT 0.500000 91.060000 15.950000  91.210000 ;
        RECT 0.500000 91.210000 15.800000  91.360000 ;
        RECT 0.500000 91.360000 15.650000  91.510000 ;
        RECT 0.500000 91.510000 15.500000  91.660000 ;
        RECT 0.500000 91.660000 15.350000  91.810000 ;
        RECT 0.500000 91.810000 15.200000  91.960000 ;
        RECT 0.500000 91.960000 15.050000  92.110000 ;
        RECT 0.500000 92.110000 14.900000  92.260000 ;
        RECT 0.500000 92.260000 14.750000  92.410000 ;
        RECT 0.500000 92.410000 14.600000  92.560000 ;
        RECT 0.500000 92.560000 14.450000  92.710000 ;
        RECT 0.500000 92.710000 14.300000  92.860000 ;
        RECT 0.500000 92.860000 14.150000  93.010000 ;
        RECT 0.500000 93.010000 14.000000  93.160000 ;
        RECT 0.500000 93.160000 13.850000  93.310000 ;
        RECT 0.500000 93.310000 13.700000  93.460000 ;
        RECT 0.500000 93.460000 13.550000  93.610000 ;
        RECT 0.500000 93.610000 13.400000  93.760000 ;
        RECT 0.500000 93.760000 13.250000  93.910000 ;
        RECT 0.500000 93.910000 13.100000  94.060000 ;
        RECT 0.500000 94.060000 12.950000  94.210000 ;
        RECT 0.500000 94.210000 12.900000  94.260000 ;
        RECT 0.500000 94.260000 12.900000 171.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000  0.000000 74.700000  84.465000 ;
        RECT 50.905000 84.465000 74.700000  84.615000 ;
        RECT 51.055000 84.615000 74.700000  84.765000 ;
        RECT 51.205000 84.765000 74.700000  84.915000 ;
        RECT 51.355000 84.915000 74.700000  85.065000 ;
        RECT 51.505000 85.065000 74.700000  85.215000 ;
        RECT 51.655000 85.215000 74.700000  85.365000 ;
        RECT 51.805000 85.365000 74.700000  85.515000 ;
        RECT 51.955000 85.515000 74.700000  85.665000 ;
        RECT 52.105000 85.665000 74.700000  85.815000 ;
        RECT 52.255000 85.815000 74.700000  85.965000 ;
        RECT 52.405000 85.965000 74.700000  86.115000 ;
        RECT 52.555000 86.115000 74.700000  86.265000 ;
        RECT 52.705000 86.265000 74.700000  86.415000 ;
        RECT 52.855000 86.415000 74.700000  86.565000 ;
        RECT 53.005000 86.565000 74.700000  86.715000 ;
        RECT 53.155000 86.715000 74.700000  86.865000 ;
        RECT 53.305000 86.865000 74.700000  87.015000 ;
        RECT 53.455000 87.015000 74.700000  87.165000 ;
        RECT 53.605000 87.165000 74.700000  87.315000 ;
        RECT 53.755000 87.315000 74.700000  87.465000 ;
        RECT 53.905000 87.465000 74.700000  87.615000 ;
        RECT 54.055000 87.615000 74.700000  87.765000 ;
        RECT 54.205000 87.765000 74.700000  87.915000 ;
        RECT 54.355000 87.915000 74.700000  88.065000 ;
        RECT 54.505000 88.065000 74.700000  88.215000 ;
        RECT 54.655000 88.215000 74.700000  88.365000 ;
        RECT 54.805000 88.365000 74.700000  88.515000 ;
        RECT 54.955000 88.515000 74.700000  88.665000 ;
        RECT 55.105000 88.665000 74.700000  88.815000 ;
        RECT 55.255000 88.815000 74.700000  88.965000 ;
        RECT 55.405000 88.965000 74.700000  89.115000 ;
        RECT 55.555000 89.115000 74.700000  89.265000 ;
        RECT 55.705000 89.265000 74.700000  89.415000 ;
        RECT 55.855000 89.415000 74.700000  89.565000 ;
        RECT 56.005000 89.565000 74.700000  89.715000 ;
        RECT 56.155000 89.715000 74.700000  89.865000 ;
        RECT 56.305000 89.865000 74.700000  90.015000 ;
        RECT 56.455000 90.015000 74.700000  90.165000 ;
        RECT 56.605000 90.165000 74.700000  90.315000 ;
        RECT 56.755000 90.315000 74.700000  90.465000 ;
        RECT 56.905000 90.465000 74.700000  90.615000 ;
        RECT 57.055000 90.615000 74.700000  90.765000 ;
        RECT 57.205000 90.765000 74.700000  90.915000 ;
        RECT 57.355000 90.915000 74.700000  91.065000 ;
        RECT 57.505000 91.065000 74.700000  91.215000 ;
        RECT 57.655000 91.215000 74.700000  91.365000 ;
        RECT 57.805000 91.365000 74.700000  91.515000 ;
        RECT 57.955000 91.515000 74.700000  91.665000 ;
        RECT 58.105000 91.665000 74.700000  91.815000 ;
        RECT 58.255000 91.815000 74.700000  91.965000 ;
        RECT 58.405000 91.965000 74.700000  92.115000 ;
        RECT 58.555000 92.115000 74.700000  92.265000 ;
        RECT 58.705000 92.265000 74.700000  92.415000 ;
        RECT 58.855000 92.415000 74.700000  92.565000 ;
        RECT 59.005000 92.565000 74.700000  92.715000 ;
        RECT 59.155000 92.715000 74.700000  92.865000 ;
        RECT 59.305000 92.865000 74.700000  93.015000 ;
        RECT 59.455000 93.015000 74.700000  93.165000 ;
        RECT 59.605000 93.165000 74.700000  93.315000 ;
        RECT 59.755000 93.315000 74.700000  93.465000 ;
        RECT 59.905000 93.465000 74.700000  93.615000 ;
        RECT 60.055000 93.615000 74.700000  93.765000 ;
        RECT 60.205000 93.765000 74.700000  93.915000 ;
        RECT 60.355000 93.915000 74.700000  94.065000 ;
        RECT 60.505000 94.065000 74.700000  94.215000 ;
        RECT 60.655000 94.215000 74.700000  94.365000 ;
        RECT 60.805000 94.365000 74.700000  94.515000 ;
        RECT 60.955000 94.515000 74.700000  94.665000 ;
        RECT 61.105000 94.665000 74.700000  94.815000 ;
        RECT 61.255000 94.815000 74.700000  94.965000 ;
        RECT 61.405000 94.965000 74.700000  95.115000 ;
        RECT 61.555000 95.115000 74.700000  95.265000 ;
        RECT 61.705000 95.265000 74.700000  95.415000 ;
        RECT 61.855000 95.415000 74.700000  95.565000 ;
        RECT 62.005000 95.565000 74.700000  95.715000 ;
        RECT 62.045000 95.715000 74.700000  95.755000 ;
        RECT 62.045000 95.755000 74.700000 172.235000 ;
    END
  END G_CORE
  PIN OGC_LVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 26.210000 0.000000 27.700000 0.170000 ;
    END
  END OGC_LVC
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT  0.500000   0.000000 20.495000   1.485000 ;
        RECT  0.500000   1.485000 20.425000   1.555000 ;
        RECT  0.500000   1.555000 20.355000   1.625000 ;
        RECT  0.500000   1.625000 20.285000   1.695000 ;
        RECT  0.500000   1.695000 20.215000   1.765000 ;
        RECT  0.500000   1.765000 20.145000   1.835000 ;
        RECT  0.500000   1.835000 20.075000   1.905000 ;
        RECT  0.500000   1.905000 20.005000   1.975000 ;
        RECT  0.500000   1.975000 19.935000   2.045000 ;
        RECT  0.500000   2.045000 19.865000   2.115000 ;
        RECT  0.500000   2.115000 19.795000   2.185000 ;
        RECT  0.500000   2.185000 19.725000   2.255000 ;
        RECT  0.500000   2.255000 19.655000   2.325000 ;
        RECT  0.500000   2.325000 19.585000   2.395000 ;
        RECT  0.500000   2.395000 19.515000   2.465000 ;
        RECT  0.500000   2.465000 19.445000   2.535000 ;
        RECT  0.500000   2.535000 19.375000   2.605000 ;
        RECT  0.500000   2.605000 19.305000   2.675000 ;
        RECT  0.500000   2.675000 19.235000   2.745000 ;
        RECT  0.500000   2.745000 19.165000   2.815000 ;
        RECT  0.500000   2.815000 19.095000   2.885000 ;
        RECT  0.500000   2.885000 19.025000   2.955000 ;
        RECT  0.500000   2.955000 18.955000   3.025000 ;
        RECT  0.500000   3.025000 18.885000   3.095000 ;
        RECT  0.500000   3.095000 18.815000   3.165000 ;
        RECT  0.500000   3.165000 18.745000   3.235000 ;
        RECT  0.500000   3.235000 18.675000   3.305000 ;
        RECT  0.500000   3.305000 18.605000   3.375000 ;
        RECT  0.500000   3.375000 18.535000   3.445000 ;
        RECT  0.500000   3.445000 18.465000   3.515000 ;
        RECT  0.500000   3.515000 18.395000   3.585000 ;
        RECT  0.500000   3.585000 18.325000   3.655000 ;
        RECT  0.500000   3.655000 18.255000   3.725000 ;
        RECT  0.500000   3.725000 18.185000   3.795000 ;
        RECT  0.500000   3.795000 18.115000   3.865000 ;
        RECT  0.500000   3.865000 18.045000   3.935000 ;
        RECT  0.500000   3.935000 17.975000   4.005000 ;
        RECT  0.500000   4.005000 17.905000   4.075000 ;
        RECT  0.500000   4.075000 17.835000   4.145000 ;
        RECT  0.500000   4.145000 17.765000   4.215000 ;
        RECT  0.500000   4.215000 17.695000   4.285000 ;
        RECT  0.500000   4.285000 17.625000   4.355000 ;
        RECT  0.500000   4.355000 17.555000   4.425000 ;
        RECT  0.500000   4.425000 17.485000   4.495000 ;
        RECT  0.500000   4.495000 17.415000   4.565000 ;
        RECT  0.500000   4.565000 17.345000   4.635000 ;
        RECT  0.500000   4.635000 17.275000   4.705000 ;
        RECT  0.500000   4.705000 17.205000   4.775000 ;
        RECT  0.500000   4.775000 17.135000   4.845000 ;
        RECT  0.500000   4.845000 17.065000   4.915000 ;
        RECT  0.500000   4.915000 16.995000   4.985000 ;
        RECT  0.500000   4.985000 16.925000   5.055000 ;
        RECT  0.500000   5.055000 16.860000   5.120000 ;
        RECT  0.500000   5.120000 16.860000   7.655000 ;
        RECT  0.500000   7.655000 10.745000   7.725000 ;
        RECT  0.500000   7.725000 10.675000   7.795000 ;
        RECT  0.500000   7.795000 10.605000   7.865000 ;
        RECT  0.500000   7.865000 10.535000   7.935000 ;
        RECT  0.500000   7.935000 10.465000   8.005000 ;
        RECT  0.500000   8.005000 10.420000   8.050000 ;
        RECT  0.500000   8.050000 10.420000   9.820000 ;
        RECT  0.500000   9.820000 10.420000   9.890000 ;
        RECT  0.500000   9.890000 10.490000   9.960000 ;
        RECT  0.500000   9.960000 10.560000  10.030000 ;
        RECT  0.500000  10.030000 10.630000  10.100000 ;
        RECT  0.500000  10.100000 10.700000  10.170000 ;
        RECT  0.500000  10.170000 10.770000  10.215000 ;
        RECT  0.500000  10.215000 55.595000  17.080000 ;
        RECT  0.500000  17.080000 21.785000  17.150000 ;
        RECT  0.500000  17.150000 21.715000  17.220000 ;
        RECT  0.500000  17.220000 21.645000  17.290000 ;
        RECT  0.500000  17.290000 21.575000  17.360000 ;
        RECT  0.500000  17.360000 21.505000  17.430000 ;
        RECT  0.500000  17.430000 21.435000  17.500000 ;
        RECT  0.500000  17.500000 21.365000  17.570000 ;
        RECT  0.500000  17.570000 21.295000  17.640000 ;
        RECT  0.500000  17.640000 21.225000  17.710000 ;
        RECT  0.500000  17.710000 21.155000  17.780000 ;
        RECT  0.500000  17.780000 21.085000  17.850000 ;
        RECT  0.500000  17.850000 21.015000  17.920000 ;
        RECT  0.500000  17.920000 20.945000  17.990000 ;
        RECT  0.500000  17.990000 20.875000  18.060000 ;
        RECT  0.500000  18.060000 20.805000  18.130000 ;
        RECT  0.500000  18.130000 20.735000  18.200000 ;
        RECT  0.500000  18.200000 20.665000  18.270000 ;
        RECT  0.500000  18.270000 20.595000  18.340000 ;
        RECT  0.500000  18.340000 20.525000  18.410000 ;
        RECT  0.500000  18.410000 20.455000  18.480000 ;
        RECT  0.500000  18.480000 20.385000  18.550000 ;
        RECT  0.500000  18.550000 20.315000  18.620000 ;
        RECT  0.500000  18.620000 20.245000  18.690000 ;
        RECT  0.500000  18.690000 20.175000  18.760000 ;
        RECT  0.500000  18.760000 20.105000  18.830000 ;
        RECT  0.500000  18.830000 20.035000  18.900000 ;
        RECT  0.500000  18.900000 19.965000  18.970000 ;
        RECT  0.500000  18.970000 19.895000  19.040000 ;
        RECT  0.500000  19.040000 19.825000  19.110000 ;
        RECT  0.500000  19.110000 19.755000  19.180000 ;
        RECT  0.500000  19.180000 19.685000  19.250000 ;
        RECT  0.500000  19.250000 19.615000  19.320000 ;
        RECT  0.500000  19.320000 19.545000  19.390000 ;
        RECT  0.500000  19.390000 19.475000  19.460000 ;
        RECT  0.500000  19.460000 19.405000  19.530000 ;
        RECT  0.500000  19.530000 19.335000  19.600000 ;
        RECT  0.500000  19.600000 19.265000  19.670000 ;
        RECT  0.500000  19.670000 19.195000  19.740000 ;
        RECT  0.500000  19.740000 19.125000  19.810000 ;
        RECT  0.500000  19.810000 19.055000  19.880000 ;
        RECT  0.500000  19.880000 18.985000  19.950000 ;
        RECT  0.500000  19.950000 18.915000  20.020000 ;
        RECT  0.500000  20.020000 18.845000  20.090000 ;
        RECT  0.500000  20.090000 18.775000  20.160000 ;
        RECT  0.500000  20.160000 18.705000  20.230000 ;
        RECT  0.500000  20.230000 18.635000  20.300000 ;
        RECT  0.500000  20.300000 18.565000  20.370000 ;
        RECT  0.500000  20.370000 18.495000  20.440000 ;
        RECT  0.500000  20.440000 18.425000  20.510000 ;
        RECT  0.500000  20.510000 18.355000  20.580000 ;
        RECT  0.500000  20.580000 18.285000  20.650000 ;
        RECT  0.500000  20.650000 18.215000  20.720000 ;
        RECT  0.500000  20.720000 18.145000  20.790000 ;
        RECT  0.500000  20.790000 18.075000  20.860000 ;
        RECT  0.500000  20.860000 18.005000  20.930000 ;
        RECT  0.500000  20.930000 17.935000  21.000000 ;
        RECT  0.500000  21.000000 17.865000  21.070000 ;
        RECT  0.500000  21.070000 17.795000  21.140000 ;
        RECT  0.500000  21.140000 17.725000  21.210000 ;
        RECT  0.500000  21.210000 17.655000  21.280000 ;
        RECT  0.500000  21.280000 17.585000  21.350000 ;
        RECT  0.500000  21.350000 17.515000  21.420000 ;
        RECT  0.500000  21.420000 17.445000  21.490000 ;
        RECT  0.500000  21.490000 17.375000  21.560000 ;
        RECT  0.500000  21.560000 17.305000  21.630000 ;
        RECT  0.500000  21.630000 17.235000  21.700000 ;
        RECT  0.500000  21.700000 17.165000  21.770000 ;
        RECT  0.500000  21.770000 17.095000  21.840000 ;
        RECT  0.500000  21.840000 17.025000  21.910000 ;
        RECT  0.500000  21.910000 16.955000  21.980000 ;
        RECT  0.500000  21.980000 16.885000  22.050000 ;
        RECT  0.500000  22.050000 16.815000  22.120000 ;
        RECT  0.500000  22.120000 16.745000  22.190000 ;
        RECT  0.500000  22.190000 16.675000  22.260000 ;
        RECT  0.500000  22.260000 16.605000  22.330000 ;
        RECT  0.500000  22.330000 16.535000  22.400000 ;
        RECT  0.500000  22.400000 16.465000  22.470000 ;
        RECT  0.500000  22.470000 16.395000  22.540000 ;
        RECT  0.500000  22.540000 16.325000  22.610000 ;
        RECT  0.500000  22.610000 16.255000  22.680000 ;
        RECT  0.500000  22.680000 16.185000  22.750000 ;
        RECT  0.500000  22.750000 16.115000  22.820000 ;
        RECT  0.500000  22.820000 16.045000  22.890000 ;
        RECT  0.500000  22.890000 15.975000  22.960000 ;
        RECT  0.500000  22.960000 15.905000  23.030000 ;
        RECT  0.500000  23.030000 15.835000  23.100000 ;
        RECT  0.500000  23.100000 15.765000  23.170000 ;
        RECT  0.500000  23.170000 15.695000  23.240000 ;
        RECT  0.500000  23.240000 15.625000  23.310000 ;
        RECT  0.500000  23.310000 15.555000  23.380000 ;
        RECT  0.500000  23.380000 15.485000  23.450000 ;
        RECT  0.500000  23.450000 15.415000  23.520000 ;
        RECT  0.500000  23.520000 15.345000  23.590000 ;
        RECT  0.500000  23.590000 15.275000  23.660000 ;
        RECT  0.500000  23.660000 15.205000  23.730000 ;
        RECT  0.500000  23.730000 15.135000  23.800000 ;
        RECT  0.500000  23.800000 15.065000  23.870000 ;
        RECT  0.500000  23.870000 14.995000  23.940000 ;
        RECT  0.500000  23.940000 14.925000  24.010000 ;
        RECT  0.500000  24.010000 14.855000  24.080000 ;
        RECT  0.500000  24.080000 14.785000  24.150000 ;
        RECT  0.500000  24.150000 14.715000  24.220000 ;
        RECT  0.500000  24.220000 14.645000  24.290000 ;
        RECT  0.500000  24.290000 14.575000  24.360000 ;
        RECT  0.500000  24.360000 14.505000  24.430000 ;
        RECT  0.500000  24.430000 14.435000  24.500000 ;
        RECT  0.500000  24.500000 14.365000  24.570000 ;
        RECT  0.500000  24.570000 14.295000  24.640000 ;
        RECT  0.500000  24.640000 14.225000  24.710000 ;
        RECT  0.500000  24.710000 14.155000  24.780000 ;
        RECT  0.500000  24.780000 14.085000  24.850000 ;
        RECT  0.500000  24.850000 14.015000  24.920000 ;
        RECT  0.500000  24.920000 13.945000  24.990000 ;
        RECT  0.500000  24.990000 13.875000  25.060000 ;
        RECT  0.500000  25.060000 13.805000  25.130000 ;
        RECT  0.500000  25.130000 13.750000  25.185000 ;
        RECT  0.500000  25.185000 13.750000  74.295000 ;
        RECT  0.500000  74.295000 13.750000  74.365000 ;
        RECT  0.500000  74.365000 13.820000  74.435000 ;
        RECT  0.500000  74.435000 13.890000  74.505000 ;
        RECT  0.500000  74.505000 13.960000 129.935000 ;
        RECT  0.500000 129.935000 13.960000 130.005000 ;
        RECT  0.500000 130.005000 14.030000 130.075000 ;
        RECT  0.500000 130.075000 14.100000 130.145000 ;
        RECT  0.500000 130.145000 14.170000 130.215000 ;
        RECT  0.500000 130.215000 14.240000 130.285000 ;
        RECT  0.500000 130.285000 14.310000 130.355000 ;
        RECT  0.500000 130.355000 14.380000 130.425000 ;
        RECT  0.500000 130.425000 14.450000 130.495000 ;
        RECT  0.500000 130.495000 14.520000 130.565000 ;
        RECT  0.500000 130.565000 14.590000 130.635000 ;
        RECT  0.500000 130.635000 14.660000 130.705000 ;
        RECT  0.500000 130.705000 14.730000 130.775000 ;
        RECT  0.500000 130.775000 14.800000 130.845000 ;
        RECT  0.500000 130.845000 14.870000 130.915000 ;
        RECT  0.500000 130.915000 14.940000 130.985000 ;
        RECT  0.500000 130.985000 68.010000 133.630000 ;
        RECT  0.500000 133.630000 14.940000 133.700000 ;
        RECT  0.500000 133.700000 14.870000 133.770000 ;
        RECT  0.500000 133.770000 14.800000 133.840000 ;
        RECT  0.500000 133.840000 14.730000 133.910000 ;
        RECT  0.500000 133.910000 14.660000 133.980000 ;
        RECT  0.500000 133.980000 14.590000 134.050000 ;
        RECT  0.500000 134.050000 14.520000 134.120000 ;
        RECT  0.500000 134.120000 14.450000 134.190000 ;
        RECT  0.500000 134.190000 14.380000 134.260000 ;
        RECT  0.500000 134.260000 14.310000 134.330000 ;
        RECT  0.500000 134.330000 14.240000 134.400000 ;
        RECT  0.500000 134.400000 14.170000 134.470000 ;
        RECT  0.500000 134.470000 14.100000 134.540000 ;
        RECT  0.500000 134.540000 14.030000 134.610000 ;
        RECT  0.500000 134.610000 13.960000 134.680000 ;
        RECT  0.500000 134.680000 13.960000 139.940000 ;
        RECT  0.500000 139.940000 13.960000 140.010000 ;
        RECT  0.500000 140.010000 14.030000 140.080000 ;
        RECT  0.500000 140.080000 14.100000 140.150000 ;
        RECT  0.500000 140.150000 14.170000 140.220000 ;
        RECT  0.500000 140.220000 14.240000 140.290000 ;
        RECT  0.500000 140.290000 14.310000 140.360000 ;
        RECT  0.500000 140.360000 14.380000 140.430000 ;
        RECT  0.500000 140.430000 14.450000 140.500000 ;
        RECT  0.500000 140.500000 14.520000 140.570000 ;
        RECT  0.500000 140.570000 14.590000 140.640000 ;
        RECT  0.500000 140.640000 14.660000 140.710000 ;
        RECT  0.500000 140.710000 14.730000 140.780000 ;
        RECT  0.500000 140.780000 14.800000 140.850000 ;
        RECT  0.500000 140.850000 14.870000 140.920000 ;
        RECT  0.500000 140.920000 14.940000 140.990000 ;
        RECT  0.500000 140.990000 68.010000 143.630000 ;
        RECT  0.500000 143.630000 14.940000 143.700000 ;
        RECT  0.500000 143.700000 14.870000 143.770000 ;
        RECT  0.500000 143.770000 14.800000 143.840000 ;
        RECT  0.500000 143.840000 14.730000 143.910000 ;
        RECT  0.500000 143.910000 14.660000 143.980000 ;
        RECT  0.500000 143.980000 14.590000 144.050000 ;
        RECT  0.500000 144.050000 14.520000 144.120000 ;
        RECT  0.500000 144.120000 14.450000 144.190000 ;
        RECT  0.500000 144.190000 14.380000 144.260000 ;
        RECT  0.500000 144.260000 14.310000 144.330000 ;
        RECT  0.500000 144.330000 14.240000 144.400000 ;
        RECT  0.500000 144.400000 14.170000 144.470000 ;
        RECT  0.500000 144.470000 14.100000 144.540000 ;
        RECT  0.500000 144.540000 14.030000 144.610000 ;
        RECT  0.500000 144.610000 13.960000 144.680000 ;
        RECT  0.500000 144.680000 13.960000 149.940000 ;
        RECT  0.500000 149.940000 13.960000 150.010000 ;
        RECT  0.500000 150.010000 14.030000 150.080000 ;
        RECT  0.500000 150.080000 14.100000 150.150000 ;
        RECT  0.500000 150.150000 14.170000 150.220000 ;
        RECT  0.500000 150.220000 14.240000 150.290000 ;
        RECT  0.500000 150.290000 14.310000 150.360000 ;
        RECT  0.500000 150.360000 14.380000 150.430000 ;
        RECT  0.500000 150.430000 14.450000 150.500000 ;
        RECT  0.500000 150.500000 14.520000 150.570000 ;
        RECT  0.500000 150.570000 14.590000 150.640000 ;
        RECT  0.500000 150.640000 14.660000 150.710000 ;
        RECT  0.500000 150.710000 14.730000 150.780000 ;
        RECT  0.500000 150.780000 14.800000 150.850000 ;
        RECT  0.500000 150.850000 14.870000 150.920000 ;
        RECT  0.500000 150.920000 14.940000 150.990000 ;
        RECT  0.500000 150.990000 68.010000 153.630000 ;
        RECT  0.500000 153.630000 14.940000 153.700000 ;
        RECT  0.500000 153.700000 14.870000 153.770000 ;
        RECT  0.500000 153.770000 14.800000 153.840000 ;
        RECT  0.500000 153.840000 14.730000 153.910000 ;
        RECT  0.500000 153.910000 14.660000 153.980000 ;
        RECT  0.500000 153.980000 14.590000 154.050000 ;
        RECT  0.500000 154.050000 14.520000 154.120000 ;
        RECT  0.500000 154.120000 14.450000 154.190000 ;
        RECT  0.500000 154.190000 14.380000 154.260000 ;
        RECT  0.500000 154.260000 14.310000 154.330000 ;
        RECT  0.500000 154.330000 14.240000 154.400000 ;
        RECT  0.500000 154.400000 14.170000 154.470000 ;
        RECT  0.500000 154.470000 14.100000 154.540000 ;
        RECT  0.500000 154.540000 14.030000 154.610000 ;
        RECT  0.500000 154.610000 13.960000 154.680000 ;
        RECT  0.500000 154.680000 13.960000 159.940000 ;
        RECT  0.500000 159.940000 13.960000 160.010000 ;
        RECT  0.500000 160.010000 14.030000 160.080000 ;
        RECT  0.500000 160.080000 14.100000 160.150000 ;
        RECT  0.500000 160.150000 14.170000 160.220000 ;
        RECT  0.500000 160.220000 14.240000 160.290000 ;
        RECT  0.500000 160.290000 14.310000 160.360000 ;
        RECT  0.500000 160.360000 14.380000 160.430000 ;
        RECT  0.500000 160.430000 14.450000 160.500000 ;
        RECT  0.500000 160.500000 14.520000 160.570000 ;
        RECT  0.500000 160.570000 14.590000 160.640000 ;
        RECT  0.500000 160.640000 14.660000 160.710000 ;
        RECT  0.500000 160.710000 14.730000 160.780000 ;
        RECT  0.500000 160.780000 14.800000 160.850000 ;
        RECT  0.500000 160.850000 14.870000 160.920000 ;
        RECT  0.500000 160.920000 14.940000 160.990000 ;
        RECT  0.500000 160.990000 68.010000 163.630000 ;
        RECT  0.500000 163.630000 14.940000 163.700000 ;
        RECT  0.500000 163.700000 14.870000 163.770000 ;
        RECT  0.500000 163.770000 14.800000 163.840000 ;
        RECT  0.500000 163.840000 14.730000 163.910000 ;
        RECT  0.500000 163.910000 14.660000 163.980000 ;
        RECT  0.500000 163.980000 14.590000 164.050000 ;
        RECT  0.500000 164.050000 14.520000 164.120000 ;
        RECT  0.500000 164.120000 14.450000 164.190000 ;
        RECT  0.500000 164.190000 14.380000 164.260000 ;
        RECT  0.500000 164.260000 14.310000 164.330000 ;
        RECT  0.500000 164.330000 14.240000 164.400000 ;
        RECT  0.500000 164.400000 14.170000 164.470000 ;
        RECT  0.500000 164.470000 14.100000 164.540000 ;
        RECT  0.500000 164.540000 14.030000 164.610000 ;
        RECT  0.500000 164.610000 13.960000 164.680000 ;
        RECT  0.500000 164.680000 13.960000 169.940000 ;
        RECT  0.500000 169.940000 13.960000 170.010000 ;
        RECT  0.500000 170.010000 14.030000 170.080000 ;
        RECT  0.500000 170.080000 14.100000 170.150000 ;
        RECT  0.500000 170.150000 14.170000 170.220000 ;
        RECT  0.500000 170.220000 14.240000 170.290000 ;
        RECT  0.500000 170.290000 14.310000 170.360000 ;
        RECT  0.500000 170.360000 14.380000 170.430000 ;
        RECT  0.500000 170.430000 14.450000 170.500000 ;
        RECT  0.500000 170.500000 14.520000 170.570000 ;
        RECT  0.500000 170.570000 14.590000 170.640000 ;
        RECT  0.500000 170.640000 14.660000 170.710000 ;
        RECT  0.500000 170.710000 14.730000 170.780000 ;
        RECT  0.500000 170.780000 14.800000 170.850000 ;
        RECT  0.500000 170.850000 14.870000 170.920000 ;
        RECT  0.500000 170.920000 14.940000 170.990000 ;
        RECT  0.500000 170.990000 68.010000 173.630000 ;
        RECT  0.500000 173.630000 14.940000 173.700000 ;
        RECT  0.500000 173.700000 14.870000 173.770000 ;
        RECT  0.500000 173.770000 14.800000 173.840000 ;
        RECT  0.500000 173.840000 14.730000 173.910000 ;
        RECT  0.500000 173.910000 14.660000 173.980000 ;
        RECT  0.500000 173.980000 14.590000 174.050000 ;
        RECT  0.500000 174.050000 14.520000 174.120000 ;
        RECT  0.500000 174.120000 14.450000 174.190000 ;
        RECT  0.500000 174.190000 14.380000 174.260000 ;
        RECT  0.500000 174.260000 14.310000 174.330000 ;
        RECT  0.500000 174.330000 14.240000 174.400000 ;
        RECT  0.500000 174.400000 14.170000 174.470000 ;
        RECT  0.500000 174.470000 14.100000 174.540000 ;
        RECT  0.500000 174.540000 14.030000 174.610000 ;
        RECT  0.500000 174.610000 13.960000 174.680000 ;
        RECT  0.500000 174.680000 13.960000 179.940000 ;
        RECT  0.500000 179.940000 13.960000 180.010000 ;
        RECT  0.500000 180.010000 14.030000 180.080000 ;
        RECT  0.500000 180.080000 14.100000 180.150000 ;
        RECT  0.500000 180.150000 14.170000 180.220000 ;
        RECT  0.500000 180.220000 14.240000 180.290000 ;
        RECT  0.500000 180.290000 14.310000 180.360000 ;
        RECT  0.500000 180.360000 14.380000 180.430000 ;
        RECT  0.500000 180.430000 14.450000 180.500000 ;
        RECT  0.500000 180.500000 14.520000 180.570000 ;
        RECT  0.500000 180.570000 14.590000 180.640000 ;
        RECT  0.500000 180.640000 14.660000 180.710000 ;
        RECT  0.500000 180.710000 14.730000 180.780000 ;
        RECT  0.500000 180.780000 14.800000 180.850000 ;
        RECT  0.500000 180.850000 14.870000 180.920000 ;
        RECT  0.500000 180.920000 14.940000 180.990000 ;
        RECT  0.500000 180.990000 68.010000 183.630000 ;
        RECT  0.500000 183.630000 14.940000 183.700000 ;
        RECT  0.500000 183.700000 14.870000 183.770000 ;
        RECT  0.500000 183.770000 14.800000 183.840000 ;
        RECT  0.500000 183.840000 14.730000 183.910000 ;
        RECT  0.500000 183.910000 14.660000 183.980000 ;
        RECT  0.500000 183.980000 14.590000 184.050000 ;
        RECT  0.500000 184.050000 14.520000 184.120000 ;
        RECT  0.500000 184.120000 14.450000 184.190000 ;
        RECT  0.500000 184.190000 14.380000 184.260000 ;
        RECT  0.500000 184.260000 14.310000 184.330000 ;
        RECT  0.500000 184.330000 14.240000 184.400000 ;
        RECT  0.500000 184.400000 14.170000 184.470000 ;
        RECT  0.500000 184.470000 14.100000 184.540000 ;
        RECT  0.500000 184.540000 14.030000 184.610000 ;
        RECT  0.500000 184.610000 13.960000 184.680000 ;
        RECT  0.500000 184.680000 13.960000 189.940000 ;
        RECT  0.500000 189.940000 13.960000 190.010000 ;
        RECT  0.500000 190.010000 14.030000 190.080000 ;
        RECT  0.500000 190.080000 14.100000 190.150000 ;
        RECT  0.500000 190.150000 14.170000 190.220000 ;
        RECT  0.500000 190.220000 14.240000 190.290000 ;
        RECT  0.500000 190.290000 14.310000 190.360000 ;
        RECT  0.500000 190.360000 14.380000 190.430000 ;
        RECT  0.500000 190.430000 14.450000 190.500000 ;
        RECT  0.500000 190.500000 14.520000 190.570000 ;
        RECT  0.500000 190.570000 14.590000 190.640000 ;
        RECT  0.500000 190.640000 14.660000 190.710000 ;
        RECT  0.500000 190.710000 14.730000 190.780000 ;
        RECT  0.500000 190.780000 14.800000 190.850000 ;
        RECT  0.500000 190.850000 14.870000 190.920000 ;
        RECT  0.500000 190.920000 14.940000 190.990000 ;
        RECT  0.500000 190.990000 68.010000 193.630000 ;
        RECT 11.635000  10.210000 55.595000  10.215000 ;
        RECT 11.695000   7.655000 16.860000   7.725000 ;
        RECT 11.700000  10.145000 55.595000  10.210000 ;
        RECT 11.765000   7.725000 16.860000   7.795000 ;
        RECT 11.765000  10.080000 55.595000  10.145000 ;
        RECT 11.805000  10.040000 17.535000  10.080000 ;
        RECT 11.835000   7.795000 16.860000   7.865000 ;
        RECT 11.875000   9.970000 17.465000  10.040000 ;
        RECT 11.905000   7.865000 16.860000   7.935000 ;
        RECT 11.945000   9.900000 17.395000   9.970000 ;
        RECT 11.975000   7.935000 16.860000   8.005000 ;
        RECT 12.015000   8.005000 16.860000   8.045000 ;
        RECT 12.015000   8.045000 16.860000   9.365000 ;
        RECT 12.015000   9.365000 16.860000   9.435000 ;
        RECT 12.015000   9.435000 16.930000   9.505000 ;
        RECT 12.015000   9.505000 17.000000   9.575000 ;
        RECT 12.015000   9.575000 17.070000   9.645000 ;
        RECT 12.015000   9.645000 17.140000   9.715000 ;
        RECT 12.015000   9.715000 17.210000   9.785000 ;
        RECT 12.015000   9.785000 17.280000   9.830000 ;
        RECT 12.015000   9.830000 17.325000   9.900000 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 16.135000 31.010000 74.700000 33.650000 ;
        RECT 16.135000 40.990000 74.700000 43.630000 ;
        RECT 16.135000 51.010000 74.700000 53.650000 ;
        RECT 16.135000 60.990000 74.700000 63.630000 ;
        RECT 16.135000 70.990000 74.700000 73.630000 ;
        RECT 54.095000  0.000000 74.700000  7.815000 ;
        RECT 54.095000 19.990000 74.700000 21.695000 ;
        RECT 54.150000 19.935000 74.700000 19.990000 ;
        RECT 54.165000  7.815000 74.700000  7.885000 ;
        RECT 54.220000 19.865000 74.700000 19.935000 ;
        RECT 54.235000  7.885000 74.700000  7.955000 ;
        RECT 54.290000 19.795000 74.700000 19.865000 ;
        RECT 54.305000  7.955000 74.700000  8.025000 ;
        RECT 54.360000 19.725000 74.700000 19.795000 ;
        RECT 54.375000  8.025000 74.700000  8.095000 ;
        RECT 54.430000 19.655000 74.700000 19.725000 ;
        RECT 54.445000  8.095000 74.700000  8.165000 ;
        RECT 54.500000 19.585000 74.700000 19.655000 ;
        RECT 54.515000  8.165000 74.700000  8.235000 ;
        RECT 54.570000 19.515000 74.700000 19.585000 ;
        RECT 54.585000  8.235000 74.700000  8.305000 ;
        RECT 54.640000 19.445000 74.700000 19.515000 ;
        RECT 54.655000  8.305000 74.700000  8.375000 ;
        RECT 54.710000 19.375000 74.700000 19.445000 ;
        RECT 54.725000  8.375000 74.700000  8.445000 ;
        RECT 54.780000 19.305000 74.700000 19.375000 ;
        RECT 54.795000  8.445000 74.700000  8.515000 ;
        RECT 54.850000 19.235000 74.700000 19.305000 ;
        RECT 54.865000  8.515000 74.700000  8.585000 ;
        RECT 54.920000 19.165000 74.700000 19.235000 ;
        RECT 54.935000  8.585000 74.700000  8.655000 ;
        RECT 54.990000 19.095000 74.700000 19.165000 ;
        RECT 55.005000  8.655000 74.700000  8.725000 ;
        RECT 55.060000 19.025000 74.700000 19.095000 ;
        RECT 55.075000  8.725000 74.700000  8.795000 ;
        RECT 55.130000 18.955000 74.700000 19.025000 ;
        RECT 55.145000  8.795000 74.700000  8.865000 ;
        RECT 55.200000 18.885000 74.700000 18.955000 ;
        RECT 55.215000  8.865000 74.700000  8.935000 ;
        RECT 55.270000 18.815000 74.700000 18.885000 ;
        RECT 55.285000  8.935000 74.700000  9.005000 ;
        RECT 55.340000 18.745000 74.700000 18.815000 ;
        RECT 55.355000  9.005000 74.700000  9.075000 ;
        RECT 55.410000 18.675000 74.700000 18.745000 ;
        RECT 55.425000  9.075000 74.700000  9.145000 ;
        RECT 55.480000 18.605000 74.700000 18.675000 ;
        RECT 55.495000  9.145000 74.700000  9.215000 ;
        RECT 55.550000 18.535000 74.700000 18.605000 ;
        RECT 55.565000  9.215000 74.700000  9.285000 ;
        RECT 55.620000 18.465000 74.700000 18.535000 ;
        RECT 55.635000  9.285000 74.700000  9.355000 ;
        RECT 55.690000 18.395000 74.700000 18.465000 ;
        RECT 55.705000  9.355000 74.700000  9.425000 ;
        RECT 55.760000 18.325000 74.700000 18.395000 ;
        RECT 55.775000  9.425000 74.700000  9.495000 ;
        RECT 55.830000 18.255000 74.700000 18.325000 ;
        RECT 55.845000  9.495000 74.700000  9.565000 ;
        RECT 55.900000 18.185000 74.700000 18.255000 ;
        RECT 55.915000  9.565000 74.700000  9.635000 ;
        RECT 55.970000 18.115000 74.700000 18.185000 ;
        RECT 55.985000  9.635000 74.700000  9.705000 ;
        RECT 56.040000 18.045000 74.700000 18.115000 ;
        RECT 56.055000  9.705000 74.700000  9.775000 ;
        RECT 56.110000 17.975000 74.700000 18.045000 ;
        RECT 56.125000  9.775000 74.700000  9.845000 ;
        RECT 56.180000 17.905000 74.700000 17.975000 ;
        RECT 56.195000  9.845000 74.700000  9.915000 ;
        RECT 56.250000  9.915000 74.700000  9.970000 ;
        RECT 56.250000  9.970000 74.700000 17.835000 ;
        RECT 56.250000 17.835000 74.700000 17.905000 ;
        RECT 62.325000 21.695000 74.700000 21.765000 ;
        RECT 62.395000 21.765000 74.700000 21.835000 ;
        RECT 62.465000 21.835000 74.700000 21.905000 ;
        RECT 62.535000 21.905000 74.700000 21.975000 ;
        RECT 62.605000 21.975000 74.700000 22.045000 ;
        RECT 62.675000 22.045000 74.700000 22.115000 ;
        RECT 62.745000 22.115000 74.700000 22.185000 ;
        RECT 62.815000 22.185000 74.700000 22.255000 ;
        RECT 62.885000 22.255000 74.700000 22.325000 ;
        RECT 62.955000 22.325000 74.700000 22.395000 ;
        RECT 63.025000 22.395000 74.700000 22.465000 ;
        RECT 63.095000 22.465000 74.700000 22.535000 ;
        RECT 63.165000 22.535000 74.700000 22.605000 ;
        RECT 63.235000 22.605000 74.700000 22.675000 ;
        RECT 63.305000 22.675000 74.700000 22.745000 ;
        RECT 63.375000 22.745000 74.700000 22.815000 ;
        RECT 63.445000 22.815000 74.700000 22.885000 ;
        RECT 63.515000 22.885000 74.700000 22.955000 ;
        RECT 63.585000 22.955000 74.700000 23.025000 ;
        RECT 63.655000 23.025000 74.700000 23.095000 ;
        RECT 63.725000 23.095000 74.700000 23.165000 ;
        RECT 63.795000 23.165000 74.700000 23.235000 ;
        RECT 63.865000 23.235000 74.700000 23.305000 ;
        RECT 63.935000 23.305000 74.700000 23.375000 ;
        RECT 64.005000 23.375000 74.700000 23.445000 ;
        RECT 64.075000 23.445000 74.700000 23.515000 ;
        RECT 64.145000 23.515000 74.700000 23.585000 ;
        RECT 64.215000 23.585000 74.700000 23.655000 ;
        RECT 64.285000 23.655000 74.700000 23.725000 ;
        RECT 64.355000 23.725000 74.700000 23.795000 ;
        RECT 64.425000 23.795000 74.700000 23.865000 ;
        RECT 64.495000 23.865000 74.700000 23.935000 ;
        RECT 64.565000 23.935000 74.700000 24.005000 ;
        RECT 64.635000 24.005000 74.700000 24.075000 ;
        RECT 64.705000 24.075000 74.700000 24.145000 ;
        RECT 64.775000 24.145000 74.700000 24.215000 ;
        RECT 64.845000 24.215000 74.700000 24.285000 ;
        RECT 64.880000 31.000000 74.700000 31.010000 ;
        RECT 64.915000 24.285000 74.700000 24.355000 ;
        RECT 64.950000 30.930000 74.700000 31.000000 ;
        RECT 64.950000 40.985000 74.700000 40.990000 ;
        RECT 64.950000 51.005000 74.700000 51.010000 ;
        RECT 64.985000 24.355000 74.700000 24.425000 ;
        RECT 65.015000 60.920000 74.700000 60.990000 ;
        RECT 65.015000 63.630000 74.700000 63.700000 ;
        RECT 65.015000 70.920000 74.700000 70.990000 ;
        RECT 65.020000 30.860000 74.700000 30.930000 ;
        RECT 65.020000 40.915000 74.700000 40.985000 ;
        RECT 65.020000 50.935000 74.700000 51.005000 ;
        RECT 65.030000 33.650000 74.700000 33.720000 ;
        RECT 65.030000 43.630000 74.700000 43.700000 ;
        RECT 65.030000 53.650000 74.700000 53.720000 ;
        RECT 65.055000 24.425000 74.700000 24.495000 ;
        RECT 65.085000 60.850000 74.700000 60.920000 ;
        RECT 65.085000 63.700000 74.700000 63.770000 ;
        RECT 65.085000 70.850000 74.700000 70.920000 ;
        RECT 65.090000 30.790000 74.700000 30.860000 ;
        RECT 65.090000 40.845000 74.700000 40.915000 ;
        RECT 65.090000 50.865000 74.700000 50.935000 ;
        RECT 65.100000 33.720000 74.700000 33.790000 ;
        RECT 65.100000 43.700000 74.700000 43.770000 ;
        RECT 65.100000 53.720000 74.700000 53.790000 ;
        RECT 65.125000 24.495000 74.700000 24.565000 ;
        RECT 65.155000 60.780000 74.700000 60.850000 ;
        RECT 65.155000 63.770000 74.700000 63.840000 ;
        RECT 65.155000 70.780000 74.700000 70.850000 ;
        RECT 65.160000 30.720000 74.700000 30.790000 ;
        RECT 65.160000 40.775000 74.700000 40.845000 ;
        RECT 65.160000 50.795000 74.700000 50.865000 ;
        RECT 65.170000 33.790000 74.700000 33.860000 ;
        RECT 65.170000 43.770000 74.700000 43.840000 ;
        RECT 65.170000 53.790000 74.700000 53.860000 ;
        RECT 65.195000 24.565000 74.700000 24.635000 ;
        RECT 65.225000 60.710000 74.700000 60.780000 ;
        RECT 65.225000 63.840000 74.700000 63.910000 ;
        RECT 65.225000 70.710000 74.700000 70.780000 ;
        RECT 65.230000 30.650000 74.700000 30.720000 ;
        RECT 65.230000 40.705000 74.700000 40.775000 ;
        RECT 65.230000 50.725000 74.700000 50.795000 ;
        RECT 65.240000 33.860000 74.700000 33.930000 ;
        RECT 65.240000 43.840000 74.700000 43.910000 ;
        RECT 65.240000 53.860000 74.700000 53.930000 ;
        RECT 65.265000 24.635000 74.700000 24.705000 ;
        RECT 65.270000 73.630000 68.740000 73.700000 ;
        RECT 65.295000 60.640000 74.700000 60.710000 ;
        RECT 65.295000 63.910000 74.700000 63.980000 ;
        RECT 65.295000 70.640000 74.700000 70.710000 ;
        RECT 65.300000 30.580000 74.700000 30.650000 ;
        RECT 65.300000 40.635000 74.700000 40.705000 ;
        RECT 65.300000 50.655000 74.700000 50.725000 ;
        RECT 65.310000 33.930000 74.700000 34.000000 ;
        RECT 65.310000 43.910000 74.700000 43.980000 ;
        RECT 65.310000 53.930000 74.700000 54.000000 ;
        RECT 65.335000 24.705000 74.700000 24.775000 ;
        RECT 65.340000 73.700000 68.670000 73.770000 ;
        RECT 65.365000 60.570000 74.700000 60.640000 ;
        RECT 65.365000 63.980000 74.700000 64.050000 ;
        RECT 65.365000 70.570000 74.700000 70.640000 ;
        RECT 65.370000 30.510000 74.700000 30.580000 ;
        RECT 65.370000 40.565000 74.700000 40.635000 ;
        RECT 65.370000 50.585000 74.700000 50.655000 ;
        RECT 65.380000 34.000000 74.700000 34.070000 ;
        RECT 65.380000 43.980000 74.700000 44.050000 ;
        RECT 65.380000 54.000000 74.700000 54.070000 ;
        RECT 65.405000 24.775000 74.700000 24.845000 ;
        RECT 65.410000 73.770000 68.600000 73.840000 ;
        RECT 65.435000 60.500000 74.700000 60.570000 ;
        RECT 65.435000 64.050000 74.700000 64.120000 ;
        RECT 65.435000 70.500000 74.700000 70.570000 ;
        RECT 65.440000 30.440000 74.700000 30.510000 ;
        RECT 65.440000 40.495000 74.700000 40.565000 ;
        RECT 65.440000 50.515000 74.700000 50.585000 ;
        RECT 65.450000 34.070000 74.700000 34.140000 ;
        RECT 65.450000 44.050000 74.700000 44.120000 ;
        RECT 65.450000 54.070000 74.700000 54.140000 ;
        RECT 65.475000 24.845000 74.700000 24.915000 ;
        RECT 65.480000 73.840000 68.530000 73.910000 ;
        RECT 65.505000 60.430000 74.700000 60.500000 ;
        RECT 65.505000 64.120000 74.700000 64.190000 ;
        RECT 65.505000 70.430000 74.700000 70.500000 ;
        RECT 65.510000 30.370000 74.700000 30.440000 ;
        RECT 65.510000 40.425000 74.700000 40.495000 ;
        RECT 65.510000 50.445000 74.700000 50.515000 ;
        RECT 65.520000 34.140000 74.700000 34.210000 ;
        RECT 65.520000 44.120000 74.700000 44.190000 ;
        RECT 65.520000 54.140000 74.700000 54.210000 ;
        RECT 65.545000 24.915000 74.700000 24.985000 ;
        RECT 65.550000 73.910000 68.460000 73.980000 ;
        RECT 65.575000 60.360000 74.700000 60.430000 ;
        RECT 65.575000 64.190000 74.700000 64.260000 ;
        RECT 65.575000 70.360000 74.700000 70.430000 ;
        RECT 65.580000 30.300000 74.700000 30.370000 ;
        RECT 65.580000 40.355000 74.700000 40.425000 ;
        RECT 65.580000 50.375000 74.700000 50.445000 ;
        RECT 65.590000 34.210000 74.700000 34.280000 ;
        RECT 65.590000 44.190000 74.700000 44.260000 ;
        RECT 65.590000 54.210000 74.700000 54.280000 ;
        RECT 65.615000 24.985000 74.700000 25.055000 ;
        RECT 65.620000 73.980000 68.390000 74.050000 ;
        RECT 65.645000 60.290000 74.700000 60.360000 ;
        RECT 65.645000 64.260000 74.700000 64.330000 ;
        RECT 65.645000 70.290000 74.700000 70.360000 ;
        RECT 65.650000 30.230000 74.700000 30.300000 ;
        RECT 65.650000 40.285000 74.700000 40.355000 ;
        RECT 65.650000 50.305000 74.700000 50.375000 ;
        RECT 65.660000 34.280000 74.700000 34.350000 ;
        RECT 65.660000 44.260000 74.700000 44.330000 ;
        RECT 65.660000 54.280000 74.700000 54.350000 ;
        RECT 65.685000 25.055000 74.700000 25.125000 ;
        RECT 65.690000 74.050000 68.320000 74.120000 ;
        RECT 65.715000 60.220000 74.700000 60.290000 ;
        RECT 65.715000 64.330000 74.700000 64.400000 ;
        RECT 65.715000 70.220000 74.700000 70.290000 ;
        RECT 65.720000 30.160000 74.700000 30.230000 ;
        RECT 65.720000 40.215000 74.700000 40.285000 ;
        RECT 65.720000 50.235000 74.700000 50.305000 ;
        RECT 65.730000 34.350000 74.700000 34.420000 ;
        RECT 65.730000 44.330000 74.700000 44.400000 ;
        RECT 65.730000 54.350000 74.700000 54.420000 ;
        RECT 65.755000 25.125000 74.700000 25.195000 ;
        RECT 65.760000 74.120000 68.250000 74.190000 ;
        RECT 65.785000 60.150000 74.700000 60.220000 ;
        RECT 65.785000 64.400000 74.700000 64.470000 ;
        RECT 65.785000 70.150000 74.700000 70.220000 ;
        RECT 65.790000 30.090000 74.700000 30.160000 ;
        RECT 65.790000 40.145000 74.700000 40.215000 ;
        RECT 65.790000 50.165000 74.700000 50.235000 ;
        RECT 65.800000 34.420000 74.700000 34.490000 ;
        RECT 65.800000 44.400000 74.700000 44.470000 ;
        RECT 65.800000 54.420000 74.700000 54.490000 ;
        RECT 65.825000 25.195000 74.700000 25.265000 ;
        RECT 65.830000 74.190000 68.180000 74.260000 ;
        RECT 65.855000 60.080000 74.700000 60.150000 ;
        RECT 65.855000 64.470000 74.700000 64.540000 ;
        RECT 65.855000 70.080000 74.700000 70.150000 ;
        RECT 65.860000 30.020000 74.700000 30.090000 ;
        RECT 65.860000 40.075000 74.700000 40.145000 ;
        RECT 65.860000 50.095000 74.700000 50.165000 ;
        RECT 65.870000 34.490000 74.700000 34.560000 ;
        RECT 65.870000 44.470000 74.700000 44.540000 ;
        RECT 65.870000 54.490000 74.700000 54.560000 ;
        RECT 65.895000 25.265000 74.700000 25.335000 ;
        RECT 65.900000 74.260000 68.110000 74.330000 ;
        RECT 65.925000 60.010000 74.700000 60.080000 ;
        RECT 65.925000 64.540000 74.700000 64.610000 ;
        RECT 65.925000 70.010000 74.700000 70.080000 ;
        RECT 65.930000 29.950000 74.700000 30.020000 ;
        RECT 65.930000 40.005000 74.700000 40.075000 ;
        RECT 65.930000 50.025000 74.700000 50.095000 ;
        RECT 65.940000 34.560000 74.700000 34.630000 ;
        RECT 65.940000 44.540000 74.700000 44.610000 ;
        RECT 65.940000 54.560000 74.700000 54.630000 ;
        RECT 65.965000 25.335000 74.700000 25.405000 ;
        RECT 65.970000 74.330000 68.040000 74.400000 ;
        RECT 65.995000 54.630000 74.700000 54.685000 ;
        RECT 65.995000 54.685000 74.700000 59.940000 ;
        RECT 65.995000 59.940000 74.700000 60.010000 ;
        RECT 65.995000 64.610000 74.700000 64.680000 ;
        RECT 65.995000 64.680000 74.700000 69.940000 ;
        RECT 65.995000 69.940000 74.700000 70.010000 ;
        RECT 66.000000 25.405000 74.700000 25.440000 ;
        RECT 66.000000 25.440000 74.700000 29.880000 ;
        RECT 66.000000 29.880000 74.700000 29.950000 ;
        RECT 66.000000 34.630000 74.700000 34.690000 ;
        RECT 66.000000 34.690000 74.700000 39.935000 ;
        RECT 66.000000 39.935000 74.700000 40.005000 ;
        RECT 66.000000 44.610000 74.700000 44.670000 ;
        RECT 66.000000 44.670000 74.700000 49.955000 ;
        RECT 66.000000 49.955000 74.700000 50.025000 ;
        RECT 66.000000 74.400000 68.010000 74.430000 ;
        RECT 66.000000 74.430000 68.010000 98.560000 ;
    END
  END SRC_BDY_LVC2
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  0.240000  17.210000  2.995000  19.200000 ;
      RECT  1.350000   1.020000  7.110000   1.190000 ;
      RECT  1.350000   1.190000  1.520000  17.040000 ;
      RECT  1.350000  17.040000  7.110000  17.210000 ;
      RECT  1.760000  19.630000  9.385000  20.140000 ;
      RECT  1.760000  20.140000  2.685000  23.060000 ;
      RECT  1.845000   3.220000  2.015000   8.960000 ;
      RECT  1.845000   9.710000  2.015000  16.610000 ;
      RECT  2.070000   1.610000  6.390000   1.780000 ;
      RECT  2.070000   9.260000  6.390000   9.430000 ;
      RECT  2.305000   2.490000  2.475000   8.960000 ;
      RECT  2.305000  10.140000  2.475000  15.440000 ;
      RECT  2.765000   3.220000  2.935000   8.960000 ;
      RECT  2.765000   9.710000  2.935000  16.610000 ;
      RECT  3.225000   2.490000  3.395000   8.960000 ;
      RECT  3.225000  10.140000  3.395000  15.440000 ;
      RECT  3.685000   3.220000  3.855000   8.960000 ;
      RECT  3.685000   9.710000  3.855000  16.610000 ;
      RECT  4.145000   2.490000  4.315000   8.960000 ;
      RECT  4.145000  10.140000  4.315000  15.440000 ;
      RECT  4.605000   3.220000  4.775000   8.960000 ;
      RECT  4.605000   9.710000  4.775000  16.610000 ;
      RECT  4.975000  22.290000 10.650000  23.010000 ;
      RECT  5.065000   2.490000  5.235000   8.960000 ;
      RECT  5.065000  10.140000  5.235000  15.440000 ;
      RECT  5.525000   3.220000  5.695000   8.960000 ;
      RECT  5.525000   9.710000  5.695000  16.610000 ;
      RECT  5.890000  23.010000 10.650000  23.015000 ;
      RECT  5.985000   2.490000  6.155000   8.960000 ;
      RECT  5.985000  10.140000  6.155000  15.440000 ;
      RECT  6.445000   2.060000  6.615000   8.960000 ;
      RECT  6.445000   9.710000  6.615000  16.610000 ;
      RECT  6.940000   1.190000  7.110000  17.040000 ;
      RECT  8.340000 196.360000  8.670000 196.420000 ;
      RECT  8.345000   1.410000 16.655000  18.350000 ;
      RECT  8.420000 195.890000  8.590000 196.360000 ;
      RECT  9.155000 106.965000 10.280000 196.850000 ;
      RECT  9.155000 196.850000 69.720000 197.380000 ;
      RECT  9.185000  23.825000 69.720000  24.355000 ;
      RECT  9.185000  24.355000 10.280000  82.980000 ;
      RECT  9.185000  82.980000 21.740000  83.150000 ;
      RECT  9.185000  83.150000 10.280000  99.490000 ;
      RECT  9.730000  99.490000 10.280000 106.965000 ;
      RECT 10.920000  83.820000 11.830000  84.585000 ;
      RECT 11.065000 168.280000 12.220000 194.935000 ;
      RECT 11.065000 194.935000 68.495000 195.885000 ;
      RECT 11.095000 144.465000 21.490000 145.315000 ;
      RECT 11.095000 145.315000 12.220000 168.280000 ;
      RECT 11.275000  25.065000 68.140000  26.015000 ;
      RECT 11.275000  26.015000 12.220000  34.040000 ;
      RECT 11.275000  36.745000 12.220000  43.620000 ;
      RECT 11.275000  46.905000 12.220000  81.575000 ;
      RECT 11.275000  81.575000 23.280000  82.085000 ;
      RECT 11.370000  34.040000 12.220000  36.745000 ;
      RECT 11.370000  43.620000 12.220000  46.905000 ;
      RECT 12.405000 184.140000 66.575000 186.620000 ;
      RECT 12.430000 184.100000 66.575000 184.140000 ;
      RECT 12.750000  75.785000 12.920000  80.300000 ;
      RECT 12.975000  81.045000 66.655000  81.215000 ;
      RECT 13.060000  44.100000 65.590000  46.620000 ;
      RECT 13.060000  64.100000 65.590000  66.620000 ;
      RECT 13.190000  34.100000 65.590000  36.620000 ;
      RECT 13.190000  54.100000 65.590000  56.620000 ;
      RECT 13.335000 174.100000 65.590000 176.620000 ;
      RECT 13.365000 145.615000 14.305000 145.620000 ;
      RECT 13.365000 145.620000 65.590000 146.620000 ;
      RECT 13.365000 154.100000 65.590000 156.620000 ;
      RECT 13.365000 164.100000 65.590000 166.620000 ;
      RECT 13.395000  26.900000 13.925000  33.570000 ;
      RECT 13.395000  36.900000 13.925000  43.570000 ;
      RECT 13.395000  46.900000 13.925000  53.570000 ;
      RECT 13.395000  56.900000 13.925000  63.570000 ;
      RECT 13.395000  66.900000 13.925000  71.725000 ;
      RECT 13.395000 186.900000 13.925000 193.570000 ;
      RECT 14.360000 194.100000 65.590000 194.270000 ;
      RECT 14.780000  26.900000 15.310000  33.570000 ;
      RECT 14.780000  36.900000 15.310000  43.570000 ;
      RECT 14.780000  46.900000 15.310000  53.570000 ;
      RECT 14.780000  56.900000 15.310000  63.570000 ;
      RECT 14.780000  66.900000 15.310000  71.725000 ;
      RECT 14.780000 186.900000 15.310000 193.570000 ;
      RECT 14.790000  26.840000 15.300000  26.900000 ;
      RECT 14.790000  33.570000 15.300000  33.630000 ;
      RECT 14.790000  36.840000 15.300000  36.900000 ;
      RECT 14.790000  43.570000 15.300000  43.630000 ;
      RECT 14.790000  46.840000 15.300000  46.900000 ;
      RECT 14.790000  53.570000 15.300000  53.630000 ;
      RECT 14.790000  56.840000 15.300000  56.900000 ;
      RECT 14.790000  63.570000 15.300000  63.630000 ;
      RECT 14.790000  66.840000 15.300000  66.900000 ;
      RECT 14.790000 186.840000 15.300000 186.900000 ;
      RECT 14.790000 193.570000 15.300000 193.630000 ;
      RECT 15.865000 146.900000 16.395000 153.570000 ;
      RECT 15.865000 156.900000 16.395000 163.570000 ;
      RECT 15.865000 166.900000 16.395000 173.570000 ;
      RECT 16.165000  26.900000 16.695000  33.570000 ;
      RECT 16.165000  36.900000 16.695000  43.570000 ;
      RECT 16.165000  46.900000 16.695000  53.570000 ;
      RECT 16.165000  56.900000 16.695000  63.570000 ;
      RECT 16.165000  66.900000 16.695000  71.725000 ;
      RECT 16.165000 176.900000 16.695000 183.570000 ;
      RECT 16.165000 186.900000 16.695000 193.570000 ;
      RECT 17.000000  17.580000 56.200000  18.350000 ;
      RECT 17.030000  75.785000 17.200000  80.300000 ;
      RECT 17.550000  26.900000 18.080000  33.570000 ;
      RECT 17.550000  36.900000 18.080000  43.570000 ;
      RECT 17.550000  46.900000 18.080000  53.570000 ;
      RECT 17.550000  56.900000 18.080000  63.570000 ;
      RECT 17.550000  66.900000 18.080000  71.725000 ;
      RECT 17.550000 176.900000 18.080000 183.570000 ;
      RECT 17.550000 186.900000 18.080000 193.570000 ;
      RECT 17.560000  26.840000 18.070000  26.900000 ;
      RECT 17.560000  33.570000 18.070000  33.630000 ;
      RECT 17.560000  36.840000 18.070000  36.900000 ;
      RECT 17.560000  43.570000 18.070000  43.630000 ;
      RECT 17.560000  46.840000 18.070000  46.900000 ;
      RECT 17.560000  53.570000 18.070000  53.630000 ;
      RECT 17.560000  56.840000 18.070000  56.900000 ;
      RECT 17.560000  63.570000 18.070000  63.630000 ;
      RECT 17.560000  66.840000 18.070000  66.900000 ;
      RECT 17.560000 176.840000 18.070000 176.900000 ;
      RECT 17.560000 183.570000 18.070000 183.630000 ;
      RECT 17.560000 186.840000 18.070000 186.900000 ;
      RECT 17.560000 193.570000 18.070000 193.630000 ;
      RECT 17.955000 146.900000 18.485000 153.570000 ;
      RECT 17.955000 156.900000 18.485000 163.570000 ;
      RECT 17.955000 166.900000 18.485000 173.570000 ;
      RECT 17.965000 146.840000 18.475000 146.900000 ;
      RECT 17.965000 153.570000 18.475000 153.630000 ;
      RECT 17.965000 156.840000 18.475000 156.900000 ;
      RECT 17.965000 163.570000 18.475000 163.630000 ;
      RECT 17.965000 166.840000 18.475000 166.900000 ;
      RECT 17.965000 173.570000 18.475000 173.630000 ;
      RECT 18.935000  26.900000 19.465000  33.570000 ;
      RECT 18.935000  36.900000 19.465000  43.570000 ;
      RECT 18.935000  46.900000 19.465000  53.570000 ;
      RECT 18.935000  56.900000 19.465000  63.570000 ;
      RECT 18.935000  66.900000 19.465000  71.725000 ;
      RECT 18.935000 176.900000 19.465000 183.570000 ;
      RECT 18.935000 186.900000 19.465000 193.570000 ;
      RECT 19.495000  83.820000 20.405000  84.585000 ;
      RECT 20.045000 146.900000 20.575000 153.570000 ;
      RECT 20.045000 156.900000 20.575000 163.570000 ;
      RECT 20.045000 166.900000 20.575000 173.570000 ;
      RECT 20.320000  26.900000 20.850000  33.570000 ;
      RECT 20.320000  36.900000 20.850000  43.570000 ;
      RECT 20.320000  46.900000 20.850000  53.570000 ;
      RECT 20.320000  56.900000 20.850000  63.570000 ;
      RECT 20.320000  66.900000 20.850000  71.725000 ;
      RECT 20.320000 176.900000 20.850000 183.570000 ;
      RECT 20.320000 186.900000 20.850000 193.570000 ;
      RECT 20.330000  26.840000 20.840000  26.900000 ;
      RECT 20.330000  33.570000 20.840000  33.630000 ;
      RECT 20.330000  36.840000 20.840000  36.900000 ;
      RECT 20.330000  43.570000 20.840000  43.630000 ;
      RECT 20.330000  46.840000 20.840000  46.900000 ;
      RECT 20.330000  53.570000 20.840000  53.630000 ;
      RECT 20.330000  56.840000 20.840000  56.900000 ;
      RECT 20.330000  63.570000 20.840000  63.630000 ;
      RECT 20.330000  66.840000 20.840000  66.900000 ;
      RECT 20.330000 176.840000 20.840000 176.900000 ;
      RECT 20.330000 183.570000 20.840000 183.630000 ;
      RECT 20.330000 186.840000 20.840000 186.900000 ;
      RECT 20.330000 193.570000 20.840000 193.630000 ;
      RECT 20.640000 100.865000 68.495000 101.035000 ;
      RECT 20.640000 101.035000 21.490000 109.275000 ;
      RECT 20.640000 109.275000 68.495000 109.445000 ;
      RECT 20.640000 109.445000 21.490000 117.770000 ;
      RECT 20.640000 117.770000 68.495000 117.940000 ;
      RECT 20.640000 117.940000 21.490000 144.465000 ;
      RECT 21.570000  83.150000 21.740000  99.925000 ;
      RECT 21.570000  99.925000 69.720000 100.095000 ;
      RECT 21.660000 128.010000 65.590000 128.515000 ;
      RECT 21.690000 134.100000 65.590000 136.620000 ;
      RECT 21.705000  26.900000 22.235000  33.570000 ;
      RECT 21.705000  36.900000 22.235000  43.570000 ;
      RECT 21.705000  46.900000 22.235000  53.570000 ;
      RECT 21.705000  56.900000 22.235000  63.570000 ;
      RECT 21.705000  66.900000 22.235000  71.725000 ;
      RECT 21.705000 176.900000 22.235000 183.570000 ;
      RECT 21.705000 186.900000 22.235000 193.570000 ;
      RECT 22.135000 146.900000 22.665000 153.570000 ;
      RECT 22.135000 156.900000 22.665000 163.570000 ;
      RECT 22.135000 166.900000 22.665000 173.570000 ;
      RECT 22.145000 146.840000 22.655000 146.900000 ;
      RECT 22.145000 153.570000 22.655000 153.630000 ;
      RECT 22.145000 156.840000 22.655000 156.900000 ;
      RECT 22.145000 163.570000 22.655000 163.630000 ;
      RECT 22.145000 166.840000 22.655000 166.900000 ;
      RECT 22.145000 173.570000 22.655000 173.630000 ;
      RECT 22.430000  82.085000 23.280000  82.180000 ;
      RECT 22.430000  82.180000 68.140000  82.350000 ;
      RECT 22.430000  82.350000 23.280000  90.675000 ;
      RECT 22.430000  90.675000 68.140000  90.845000 ;
      RECT 22.430000  90.845000 23.280000  97.890000 ;
      RECT 22.770000  97.890000 23.280000  98.990000 ;
      RECT 22.770000  98.990000 68.140000  99.160000 ;
      RECT 23.090000  26.900000 23.620000  33.570000 ;
      RECT 23.090000  36.900000 23.620000  43.570000 ;
      RECT 23.090000  46.900000 23.620000  53.570000 ;
      RECT 23.090000  56.900000 23.620000  63.570000 ;
      RECT 23.090000  66.900000 23.620000  71.725000 ;
      RECT 23.090000 176.900000 23.620000 183.570000 ;
      RECT 23.090000 186.900000 23.620000 193.570000 ;
      RECT 23.100000  26.840000 23.610000  26.900000 ;
      RECT 23.100000  33.570000 23.610000  33.630000 ;
      RECT 23.100000  36.840000 23.610000  36.900000 ;
      RECT 23.100000  43.570000 23.610000  43.630000 ;
      RECT 23.100000  46.840000 23.610000  46.900000 ;
      RECT 23.100000  53.570000 23.610000  53.630000 ;
      RECT 23.100000  56.840000 23.610000  56.900000 ;
      RECT 23.100000  63.570000 23.610000  63.630000 ;
      RECT 23.100000  66.840000 23.610000  66.900000 ;
      RECT 23.100000 176.840000 23.610000 176.900000 ;
      RECT 23.100000 183.570000 23.610000 183.630000 ;
      RECT 23.100000 186.840000 23.610000 186.900000 ;
      RECT 23.100000 193.570000 23.610000 193.630000 ;
      RECT 23.405000 144.100000 65.590000 145.620000 ;
      RECT 23.635000 101.385000 24.045000 108.175000 ;
      RECT 23.635000 109.880000 24.045000 115.550000 ;
      RECT 23.635000 120.080000 24.045000 125.295000 ;
      RECT 23.685000  82.785000 24.215000  89.575000 ;
      RECT 23.685000  91.280000 24.215000  98.070000 ;
      RECT 23.805000 115.550000 24.045000 116.670000 ;
      RECT 23.805000 118.955000 24.045000 120.080000 ;
      RECT 23.805000 125.295000 24.045000 125.745000 ;
      RECT 24.225000 128.730000 24.755000 133.760000 ;
      RECT 24.225000 136.900000 24.755000 143.570000 ;
      RECT 24.225000 146.900000 24.755000 153.570000 ;
      RECT 24.225000 156.900000 24.755000 163.570000 ;
      RECT 24.225000 166.900000 24.755000 173.570000 ;
      RECT 24.475000  26.900000 25.005000  33.570000 ;
      RECT 24.475000  36.900000 25.005000  43.570000 ;
      RECT 24.475000  46.900000 25.005000  53.570000 ;
      RECT 24.475000  56.900000 25.005000  63.570000 ;
      RECT 24.475000  66.900000 25.005000  71.725000 ;
      RECT 24.475000 176.900000 25.005000 183.570000 ;
      RECT 24.475000 186.900000 25.005000 193.570000 ;
      RECT 24.615000  90.045000 66.655000  90.215000 ;
      RECT 24.615000  98.540000 66.655000  98.710000 ;
      RECT 24.670000 108.645000 66.655000 108.815000 ;
      RECT 24.670000 117.140000 66.655000 117.310000 ;
      RECT 24.670000 118.315000 66.655000 118.485000 ;
      RECT 25.310000  75.785000 25.480000  80.300000 ;
      RECT 25.310000  82.915000 25.480000  89.020000 ;
      RECT 25.310000  91.930000 25.480000  96.925000 ;
      RECT 25.365000 101.385000 25.535000 106.255000 ;
      RECT 25.365000 110.450000 25.535000 115.330000 ;
      RECT 25.365000 120.080000 25.535000 124.860000 ;
      RECT 25.860000  26.900000 26.390000  33.570000 ;
      RECT 25.860000  36.900000 26.390000  43.570000 ;
      RECT 25.860000  46.900000 26.390000  53.570000 ;
      RECT 25.860000  56.900000 26.390000  63.570000 ;
      RECT 25.860000  66.900000 26.390000  71.725000 ;
      RECT 25.860000 176.900000 26.390000 183.570000 ;
      RECT 25.860000 186.900000 26.390000 193.570000 ;
      RECT 25.870000  26.840000 26.380000  26.900000 ;
      RECT 25.870000  33.570000 26.380000  33.630000 ;
      RECT 25.870000  36.840000 26.380000  36.900000 ;
      RECT 25.870000  43.570000 26.380000  43.630000 ;
      RECT 25.870000  46.840000 26.380000  46.900000 ;
      RECT 25.870000  53.570000 26.380000  53.630000 ;
      RECT 25.870000  56.840000 26.380000  56.900000 ;
      RECT 25.870000  63.570000 26.380000  63.630000 ;
      RECT 25.870000  66.840000 26.380000  66.900000 ;
      RECT 25.870000 176.840000 26.380000 176.900000 ;
      RECT 25.870000 183.570000 26.380000 183.630000 ;
      RECT 25.870000 186.840000 26.380000 186.900000 ;
      RECT 25.870000 193.570000 26.380000 193.630000 ;
      RECT 26.315000 128.730000 26.845000 133.715000 ;
      RECT 26.315000 136.900000 26.845000 143.570000 ;
      RECT 26.315000 146.900000 26.845000 153.570000 ;
      RECT 26.315000 156.900000 26.845000 163.570000 ;
      RECT 26.315000 166.900000 26.845000 173.570000 ;
      RECT 26.325000 136.840000 26.835000 136.900000 ;
      RECT 26.325000 143.570000 26.835000 143.630000 ;
      RECT 26.325000 146.840000 26.835000 146.900000 ;
      RECT 26.325000 153.570000 26.835000 153.630000 ;
      RECT 26.325000 156.840000 26.835000 156.900000 ;
      RECT 26.325000 163.570000 26.835000 163.630000 ;
      RECT 26.325000 166.840000 26.835000 166.900000 ;
      RECT 26.325000 173.570000 26.835000 173.630000 ;
      RECT 27.245000  26.900000 27.775000  33.570000 ;
      RECT 27.245000  36.900000 27.775000  43.570000 ;
      RECT 27.245000  46.900000 27.775000  53.570000 ;
      RECT 27.245000  56.900000 27.775000  63.570000 ;
      RECT 27.245000  66.900000 27.775000  71.725000 ;
      RECT 27.245000 176.900000 27.775000 183.570000 ;
      RECT 27.245000 186.900000 27.775000 193.570000 ;
      RECT 28.405000 128.860000 28.935000 133.760000 ;
      RECT 28.405000 136.900000 28.935000 143.570000 ;
      RECT 28.405000 146.900000 28.935000 153.570000 ;
      RECT 28.405000 156.900000 28.935000 163.570000 ;
      RECT 28.405000 166.900000 28.935000 173.570000 ;
      RECT 28.630000  26.900000 29.160000  33.570000 ;
      RECT 28.630000  36.900000 29.160000  43.570000 ;
      RECT 28.630000  46.900000 29.160000  53.570000 ;
      RECT 28.630000  56.900000 29.160000  63.570000 ;
      RECT 28.630000  66.900000 29.160000  71.725000 ;
      RECT 28.630000 176.900000 29.160000 183.570000 ;
      RECT 28.630000 186.900000 29.160000 193.570000 ;
      RECT 28.640000  26.840000 29.150000  26.900000 ;
      RECT 28.640000  33.570000 29.150000  33.630000 ;
      RECT 28.640000  36.840000 29.150000  36.900000 ;
      RECT 28.640000  43.570000 29.150000  43.630000 ;
      RECT 28.640000  46.840000 29.150000  46.900000 ;
      RECT 28.640000  53.570000 29.150000  53.630000 ;
      RECT 28.640000  56.840000 29.150000  56.900000 ;
      RECT 28.640000  63.570000 29.150000  63.630000 ;
      RECT 28.640000  66.840000 29.150000  66.900000 ;
      RECT 28.640000 176.840000 29.150000 176.900000 ;
      RECT 28.640000 183.570000 29.150000 183.630000 ;
      RECT 28.640000 186.840000 29.150000 186.900000 ;
      RECT 28.640000 193.570000 29.150000 193.630000 ;
      RECT 30.015000  26.900000 30.545000  33.570000 ;
      RECT 30.015000  36.900000 30.545000  43.570000 ;
      RECT 30.015000  46.900000 30.545000  53.570000 ;
      RECT 30.015000  56.900000 30.545000  63.570000 ;
      RECT 30.015000  66.900000 30.545000  71.725000 ;
      RECT 30.015000 176.900000 30.545000 183.570000 ;
      RECT 30.015000 186.900000 30.545000 193.570000 ;
      RECT 30.495000 128.730000 31.025000 133.715000 ;
      RECT 30.495000 136.900000 31.025000 143.570000 ;
      RECT 30.495000 146.900000 31.025000 153.570000 ;
      RECT 30.495000 156.900000 31.025000 163.570000 ;
      RECT 30.495000 166.900000 31.025000 173.570000 ;
      RECT 30.505000 136.840000 31.015000 136.900000 ;
      RECT 30.505000 143.570000 31.015000 143.630000 ;
      RECT 30.505000 146.840000 31.015000 146.900000 ;
      RECT 30.505000 153.570000 31.015000 153.630000 ;
      RECT 30.505000 156.840000 31.015000 156.900000 ;
      RECT 30.505000 163.570000 31.015000 163.630000 ;
      RECT 30.505000 166.840000 31.015000 166.900000 ;
      RECT 30.505000 173.570000 31.015000 173.630000 ;
      RECT 31.400000  26.900000 31.930000  33.570000 ;
      RECT 31.400000  36.900000 31.930000  43.570000 ;
      RECT 31.400000  46.900000 31.930000  53.570000 ;
      RECT 31.400000  56.900000 31.930000  63.570000 ;
      RECT 31.400000  66.900000 31.930000  71.725000 ;
      RECT 31.400000 176.900000 31.930000 183.570000 ;
      RECT 31.400000 186.900000 31.930000 193.570000 ;
      RECT 31.410000  26.840000 31.920000  26.900000 ;
      RECT 31.410000  33.570000 31.920000  33.630000 ;
      RECT 31.410000  36.840000 31.920000  36.900000 ;
      RECT 31.410000  43.570000 31.920000  43.630000 ;
      RECT 31.410000  46.840000 31.920000  46.900000 ;
      RECT 31.410000  53.570000 31.920000  53.630000 ;
      RECT 31.410000  56.840000 31.920000  56.900000 ;
      RECT 31.410000  63.570000 31.920000  63.630000 ;
      RECT 31.410000  66.840000 31.920000  66.900000 ;
      RECT 31.410000 176.840000 31.920000 176.900000 ;
      RECT 31.410000 183.570000 31.920000 183.630000 ;
      RECT 31.410000 186.840000 31.920000 186.900000 ;
      RECT 31.410000 193.570000 31.920000 193.630000 ;
      RECT 32.585000 128.730000 33.115000 133.755000 ;
      RECT 32.585000 136.900000 33.115000 143.570000 ;
      RECT 32.585000 146.900000 33.115000 153.570000 ;
      RECT 32.585000 156.900000 33.115000 163.570000 ;
      RECT 32.585000 166.900000 33.115000 173.570000 ;
      RECT 32.785000  26.900000 33.315000  33.570000 ;
      RECT 32.785000  36.900000 33.315000  43.570000 ;
      RECT 32.785000  46.900000 33.315000  53.570000 ;
      RECT 32.785000  56.900000 33.315000  63.570000 ;
      RECT 32.785000  66.900000 33.315000  71.725000 ;
      RECT 32.785000 176.900000 33.315000 183.570000 ;
      RECT 32.785000 186.900000 33.315000 193.570000 ;
      RECT 33.590000  75.785000 33.760000  80.300000 ;
      RECT 33.590000  82.915000 33.760000  89.020000 ;
      RECT 33.590000  91.930000 33.760000  96.925000 ;
      RECT 33.590000 101.385000 33.760000 106.255000 ;
      RECT 33.590000 110.450000 33.760000 115.270000 ;
      RECT 33.595000 120.080000 33.765000 124.860000 ;
      RECT 34.170000  26.900000 34.700000  33.570000 ;
      RECT 34.170000  36.900000 34.700000  43.570000 ;
      RECT 34.170000  46.900000 34.700000  53.570000 ;
      RECT 34.170000  56.900000 34.700000  63.570000 ;
      RECT 34.170000  66.900000 34.700000  71.725000 ;
      RECT 34.170000 176.900000 34.700000 183.570000 ;
      RECT 34.170000 186.900000 34.700000 193.570000 ;
      RECT 34.180000  26.840000 34.690000  26.900000 ;
      RECT 34.180000  33.570000 34.690000  33.630000 ;
      RECT 34.180000  36.840000 34.690000  36.900000 ;
      RECT 34.180000  43.570000 34.690000  43.630000 ;
      RECT 34.180000  46.840000 34.690000  46.900000 ;
      RECT 34.180000  53.570000 34.690000  53.630000 ;
      RECT 34.180000  56.840000 34.690000  56.900000 ;
      RECT 34.180000  63.570000 34.690000  63.630000 ;
      RECT 34.180000  66.840000 34.690000  66.900000 ;
      RECT 34.180000 176.840000 34.690000 176.900000 ;
      RECT 34.180000 183.570000 34.690000 183.630000 ;
      RECT 34.180000 186.840000 34.690000 186.900000 ;
      RECT 34.180000 193.570000 34.690000 193.630000 ;
      RECT 34.675000 128.730000 35.205000 133.840000 ;
      RECT 34.675000 136.900000 35.205000 143.570000 ;
      RECT 34.675000 146.900000 35.205000 153.570000 ;
      RECT 34.675000 156.900000 35.205000 163.570000 ;
      RECT 34.675000 166.900000 35.205000 173.570000 ;
      RECT 34.685000 136.840000 35.195000 136.900000 ;
      RECT 34.685000 143.570000 35.195000 143.630000 ;
      RECT 34.685000 146.840000 35.195000 146.900000 ;
      RECT 34.685000 153.570000 35.195000 153.630000 ;
      RECT 34.685000 156.840000 35.195000 156.900000 ;
      RECT 34.685000 163.570000 35.195000 163.630000 ;
      RECT 34.685000 166.840000 35.195000 166.900000 ;
      RECT 34.685000 173.570000 35.195000 173.630000 ;
      RECT 35.555000  26.900000 36.085000  33.570000 ;
      RECT 35.555000  36.900000 36.085000  43.570000 ;
      RECT 35.555000  46.900000 36.085000  53.570000 ;
      RECT 35.555000  56.900000 36.085000  63.570000 ;
      RECT 35.555000  66.900000 36.085000  71.725000 ;
      RECT 35.555000 176.900000 36.085000 183.570000 ;
      RECT 35.555000 186.900000 36.085000 193.570000 ;
      RECT 36.765000 128.730000 37.295000 133.755000 ;
      RECT 36.765000 136.900000 37.295000 143.570000 ;
      RECT 36.765000 146.900000 37.295000 153.570000 ;
      RECT 36.765000 156.900000 37.295000 163.570000 ;
      RECT 36.765000 166.900000 37.295000 173.570000 ;
      RECT 36.940000  26.900000 37.470000  33.570000 ;
      RECT 36.940000  36.900000 37.470000  43.570000 ;
      RECT 36.940000  46.900000 37.470000  53.570000 ;
      RECT 36.940000  56.900000 37.470000  63.570000 ;
      RECT 36.940000  66.900000 37.470000  71.725000 ;
      RECT 36.940000 176.900000 37.470000 183.570000 ;
      RECT 36.940000 186.900000 37.470000 193.570000 ;
      RECT 36.950000  26.840000 37.460000  26.900000 ;
      RECT 36.950000  33.570000 37.460000  33.630000 ;
      RECT 36.950000  36.840000 37.460000  36.900000 ;
      RECT 36.950000  43.570000 37.460000  43.630000 ;
      RECT 36.950000  46.840000 37.460000  46.900000 ;
      RECT 36.950000  53.570000 37.460000  53.630000 ;
      RECT 36.950000  56.840000 37.460000  56.900000 ;
      RECT 36.950000  63.570000 37.460000  63.630000 ;
      RECT 36.950000  66.840000 37.460000  66.900000 ;
      RECT 36.950000 176.840000 37.460000 176.900000 ;
      RECT 36.950000 183.570000 37.460000 183.630000 ;
      RECT 36.950000 186.840000 37.460000 186.900000 ;
      RECT 36.950000 193.570000 37.460000 193.630000 ;
      RECT 38.325000  26.900000 38.855000  33.570000 ;
      RECT 38.325000  36.900000 38.855000  43.570000 ;
      RECT 38.325000  46.900000 38.855000  53.570000 ;
      RECT 38.325000  56.900000 38.855000  63.570000 ;
      RECT 38.325000  66.900000 38.855000  71.725000 ;
      RECT 38.325000 176.900000 38.855000 183.570000 ;
      RECT 38.325000 186.900000 38.855000 193.570000 ;
      RECT 38.855000 128.730000 39.385000 133.925000 ;
      RECT 38.855000 136.900000 39.385000 143.570000 ;
      RECT 38.855000 146.900000 39.385000 153.570000 ;
      RECT 38.855000 156.900000 39.385000 163.570000 ;
      RECT 38.855000 166.900000 39.385000 173.570000 ;
      RECT 38.865000 136.840000 39.375000 136.900000 ;
      RECT 38.865000 143.570000 39.375000 143.630000 ;
      RECT 38.865000 146.840000 39.375000 146.900000 ;
      RECT 38.865000 153.570000 39.375000 153.630000 ;
      RECT 38.865000 156.840000 39.375000 156.900000 ;
      RECT 38.865000 163.570000 39.375000 163.630000 ;
      RECT 38.865000 166.840000 39.375000 166.900000 ;
      RECT 38.865000 173.570000 39.375000 173.630000 ;
      RECT 39.710000  26.900000 40.240000  33.570000 ;
      RECT 39.710000  36.900000 40.240000  43.570000 ;
      RECT 39.710000  46.900000 40.240000  53.570000 ;
      RECT 39.710000  56.900000 40.240000  63.570000 ;
      RECT 39.710000  66.900000 40.240000  71.725000 ;
      RECT 39.710000 176.900000 40.240000 183.570000 ;
      RECT 39.710000 186.900000 40.240000 193.570000 ;
      RECT 39.720000  26.840000 40.230000  26.900000 ;
      RECT 39.720000  33.570000 40.230000  33.630000 ;
      RECT 39.720000  36.840000 40.230000  36.900000 ;
      RECT 39.720000  43.570000 40.230000  43.630000 ;
      RECT 39.720000  46.840000 40.230000  46.900000 ;
      RECT 39.720000  53.570000 40.230000  53.630000 ;
      RECT 39.720000  56.840000 40.230000  56.900000 ;
      RECT 39.720000  63.570000 40.230000  63.630000 ;
      RECT 39.720000  66.840000 40.230000  66.900000 ;
      RECT 39.720000 176.840000 40.230000 176.900000 ;
      RECT 39.720000 183.570000 40.230000 183.630000 ;
      RECT 39.720000 186.840000 40.230000 186.900000 ;
      RECT 39.720000 193.570000 40.230000 193.630000 ;
      RECT 40.945000 128.730000 41.475000 133.755000 ;
      RECT 40.945000 136.900000 41.475000 143.570000 ;
      RECT 40.945000 146.900000 41.475000 153.570000 ;
      RECT 40.945000 156.900000 41.475000 163.570000 ;
      RECT 40.945000 166.900000 41.475000 173.570000 ;
      RECT 41.095000  26.900000 41.625000  33.570000 ;
      RECT 41.095000  36.900000 41.625000  43.570000 ;
      RECT 41.095000  46.900000 41.625000  53.570000 ;
      RECT 41.095000  56.900000 41.625000  63.570000 ;
      RECT 41.095000  66.900000 41.625000  71.725000 ;
      RECT 41.095000 176.900000 41.625000 183.570000 ;
      RECT 41.095000 186.900000 41.625000 193.570000 ;
      RECT 41.870000  75.785000 42.040000  80.300000 ;
      RECT 41.870000  82.915000 42.040000  89.020000 ;
      RECT 41.870000  91.930000 42.040000  96.925000 ;
      RECT 41.870000 101.385000 42.040000 106.255000 ;
      RECT 41.870000 110.450000 42.040000 115.270000 ;
      RECT 41.870000 120.080000 42.040000 124.860000 ;
      RECT 42.480000  26.900000 43.010000  33.570000 ;
      RECT 42.480000  36.900000 43.010000  43.570000 ;
      RECT 42.480000  46.900000 43.010000  53.570000 ;
      RECT 42.480000  56.900000 43.010000  63.570000 ;
      RECT 42.480000  66.900000 43.010000  71.725000 ;
      RECT 42.480000 176.900000 43.010000 183.570000 ;
      RECT 42.480000 186.900000 43.010000 193.570000 ;
      RECT 42.490000  26.840000 43.000000  26.900000 ;
      RECT 42.490000  33.570000 43.000000  33.630000 ;
      RECT 42.490000  36.840000 43.000000  36.900000 ;
      RECT 42.490000  43.570000 43.000000  43.630000 ;
      RECT 42.490000  46.840000 43.000000  46.900000 ;
      RECT 42.490000  53.570000 43.000000  53.630000 ;
      RECT 42.490000  56.840000 43.000000  56.900000 ;
      RECT 42.490000  63.570000 43.000000  63.630000 ;
      RECT 42.490000  66.840000 43.000000  66.900000 ;
      RECT 42.490000 176.840000 43.000000 176.900000 ;
      RECT 42.490000 183.570000 43.000000 183.630000 ;
      RECT 42.490000 186.840000 43.000000 186.900000 ;
      RECT 42.490000 193.570000 43.000000 193.630000 ;
      RECT 43.035000 128.730000 43.565000 133.925000 ;
      RECT 43.035000 136.900000 43.565000 143.570000 ;
      RECT 43.035000 146.900000 43.565000 153.570000 ;
      RECT 43.035000 156.900000 43.565000 163.570000 ;
      RECT 43.035000 166.900000 43.565000 173.570000 ;
      RECT 43.045000 136.840000 43.555000 136.900000 ;
      RECT 43.045000 143.570000 43.555000 143.630000 ;
      RECT 43.045000 146.840000 43.555000 146.900000 ;
      RECT 43.045000 153.570000 43.555000 153.630000 ;
      RECT 43.045000 156.840000 43.555000 156.900000 ;
      RECT 43.045000 163.570000 43.555000 163.630000 ;
      RECT 43.045000 166.840000 43.555000 166.900000 ;
      RECT 43.045000 173.570000 43.555000 173.630000 ;
      RECT 43.865000  26.900000 44.395000  33.570000 ;
      RECT 43.865000  36.900000 44.395000  43.570000 ;
      RECT 43.865000  46.900000 44.395000  53.570000 ;
      RECT 43.865000  56.900000 44.395000  63.570000 ;
      RECT 43.865000  66.900000 44.395000  71.725000 ;
      RECT 43.865000 176.900000 44.395000 183.570000 ;
      RECT 43.865000 186.900000 44.395000 193.570000 ;
      RECT 45.125000 128.730000 45.655000 133.755000 ;
      RECT 45.125000 136.900000 45.655000 143.570000 ;
      RECT 45.125000 146.900000 45.655000 153.570000 ;
      RECT 45.125000 156.900000 45.655000 163.570000 ;
      RECT 45.125000 166.900000 45.655000 173.570000 ;
      RECT 45.250000  26.900000 45.780000  33.570000 ;
      RECT 45.250000  36.900000 45.780000  43.570000 ;
      RECT 45.250000  46.900000 45.780000  53.570000 ;
      RECT 45.250000  56.900000 45.780000  63.570000 ;
      RECT 45.250000  66.900000 45.780000  71.725000 ;
      RECT 45.250000 176.900000 45.780000 183.570000 ;
      RECT 45.250000 186.900000 45.780000 193.570000 ;
      RECT 45.260000  26.840000 45.770000  26.900000 ;
      RECT 45.260000  33.570000 45.770000  33.630000 ;
      RECT 45.260000  36.840000 45.770000  36.900000 ;
      RECT 45.260000  43.570000 45.770000  43.630000 ;
      RECT 45.260000  46.840000 45.770000  46.900000 ;
      RECT 45.260000  53.570000 45.770000  53.630000 ;
      RECT 45.260000  56.840000 45.770000  56.900000 ;
      RECT 45.260000  63.570000 45.770000  63.630000 ;
      RECT 45.260000  66.840000 45.770000  66.900000 ;
      RECT 45.260000 176.840000 45.770000 176.900000 ;
      RECT 45.260000 183.570000 45.770000 183.630000 ;
      RECT 45.260000 186.840000 45.770000 186.900000 ;
      RECT 45.260000 193.570000 45.770000 193.630000 ;
      RECT 46.635000  26.900000 47.165000  33.570000 ;
      RECT 46.635000  36.900000 47.165000  43.570000 ;
      RECT 46.635000  46.900000 47.165000  53.570000 ;
      RECT 46.635000  56.900000 47.165000  63.570000 ;
      RECT 46.635000  66.900000 47.165000  71.725000 ;
      RECT 46.635000 176.900000 47.165000 183.570000 ;
      RECT 46.635000 186.900000 47.165000 193.570000 ;
      RECT 47.215000 128.730000 47.745000 133.925000 ;
      RECT 47.215000 136.900000 47.745000 143.570000 ;
      RECT 47.215000 146.900000 47.745000 153.570000 ;
      RECT 47.215000 156.900000 47.745000 163.570000 ;
      RECT 47.215000 166.900000 47.745000 173.570000 ;
      RECT 47.225000 136.840000 47.735000 136.900000 ;
      RECT 47.225000 143.570000 47.735000 143.630000 ;
      RECT 47.225000 146.840000 47.735000 146.900000 ;
      RECT 47.225000 153.570000 47.735000 153.630000 ;
      RECT 47.225000 156.840000 47.735000 156.900000 ;
      RECT 47.225000 163.570000 47.735000 163.630000 ;
      RECT 47.225000 166.840000 47.735000 166.900000 ;
      RECT 47.225000 173.570000 47.735000 173.630000 ;
      RECT 48.020000  26.900000 48.550000  33.570000 ;
      RECT 48.020000  36.900000 48.550000  43.570000 ;
      RECT 48.020000  46.900000 48.550000  53.570000 ;
      RECT 48.020000  56.900000 48.550000  63.570000 ;
      RECT 48.020000  66.900000 48.550000  71.725000 ;
      RECT 48.020000 176.900000 48.550000 183.570000 ;
      RECT 48.020000 186.900000 48.550000 193.570000 ;
      RECT 48.030000  26.840000 48.540000  26.900000 ;
      RECT 48.030000  33.570000 48.540000  33.630000 ;
      RECT 48.030000  36.840000 48.540000  36.900000 ;
      RECT 48.030000  43.570000 48.540000  43.630000 ;
      RECT 48.030000  46.840000 48.540000  46.900000 ;
      RECT 48.030000  53.570000 48.540000  53.630000 ;
      RECT 48.030000  56.840000 48.540000  56.900000 ;
      RECT 48.030000  63.570000 48.540000  63.630000 ;
      RECT 48.030000  66.840000 48.540000  66.900000 ;
      RECT 48.030000 176.840000 48.540000 176.900000 ;
      RECT 48.030000 183.570000 48.540000 183.630000 ;
      RECT 48.030000 186.840000 48.540000 186.900000 ;
      RECT 48.030000 193.570000 48.540000 193.630000 ;
      RECT 49.305000 128.730000 49.835000 133.755000 ;
      RECT 49.305000 136.900000 49.835000 143.570000 ;
      RECT 49.305000 146.900000 49.835000 153.570000 ;
      RECT 49.305000 156.900000 49.835000 163.570000 ;
      RECT 49.305000 166.900000 49.835000 173.570000 ;
      RECT 49.405000  26.900000 49.935000  33.570000 ;
      RECT 49.405000  36.900000 49.935000  43.570000 ;
      RECT 49.405000  46.900000 49.935000  53.570000 ;
      RECT 49.405000  56.900000 49.935000  63.570000 ;
      RECT 49.405000  66.900000 49.935000  71.725000 ;
      RECT 49.405000 176.900000 49.935000 183.570000 ;
      RECT 49.405000 186.900000 49.935000 193.570000 ;
      RECT 50.150000  75.785000 50.320000  80.300000 ;
      RECT 50.150000  82.915000 50.320000  89.020000 ;
      RECT 50.150000  91.930000 50.320000  96.925000 ;
      RECT 50.150000 101.385000 50.320000 106.255000 ;
      RECT 50.150000 110.450000 50.320000 115.270000 ;
      RECT 50.150000 120.080000 50.320000 124.860000 ;
      RECT 50.790000  26.900000 51.320000  33.570000 ;
      RECT 50.790000  36.900000 51.320000  43.570000 ;
      RECT 50.790000  46.900000 51.320000  53.570000 ;
      RECT 50.790000  56.900000 51.320000  63.570000 ;
      RECT 50.790000  66.900000 51.320000  71.725000 ;
      RECT 50.790000 176.900000 51.320000 183.570000 ;
      RECT 50.790000 186.900000 51.320000 193.570000 ;
      RECT 50.800000  26.840000 51.310000  26.900000 ;
      RECT 50.800000  33.570000 51.310000  33.630000 ;
      RECT 50.800000  36.840000 51.310000  36.900000 ;
      RECT 50.800000  43.570000 51.310000  43.630000 ;
      RECT 50.800000  46.840000 51.310000  46.900000 ;
      RECT 50.800000  53.570000 51.310000  53.630000 ;
      RECT 50.800000  56.840000 51.310000  56.900000 ;
      RECT 50.800000  63.570000 51.310000  63.630000 ;
      RECT 50.800000  66.840000 51.310000  66.900000 ;
      RECT 50.800000 176.840000 51.310000 176.900000 ;
      RECT 50.800000 183.570000 51.310000 183.630000 ;
      RECT 50.800000 186.840000 51.310000 186.900000 ;
      RECT 50.800000 193.570000 51.310000 193.630000 ;
      RECT 51.395000 128.730000 51.925000 133.925000 ;
      RECT 51.395000 136.900000 51.925000 143.570000 ;
      RECT 51.395000 146.900000 51.925000 153.570000 ;
      RECT 51.395000 156.900000 51.925000 163.570000 ;
      RECT 51.395000 166.900000 51.925000 173.570000 ;
      RECT 51.405000 136.840000 51.915000 136.900000 ;
      RECT 51.405000 143.570000 51.915000 143.630000 ;
      RECT 51.405000 146.840000 51.915000 146.900000 ;
      RECT 51.405000 153.570000 51.915000 153.630000 ;
      RECT 51.405000 156.840000 51.915000 156.900000 ;
      RECT 51.405000 163.570000 51.915000 163.630000 ;
      RECT 51.405000 166.840000 51.915000 166.900000 ;
      RECT 51.405000 173.570000 51.915000 173.630000 ;
      RECT 52.175000  26.900000 52.705000  33.570000 ;
      RECT 52.175000  36.900000 52.705000  43.570000 ;
      RECT 52.175000  46.900000 52.705000  53.570000 ;
      RECT 52.175000  56.900000 52.705000  63.570000 ;
      RECT 52.175000  66.900000 52.705000  71.725000 ;
      RECT 52.175000 176.900000 52.705000 183.570000 ;
      RECT 52.175000 186.900000 52.705000 193.570000 ;
      RECT 53.485000 128.730000 54.015000 133.755000 ;
      RECT 53.485000 136.900000 54.015000 143.570000 ;
      RECT 53.485000 146.900000 54.015000 153.570000 ;
      RECT 53.485000 156.900000 54.015000 163.570000 ;
      RECT 53.485000 166.900000 54.015000 173.570000 ;
      RECT 53.560000  26.900000 54.090000  33.570000 ;
      RECT 53.560000  36.900000 54.090000  43.570000 ;
      RECT 53.560000  46.900000 54.090000  53.570000 ;
      RECT 53.560000  56.900000 54.090000  63.570000 ;
      RECT 53.560000  66.900000 54.090000  71.725000 ;
      RECT 53.560000 176.900000 54.090000 183.570000 ;
      RECT 53.560000 186.900000 54.090000 193.570000 ;
      RECT 53.570000  26.840000 54.080000  26.900000 ;
      RECT 53.570000  33.570000 54.080000  33.630000 ;
      RECT 53.570000  36.840000 54.080000  36.900000 ;
      RECT 53.570000  43.570000 54.080000  43.630000 ;
      RECT 53.570000  46.840000 54.080000  46.900000 ;
      RECT 53.570000  53.570000 54.080000  53.630000 ;
      RECT 53.570000  56.840000 54.080000  56.900000 ;
      RECT 53.570000  63.570000 54.080000  63.630000 ;
      RECT 53.570000  66.840000 54.080000  66.900000 ;
      RECT 53.570000 176.840000 54.080000 176.900000 ;
      RECT 53.570000 183.570000 54.080000 183.630000 ;
      RECT 53.570000 186.840000 54.080000 186.900000 ;
      RECT 53.570000 193.570000 54.080000 193.630000 ;
      RECT 54.945000  26.900000 55.475000  33.570000 ;
      RECT 54.945000  36.900000 55.475000  43.570000 ;
      RECT 54.945000  46.900000 55.475000  53.570000 ;
      RECT 54.945000  56.900000 55.475000  63.570000 ;
      RECT 54.945000  66.900000 55.475000  71.725000 ;
      RECT 54.945000 176.900000 55.475000 183.570000 ;
      RECT 54.945000 186.900000 55.475000 193.570000 ;
      RECT 55.575000 128.730000 56.105000 133.925000 ;
      RECT 55.575000 136.900000 56.105000 143.570000 ;
      RECT 55.575000 146.900000 56.105000 153.570000 ;
      RECT 55.575000 156.900000 56.105000 163.570000 ;
      RECT 55.575000 166.900000 56.105000 173.570000 ;
      RECT 55.585000 136.840000 56.095000 136.900000 ;
      RECT 55.585000 143.570000 56.095000 143.630000 ;
      RECT 55.585000 146.840000 56.095000 146.900000 ;
      RECT 55.585000 153.570000 56.095000 153.630000 ;
      RECT 55.585000 156.840000 56.095000 156.900000 ;
      RECT 55.585000 163.570000 56.095000 163.630000 ;
      RECT 55.585000 166.840000 56.095000 166.900000 ;
      RECT 55.585000 173.570000 56.095000 173.630000 ;
      RECT 56.330000  26.900000 56.860000  33.570000 ;
      RECT 56.330000  36.900000 56.860000  43.570000 ;
      RECT 56.330000  46.900000 56.860000  53.570000 ;
      RECT 56.330000  56.900000 56.860000  63.570000 ;
      RECT 56.330000  66.900000 56.860000  71.725000 ;
      RECT 56.330000 176.900000 56.860000 183.570000 ;
      RECT 56.330000 186.900000 56.860000 193.570000 ;
      RECT 56.340000  26.840000 56.850000  26.900000 ;
      RECT 56.340000  33.570000 56.850000  33.630000 ;
      RECT 56.340000  36.840000 56.850000  36.900000 ;
      RECT 56.340000  43.570000 56.850000  43.630000 ;
      RECT 56.340000  46.840000 56.850000  46.900000 ;
      RECT 56.340000  53.570000 56.850000  53.630000 ;
      RECT 56.340000  56.840000 56.850000  56.900000 ;
      RECT 56.340000  63.570000 56.850000  63.630000 ;
      RECT 56.340000  66.840000 56.850000  66.900000 ;
      RECT 56.340000 176.840000 56.850000 176.900000 ;
      RECT 56.340000 183.570000 56.850000 183.630000 ;
      RECT 56.340000 186.840000 56.850000 186.900000 ;
      RECT 56.340000 193.570000 56.850000 193.630000 ;
      RECT 56.980000  16.365000 57.510000  16.895000 ;
      RECT 57.665000 128.730000 58.195000 133.755000 ;
      RECT 57.665000 136.900000 58.195000 143.570000 ;
      RECT 57.665000 146.900000 58.195000 153.570000 ;
      RECT 57.665000 156.900000 58.195000 163.570000 ;
      RECT 57.665000 166.900000 58.195000 173.570000 ;
      RECT 57.715000  26.900000 58.245000  33.570000 ;
      RECT 57.715000  36.900000 58.245000  43.570000 ;
      RECT 57.715000  46.900000 58.245000  53.570000 ;
      RECT 57.715000  56.900000 58.245000  63.570000 ;
      RECT 57.715000  66.900000 58.245000  71.725000 ;
      RECT 57.715000 176.900000 58.245000 183.570000 ;
      RECT 57.715000 186.900000 58.245000 193.570000 ;
      RECT 58.430000  75.785000 58.600000  80.300000 ;
      RECT 58.430000  82.915000 58.600000  89.020000 ;
      RECT 58.430000  91.930000 58.600000  96.925000 ;
      RECT 58.430000 101.385000 58.600000 106.255000 ;
      RECT 58.430000 110.450000 58.600000 115.270000 ;
      RECT 58.430000 120.080000 58.600000 124.860000 ;
      RECT 59.100000  26.900000 59.630000  33.570000 ;
      RECT 59.100000  36.900000 59.630000  43.570000 ;
      RECT 59.100000  46.900000 59.630000  53.570000 ;
      RECT 59.100000  56.900000 59.630000  63.570000 ;
      RECT 59.100000  66.900000 59.630000  71.725000 ;
      RECT 59.100000 176.900000 59.630000 183.570000 ;
      RECT 59.100000 186.900000 59.630000 193.570000 ;
      RECT 59.110000  26.840000 59.620000  26.900000 ;
      RECT 59.110000  33.570000 59.620000  33.630000 ;
      RECT 59.110000  36.840000 59.620000  36.900000 ;
      RECT 59.110000  43.570000 59.620000  43.630000 ;
      RECT 59.110000  46.840000 59.620000  46.900000 ;
      RECT 59.110000  53.570000 59.620000  53.630000 ;
      RECT 59.110000  56.840000 59.620000  56.900000 ;
      RECT 59.110000  63.570000 59.620000  63.630000 ;
      RECT 59.110000  66.840000 59.620000  66.900000 ;
      RECT 59.110000 176.840000 59.620000 176.900000 ;
      RECT 59.110000 183.570000 59.620000 183.630000 ;
      RECT 59.110000 186.840000 59.620000 186.900000 ;
      RECT 59.110000 193.570000 59.620000 193.630000 ;
      RECT 59.755000 128.730000 60.285000 133.925000 ;
      RECT 59.755000 136.900000 60.285000 143.570000 ;
      RECT 59.755000 146.900000 60.285000 153.570000 ;
      RECT 59.755000 156.900000 60.285000 163.570000 ;
      RECT 59.755000 166.900000 60.285000 173.570000 ;
      RECT 59.765000 136.840000 60.275000 136.900000 ;
      RECT 59.765000 143.570000 60.275000 143.630000 ;
      RECT 59.765000 146.840000 60.275000 146.900000 ;
      RECT 59.765000 153.570000 60.275000 153.630000 ;
      RECT 59.765000 156.840000 60.275000 156.900000 ;
      RECT 59.765000 163.570000 60.275000 163.630000 ;
      RECT 59.765000 166.840000 60.275000 166.900000 ;
      RECT 59.765000 173.570000 60.275000 173.630000 ;
      RECT 60.485000  26.900000 61.015000  33.570000 ;
      RECT 60.485000  36.900000 61.015000  43.570000 ;
      RECT 60.485000  46.900000 61.015000  53.570000 ;
      RECT 60.485000  56.900000 61.015000  63.570000 ;
      RECT 60.485000  66.900000 61.015000  71.725000 ;
      RECT 60.485000 176.900000 61.015000 183.570000 ;
      RECT 60.485000 186.900000 61.015000 193.570000 ;
      RECT 61.845000 128.730000 62.375000 133.755000 ;
      RECT 61.845000 136.900000 62.375000 143.570000 ;
      RECT 61.845000 146.900000 62.375000 153.570000 ;
      RECT 61.845000 156.900000 62.375000 163.570000 ;
      RECT 61.845000 166.900000 62.375000 173.570000 ;
      RECT 61.870000  26.900000 62.400000  33.570000 ;
      RECT 61.870000  36.900000 62.400000  43.570000 ;
      RECT 61.870000  46.900000 62.400000  53.570000 ;
      RECT 61.870000  56.900000 62.400000  63.570000 ;
      RECT 61.870000  66.900000 62.400000  71.725000 ;
      RECT 61.870000 176.900000 62.400000 183.570000 ;
      RECT 61.870000 186.900000 62.400000 193.570000 ;
      RECT 61.880000  26.840000 62.390000  26.900000 ;
      RECT 61.880000  33.570000 62.390000  33.630000 ;
      RECT 61.880000  36.840000 62.390000  36.900000 ;
      RECT 61.880000  43.570000 62.390000  43.630000 ;
      RECT 61.880000  46.840000 62.390000  46.900000 ;
      RECT 61.880000  53.570000 62.390000  53.630000 ;
      RECT 61.880000  56.840000 62.390000  56.900000 ;
      RECT 61.880000  63.570000 62.390000  63.630000 ;
      RECT 61.880000  66.840000 62.390000  66.900000 ;
      RECT 61.880000 176.840000 62.390000 176.900000 ;
      RECT 61.880000 183.570000 62.390000 183.630000 ;
      RECT 61.880000 186.840000 62.390000 186.900000 ;
      RECT 61.880000 193.570000 62.390000 193.630000 ;
      RECT 63.255000  26.900000 63.785000  33.570000 ;
      RECT 63.255000  36.900000 63.785000  43.570000 ;
      RECT 63.255000  46.900000 63.785000  53.570000 ;
      RECT 63.255000  56.900000 63.785000  63.570000 ;
      RECT 63.255000  66.900000 63.785000  71.725000 ;
      RECT 63.255000 176.900000 63.785000 183.570000 ;
      RECT 63.255000 186.900000 63.785000 193.570000 ;
      RECT 63.935000 128.730000 64.465000 133.925000 ;
      RECT 63.935000 136.900000 64.465000 143.570000 ;
      RECT 63.935000 146.900000 64.465000 153.570000 ;
      RECT 63.935000 156.900000 64.465000 163.570000 ;
      RECT 63.935000 166.900000 64.465000 173.570000 ;
      RECT 63.945000 136.840000 64.455000 136.900000 ;
      RECT 63.945000 143.570000 64.455000 143.630000 ;
      RECT 63.945000 146.840000 64.455000 146.900000 ;
      RECT 63.945000 153.570000 64.455000 153.630000 ;
      RECT 63.945000 156.840000 64.455000 156.900000 ;
      RECT 63.945000 163.570000 64.455000 163.630000 ;
      RECT 63.945000 166.840000 64.455000 166.900000 ;
      RECT 63.945000 173.570000 64.455000 173.630000 ;
      RECT 64.640000  26.900000 65.170000  33.570000 ;
      RECT 64.640000  36.900000 65.170000  43.570000 ;
      RECT 64.640000  46.900000 65.170000  53.570000 ;
      RECT 64.640000  56.900000 65.170000  63.570000 ;
      RECT 64.640000  66.900000 65.170000  71.725000 ;
      RECT 64.640000 176.900000 65.170000 183.570000 ;
      RECT 64.640000 186.900000 65.170000 193.570000 ;
      RECT 64.650000  26.840000 65.160000  26.900000 ;
      RECT 64.650000  33.570000 65.160000  33.630000 ;
      RECT 64.650000  36.840000 65.160000  36.900000 ;
      RECT 64.650000  43.570000 65.160000  43.630000 ;
      RECT 64.650000  46.840000 65.160000  46.900000 ;
      RECT 64.650000  53.570000 65.160000  53.630000 ;
      RECT 64.650000  56.840000 65.160000  56.900000 ;
      RECT 64.650000  63.570000 65.160000  63.630000 ;
      RECT 64.650000  66.840000 65.160000  66.900000 ;
      RECT 64.650000 176.840000 65.160000 176.900000 ;
      RECT 64.650000 183.570000 65.160000 183.630000 ;
      RECT 64.650000 186.840000 65.160000 186.900000 ;
      RECT 64.650000 193.570000 65.160000 193.630000 ;
      RECT 66.025000  26.900000 66.555000  33.570000 ;
      RECT 66.025000  36.900000 66.555000  43.570000 ;
      RECT 66.025000  46.900000 66.555000  53.570000 ;
      RECT 66.025000  56.900000 66.555000  63.570000 ;
      RECT 66.025000  66.900000 66.555000  71.725000 ;
      RECT 66.025000 128.730000 66.555000 133.755000 ;
      RECT 66.025000 136.900000 66.555000 143.570000 ;
      RECT 66.025000 146.900000 66.555000 153.570000 ;
      RECT 66.025000 156.900000 66.555000 163.570000 ;
      RECT 66.025000 166.900000 66.555000 173.570000 ;
      RECT 66.025000 176.900000 66.555000 183.570000 ;
      RECT 66.025000 186.900000 66.555000 193.570000 ;
      RECT 66.700000   1.205000 67.230000   1.735000 ;
      RECT 66.710000  75.785000 66.880000  80.535000 ;
      RECT 66.710000  82.785000 66.880000  89.375000 ;
      RECT 66.710000  91.280000 66.880000  97.870000 ;
      RECT 66.710000 101.385000 66.880000 106.255000 ;
      RECT 66.710000 110.450000 66.880000 115.270000 ;
      RECT 66.710000 120.080000 66.880000 124.860000 ;
      RECT 67.290000  26.015000 68.140000  82.180000 ;
      RECT 67.290000  82.350000 68.140000  90.675000 ;
      RECT 67.290000  90.845000 68.140000  98.990000 ;
      RECT 67.575000 101.035000 68.495000 109.275000 ;
      RECT 67.575000 109.445000 68.495000 117.770000 ;
      RECT 67.575000 117.940000 68.495000 194.935000 ;
      RECT 67.610000   1.080000 73.375000   1.250000 ;
      RECT 67.615000   1.250000 67.785000  17.100000 ;
      RECT 67.615000  17.100000 73.375000  17.270000 ;
      RECT 68.110000   3.280000 68.280000   9.020000 ;
      RECT 68.110000   9.770000 68.280000  16.670000 ;
      RECT 68.335000   1.670000 72.655000   1.840000 ;
      RECT 68.335000   9.320000 72.655000   9.490000 ;
      RECT 68.570000   2.550000 68.740000   9.020000 ;
      RECT 68.570000  10.200000 68.740000  15.660000 ;
      RECT 69.030000   3.280000 69.200000   9.020000 ;
      RECT 69.030000   9.770000 69.200000  16.670000 ;
      RECT 69.190000  24.355000 69.720000  99.925000 ;
      RECT 69.190000 100.095000 69.720000 196.850000 ;
      RECT 69.490000   2.550000 69.660000   9.020000 ;
      RECT 69.490000  10.200000 69.660000  15.660000 ;
      RECT 69.530000  19.010000 70.265000  19.610000 ;
      RECT 69.950000   3.280000 70.120000   9.020000 ;
      RECT 69.950000   9.770000 70.120000  16.670000 ;
      RECT 70.410000   2.550000 70.580000   9.020000 ;
      RECT 70.410000  10.200000 70.580000  15.660000 ;
      RECT 70.495000  17.960000 71.095000  18.695000 ;
      RECT 70.870000   3.280000 71.040000   9.020000 ;
      RECT 70.870000   9.770000 71.040000  16.670000 ;
      RECT 71.330000   2.550000 71.500000   9.020000 ;
      RECT 71.330000  10.200000 71.500000  15.660000 ;
      RECT 71.790000   3.280000 71.960000   9.020000 ;
      RECT 71.790000   9.770000 71.960000  16.670000 ;
      RECT 72.250000   2.550000 72.420000   9.020000 ;
      RECT 72.250000  10.200000 72.420000  15.660000 ;
      RECT 72.710000   2.120000 72.880000   9.020000 ;
      RECT 72.710000   9.770000 72.880000  16.670000 ;
      RECT 73.205000   1.250000 73.375000  17.100000 ;
      RECT 73.875000 196.920000 74.755000 197.780000 ;
    LAYER met1 ;
      RECT  0.000000   0.000000 25.930000   0.295000 ;
      RECT  0.000000   0.000000 26.070000   0.310000 ;
      RECT  0.000000   0.295000 25.930000   0.310000 ;
      RECT  0.000000   0.310000 25.945000   0.325000 ;
      RECT  0.000000   0.310000 75.000000 198.000000 ;
      RECT  0.000000   0.325000 75.000000   3.330000 ;
      RECT  0.000000   3.330000  3.005000 194.995000 ;
      RECT  0.000000 194.995000 75.000000 198.000000 ;
      RECT  3.000000   3.002000 24.390000   3.070000 ;
      RECT  3.000000   3.002000 24.390000   3.070000 ;
      RECT  3.000000   3.070000 24.460000   3.140000 ;
      RECT  3.000000   3.070000 24.460000   3.140000 ;
      RECT  3.000000   3.140000 24.530000   3.210000 ;
      RECT  3.000000   3.140000 24.530000   3.210000 ;
      RECT  3.000000   3.210000 24.600000   3.280000 ;
      RECT  3.000000   3.210000 24.600000   3.280000 ;
      RECT  3.000000   3.280000 24.670000   3.325000 ;
      RECT  3.000000   3.280000 24.670000   3.325000 ;
      RECT  3.000000   3.325000 72.000000 195.000000 ;
      RECT 27.840000   0.000000 75.000000   0.310000 ;
      RECT 27.950000   0.320000 75.000000   0.325000 ;
      RECT 27.965000   0.305000 75.000000   0.320000 ;
      RECT 27.980000   0.000000 75.000000   0.290000 ;
      RECT 27.980000   0.290000 75.000000   0.305000 ;
      RECT 30.950000   3.000000 72.000000   6.330000 ;
      RECT 71.995000   3.330000 75.000000 194.995000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  0.220000 193.910000 ;
      RECT  0.000000   0.000000  0.220000 193.910000 ;
      RECT  0.000000 193.910000 75.000000 198.000000 ;
      RECT  0.000000 193.910000 75.000000 198.000000 ;
      RECT 10.700000   8.165000 11.735000   9.705000 ;
      RECT 10.700000   8.165000 11.735000   9.705000 ;
      RECT 10.700000   9.705000 11.735000   9.715000 ;
      RECT 10.705000   8.160000 11.735000   8.165000 ;
      RECT 10.705000   8.160000 11.735000   8.165000 ;
      RECT 10.705000   9.705000 11.735000   9.710000 ;
      RECT 10.710000   9.710000 11.735000   9.715000 ;
      RECT 10.710000   9.715000 11.515000   9.935000 ;
      RECT 10.720000   8.145000 11.720000   8.160000 ;
      RECT 10.780000   9.715000 11.665000   9.785000 ;
      RECT 10.790000   8.075000 11.650000   8.145000 ;
      RECT 10.850000   9.785000 11.595000   9.855000 ;
      RECT 10.860000   8.005000 11.580000   8.075000 ;
      RECT 10.920000   9.855000 11.525000   9.925000 ;
      RECT 10.930000   7.935000 11.510000   8.005000 ;
      RECT 10.930000   7.935000 11.735000   8.160000 ;
      RECT 10.930000   9.925000 11.515000   9.935000 ;
      RECT 14.030000  25.300000 65.465000  25.370000 ;
      RECT 14.030000  25.300000 65.465000  25.370000 ;
      RECT 14.030000  25.300000 65.860000  25.500000 ;
      RECT 14.030000  25.370000 65.535000  25.440000 ;
      RECT 14.030000  25.370000 65.535000  25.440000 ;
      RECT 14.030000  25.440000 65.605000  25.510000 ;
      RECT 14.030000  25.440000 65.605000  25.510000 ;
      RECT 14.030000  25.500000 65.860000  29.820000 ;
      RECT 14.030000  25.510000 65.675000  25.555000 ;
      RECT 14.030000  25.510000 65.675000  25.555000 ;
      RECT 14.030000  25.555000 65.720000  29.765000 ;
      RECT 14.030000  29.765000 65.650000  29.835000 ;
      RECT 14.030000  29.765000 65.650000  29.835000 ;
      RECT 14.030000  29.820000 64.810000  30.870000 ;
      RECT 14.030000  29.835000 65.580000  29.905000 ;
      RECT 14.030000  29.835000 65.580000  29.905000 ;
      RECT 14.030000  29.905000 65.510000  29.975000 ;
      RECT 14.030000  29.905000 65.510000  29.975000 ;
      RECT 14.030000  29.975000 65.440000  30.045000 ;
      RECT 14.030000  29.975000 65.440000  30.045000 ;
      RECT 14.030000  30.045000 65.370000  30.115000 ;
      RECT 14.030000  30.045000 65.370000  30.115000 ;
      RECT 14.030000  30.115000 65.300000  30.185000 ;
      RECT 14.030000  30.115000 65.300000  30.185000 ;
      RECT 14.030000  30.185000 65.230000  30.255000 ;
      RECT 14.030000  30.185000 65.230000  30.255000 ;
      RECT 14.030000  30.255000 65.160000  30.325000 ;
      RECT 14.030000  30.255000 65.160000  30.325000 ;
      RECT 14.030000  30.325000 65.090000  30.395000 ;
      RECT 14.030000  30.325000 65.090000  30.395000 ;
      RECT 14.030000  30.395000 65.020000  30.465000 ;
      RECT 14.030000  30.395000 65.020000  30.465000 ;
      RECT 14.030000  30.465000 64.950000  30.535000 ;
      RECT 14.030000  30.465000 64.950000  30.535000 ;
      RECT 14.030000  30.535000 64.880000  30.605000 ;
      RECT 14.030000  30.535000 64.880000  30.605000 ;
      RECT 14.030000  30.605000 64.810000  30.675000 ;
      RECT 14.030000  30.605000 64.810000  30.675000 ;
      RECT 14.030000  30.675000 64.755000  30.730000 ;
      RECT 14.030000  30.675000 64.755000  30.730000 ;
      RECT 14.030000  30.730000 15.855000  33.930000 ;
      RECT 14.030000  30.870000 15.995000  33.790000 ;
      RECT 14.030000  33.790000 65.860000  34.750000 ;
      RECT 14.030000  33.930000 64.845000  34.000000 ;
      RECT 14.030000  33.930000 64.845000  34.000000 ;
      RECT 14.030000  34.000000 64.915000  34.070000 ;
      RECT 14.030000  34.000000 64.915000  34.070000 ;
      RECT 14.030000  34.070000 64.985000  34.140000 ;
      RECT 14.030000  34.070000 64.985000  34.140000 ;
      RECT 14.030000  34.140000 65.055000  34.210000 ;
      RECT 14.030000  34.140000 65.055000  34.210000 ;
      RECT 14.030000  34.210000 65.125000  34.280000 ;
      RECT 14.030000  34.210000 65.125000  34.280000 ;
      RECT 14.030000  34.280000 65.195000  34.350000 ;
      RECT 14.030000  34.280000 65.195000  34.350000 ;
      RECT 14.030000  34.350000 65.265000  34.420000 ;
      RECT 14.030000  34.350000 65.265000  34.420000 ;
      RECT 14.030000  34.420000 65.335000  34.490000 ;
      RECT 14.030000  34.420000 65.335000  34.490000 ;
      RECT 14.030000  34.490000 65.405000  34.560000 ;
      RECT 14.030000  34.490000 65.405000  34.560000 ;
      RECT 14.030000  34.560000 65.475000  34.630000 ;
      RECT 14.030000  34.560000 65.475000  34.630000 ;
      RECT 14.030000  34.630000 65.545000  34.700000 ;
      RECT 14.030000  34.630000 65.545000  34.700000 ;
      RECT 14.030000  34.700000 65.615000  34.770000 ;
      RECT 14.030000  34.700000 65.615000  34.770000 ;
      RECT 14.030000  34.750000 65.860000  39.875000 ;
      RECT 14.030000  34.770000 65.685000  34.805000 ;
      RECT 14.030000  34.770000 65.685000  34.805000 ;
      RECT 14.030000  34.805000 65.720000  39.820000 ;
      RECT 14.030000  39.820000 65.650000  39.890000 ;
      RECT 14.030000  39.820000 65.650000  39.890000 ;
      RECT 14.030000  39.875000 64.885000  40.850000 ;
      RECT 14.030000  39.890000 65.580000  39.960000 ;
      RECT 14.030000  39.890000 65.580000  39.960000 ;
      RECT 14.030000  39.960000 65.510000  40.030000 ;
      RECT 14.030000  39.960000 65.510000  40.030000 ;
      RECT 14.030000  40.030000 65.440000  40.100000 ;
      RECT 14.030000  40.030000 65.440000  40.100000 ;
      RECT 14.030000  40.100000 65.370000  40.170000 ;
      RECT 14.030000  40.100000 65.370000  40.170000 ;
      RECT 14.030000  40.170000 65.300000  40.240000 ;
      RECT 14.030000  40.170000 65.300000  40.240000 ;
      RECT 14.030000  40.240000 65.230000  40.310000 ;
      RECT 14.030000  40.240000 65.230000  40.310000 ;
      RECT 14.030000  40.310000 65.160000  40.380000 ;
      RECT 14.030000  40.310000 65.160000  40.380000 ;
      RECT 14.030000  40.380000 65.090000  40.450000 ;
      RECT 14.030000  40.380000 65.090000  40.450000 ;
      RECT 14.030000  40.450000 65.020000  40.520000 ;
      RECT 14.030000  40.450000 65.020000  40.520000 ;
      RECT 14.030000  40.520000 64.950000  40.590000 ;
      RECT 14.030000  40.520000 64.950000  40.590000 ;
      RECT 14.030000  40.590000 64.880000  40.660000 ;
      RECT 14.030000  40.590000 64.880000  40.660000 ;
      RECT 14.030000  40.660000 64.830000  40.710000 ;
      RECT 14.030000  40.660000 64.830000  40.710000 ;
      RECT 14.030000  40.710000 15.855000  43.910000 ;
      RECT 14.030000  40.850000 15.995000  43.770000 ;
      RECT 14.030000  43.770000 65.860000  44.730000 ;
      RECT 14.030000  43.910000 64.845000  43.980000 ;
      RECT 14.030000  43.910000 64.845000  43.980000 ;
      RECT 14.030000  43.980000 64.915000  44.050000 ;
      RECT 14.030000  43.980000 64.915000  44.050000 ;
      RECT 14.030000  44.050000 64.985000  44.120000 ;
      RECT 14.030000  44.050000 64.985000  44.120000 ;
      RECT 14.030000  44.120000 65.055000  44.190000 ;
      RECT 14.030000  44.120000 65.055000  44.190000 ;
      RECT 14.030000  44.190000 65.125000  44.260000 ;
      RECT 14.030000  44.190000 65.125000  44.260000 ;
      RECT 14.030000  44.260000 65.195000  44.330000 ;
      RECT 14.030000  44.260000 65.195000  44.330000 ;
      RECT 14.030000  44.330000 65.265000  44.400000 ;
      RECT 14.030000  44.330000 65.265000  44.400000 ;
      RECT 14.030000  44.400000 65.335000  44.470000 ;
      RECT 14.030000  44.400000 65.335000  44.470000 ;
      RECT 14.030000  44.470000 65.405000  44.540000 ;
      RECT 14.030000  44.470000 65.405000  44.540000 ;
      RECT 14.030000  44.540000 65.475000  44.610000 ;
      RECT 14.030000  44.540000 65.475000  44.610000 ;
      RECT 14.030000  44.610000 65.545000  44.680000 ;
      RECT 14.030000  44.610000 65.545000  44.680000 ;
      RECT 14.030000  44.680000 65.615000  44.750000 ;
      RECT 14.030000  44.680000 65.615000  44.750000 ;
      RECT 14.030000  44.730000 65.860000  49.895000 ;
      RECT 14.030000  44.750000 65.685000  44.785000 ;
      RECT 14.030000  44.750000 65.685000  44.785000 ;
      RECT 14.030000  44.785000 65.720000  49.840000 ;
      RECT 14.030000  49.840000 65.650000  49.910000 ;
      RECT 14.030000  49.840000 65.650000  49.910000 ;
      RECT 14.030000  49.895000 64.885000  50.870000 ;
      RECT 14.030000  49.910000 65.580000  49.980000 ;
      RECT 14.030000  49.910000 65.580000  49.980000 ;
      RECT 14.030000  49.980000 65.510000  50.050000 ;
      RECT 14.030000  49.980000 65.510000  50.050000 ;
      RECT 14.030000  50.050000 65.440000  50.120000 ;
      RECT 14.030000  50.050000 65.440000  50.120000 ;
      RECT 14.030000  50.120000 65.370000  50.190000 ;
      RECT 14.030000  50.120000 65.370000  50.190000 ;
      RECT 14.030000  50.190000 65.300000  50.260000 ;
      RECT 14.030000  50.190000 65.300000  50.260000 ;
      RECT 14.030000  50.260000 65.230000  50.330000 ;
      RECT 14.030000  50.260000 65.230000  50.330000 ;
      RECT 14.030000  50.330000 65.160000  50.400000 ;
      RECT 14.030000  50.330000 65.160000  50.400000 ;
      RECT 14.030000  50.400000 65.090000  50.470000 ;
      RECT 14.030000  50.400000 65.090000  50.470000 ;
      RECT 14.030000  50.470000 65.020000  50.540000 ;
      RECT 14.030000  50.470000 65.020000  50.540000 ;
      RECT 14.030000  50.540000 64.950000  50.610000 ;
      RECT 14.030000  50.540000 64.950000  50.610000 ;
      RECT 14.030000  50.610000 64.880000  50.680000 ;
      RECT 14.030000  50.610000 64.880000  50.680000 ;
      RECT 14.030000  50.680000 64.830000  50.730000 ;
      RECT 14.030000  50.680000 64.830000  50.730000 ;
      RECT 14.030000  50.730000 15.855000  53.930000 ;
      RECT 14.030000  50.870000 15.995000  53.790000 ;
      RECT 14.030000  53.790000 65.855000  54.745000 ;
      RECT 14.030000  53.930000 64.845000  54.000000 ;
      RECT 14.030000  53.930000 64.845000  54.000000 ;
      RECT 14.030000  54.000000 64.915000  54.070000 ;
      RECT 14.030000  54.000000 64.915000  54.070000 ;
      RECT 14.030000  54.070000 64.985000  54.140000 ;
      RECT 14.030000  54.070000 64.985000  54.140000 ;
      RECT 14.030000  54.140000 65.055000  54.210000 ;
      RECT 14.030000  54.140000 65.055000  54.210000 ;
      RECT 14.030000  54.210000 65.125000  54.280000 ;
      RECT 14.030000  54.210000 65.125000  54.280000 ;
      RECT 14.030000  54.280000 65.195000  54.350000 ;
      RECT 14.030000  54.280000 65.195000  54.350000 ;
      RECT 14.030000  54.350000 65.265000  54.420000 ;
      RECT 14.030000  54.350000 65.265000  54.420000 ;
      RECT 14.030000  54.420000 65.335000  54.490000 ;
      RECT 14.030000  54.420000 65.335000  54.490000 ;
      RECT 14.030000  54.490000 65.405000  54.560000 ;
      RECT 14.030000  54.490000 65.405000  54.560000 ;
      RECT 14.030000  54.560000 65.475000  54.630000 ;
      RECT 14.030000  54.560000 65.475000  54.630000 ;
      RECT 14.030000  54.630000 65.545000  54.700000 ;
      RECT 14.030000  54.630000 65.545000  54.700000 ;
      RECT 14.030000  54.700000 65.615000  54.770000 ;
      RECT 14.030000  54.700000 65.615000  54.770000 ;
      RECT 14.030000  54.745000 65.855000  59.880000 ;
      RECT 14.030000  54.770000 65.685000  54.800000 ;
      RECT 14.030000  54.770000 65.685000  54.800000 ;
      RECT 14.030000  54.800000 65.715000  59.825000 ;
      RECT 14.030000  59.825000 65.645000  59.895000 ;
      RECT 14.030000  59.825000 65.645000  59.895000 ;
      RECT 14.030000  59.880000 64.885000  60.850000 ;
      RECT 14.030000  59.895000 65.575000  59.965000 ;
      RECT 14.030000  59.895000 65.575000  59.965000 ;
      RECT 14.030000  59.965000 65.505000  60.035000 ;
      RECT 14.030000  59.965000 65.505000  60.035000 ;
      RECT 14.030000  60.035000 65.435000  60.105000 ;
      RECT 14.030000  60.035000 65.435000  60.105000 ;
      RECT 14.030000  60.105000 65.365000  60.175000 ;
      RECT 14.030000  60.105000 65.365000  60.175000 ;
      RECT 14.030000  60.175000 65.295000  60.245000 ;
      RECT 14.030000  60.175000 65.295000  60.245000 ;
      RECT 14.030000  60.245000 65.225000  60.315000 ;
      RECT 14.030000  60.245000 65.225000  60.315000 ;
      RECT 14.030000  60.315000 65.155000  60.385000 ;
      RECT 14.030000  60.315000 65.155000  60.385000 ;
      RECT 14.030000  60.385000 65.085000  60.455000 ;
      RECT 14.030000  60.385000 65.085000  60.455000 ;
      RECT 14.030000  60.455000 65.015000  60.525000 ;
      RECT 14.030000  60.455000 65.015000  60.525000 ;
      RECT 14.030000  60.525000 64.945000  60.595000 ;
      RECT 14.030000  60.525000 64.945000  60.595000 ;
      RECT 14.030000  60.595000 64.875000  60.665000 ;
      RECT 14.030000  60.595000 64.875000  60.665000 ;
      RECT 14.030000  60.665000 64.830000  60.710000 ;
      RECT 14.030000  60.665000 64.830000  60.710000 ;
      RECT 14.030000  60.710000 15.855000  63.910000 ;
      RECT 14.030000  60.850000 15.995000  63.770000 ;
      RECT 14.030000  63.770000 65.855000  64.735000 ;
      RECT 14.030000  63.910000 64.830000  63.980000 ;
      RECT 14.030000  63.910000 64.830000  63.980000 ;
      RECT 14.030000  63.980000 64.900000  64.050000 ;
      RECT 14.030000  63.980000 64.900000  64.050000 ;
      RECT 14.030000  64.050000 64.970000  64.120000 ;
      RECT 14.030000  64.050000 64.970000  64.120000 ;
      RECT 14.030000  64.120000 65.040000  64.190000 ;
      RECT 14.030000  64.120000 65.040000  64.190000 ;
      RECT 14.030000  64.190000 65.110000  64.260000 ;
      RECT 14.030000  64.190000 65.110000  64.260000 ;
      RECT 14.030000  64.260000 65.180000  64.330000 ;
      RECT 14.030000  64.260000 65.180000  64.330000 ;
      RECT 14.030000  64.330000 65.250000  64.400000 ;
      RECT 14.030000  64.330000 65.250000  64.400000 ;
      RECT 14.030000  64.400000 65.320000  64.470000 ;
      RECT 14.030000  64.400000 65.320000  64.470000 ;
      RECT 14.030000  64.470000 65.390000  64.540000 ;
      RECT 14.030000  64.470000 65.390000  64.540000 ;
      RECT 14.030000  64.540000 65.460000  64.610000 ;
      RECT 14.030000  64.540000 65.460000  64.610000 ;
      RECT 14.030000  64.610000 65.530000  64.680000 ;
      RECT 14.030000  64.610000 65.530000  64.680000 ;
      RECT 14.030000  64.680000 65.600000  64.750000 ;
      RECT 14.030000  64.680000 65.600000  64.750000 ;
      RECT 14.030000  64.735000 65.855000  69.880000 ;
      RECT 14.030000  64.750000 65.670000  64.795000 ;
      RECT 14.030000  64.750000 65.670000  64.795000 ;
      RECT 14.030000  64.795000 65.715000  69.825000 ;
      RECT 14.030000  69.825000 65.645000  69.895000 ;
      RECT 14.030000  69.825000 65.645000  69.895000 ;
      RECT 14.030000  69.880000 64.885000  70.850000 ;
      RECT 14.030000  69.895000 65.575000  69.965000 ;
      RECT 14.030000  69.895000 65.575000  69.965000 ;
      RECT 14.030000  69.965000 65.505000  70.035000 ;
      RECT 14.030000  69.965000 65.505000  70.035000 ;
      RECT 14.030000  70.035000 65.435000  70.105000 ;
      RECT 14.030000  70.035000 65.435000  70.105000 ;
      RECT 14.030000  70.105000 65.365000  70.175000 ;
      RECT 14.030000  70.105000 65.365000  70.175000 ;
      RECT 14.030000  70.175000 65.295000  70.245000 ;
      RECT 14.030000  70.175000 65.295000  70.245000 ;
      RECT 14.030000  70.245000 65.225000  70.315000 ;
      RECT 14.030000  70.245000 65.225000  70.315000 ;
      RECT 14.030000  70.315000 65.155000  70.385000 ;
      RECT 14.030000  70.315000 65.155000  70.385000 ;
      RECT 14.030000  70.385000 65.085000  70.455000 ;
      RECT 14.030000  70.385000 65.085000  70.455000 ;
      RECT 14.030000  70.455000 65.015000  70.525000 ;
      RECT 14.030000  70.455000 65.015000  70.525000 ;
      RECT 14.030000  70.525000 64.945000  70.595000 ;
      RECT 14.030000  70.525000 64.945000  70.595000 ;
      RECT 14.030000  70.595000 64.875000  70.665000 ;
      RECT 14.030000  70.595000 64.875000  70.665000 ;
      RECT 14.030000  70.665000 64.830000  70.710000 ;
      RECT 14.030000  70.665000 64.830000  70.710000 ;
      RECT 14.030000  70.710000 15.855000  73.910000 ;
      RECT 14.030000  70.850000 15.995000  73.770000 ;
      RECT 14.030000  73.770000 65.550000  74.180000 ;
      RECT 14.030000  73.910000 65.085000  73.980000 ;
      RECT 14.030000  73.980000 65.155000  74.050000 ;
      RECT 14.030000  74.050000 65.225000  74.120000 ;
      RECT 14.030000  74.120000 65.295000  74.180000 ;
      RECT 14.030000  74.180000 65.760000  74.390000 ;
      RECT 14.065000  25.265000 65.430000  25.300000 ;
      RECT 14.065000  25.265000 65.430000  25.300000 ;
      RECT 14.100000  74.180000 65.350000  74.250000 ;
      RECT 14.135000  25.195000 65.360000  25.265000 ;
      RECT 14.135000  25.195000 65.360000  25.265000 ;
      RECT 14.170000  74.250000 65.425000  74.320000 ;
      RECT 14.205000  25.125000 65.290000  25.195000 ;
      RECT 14.205000  25.125000 65.290000  25.195000 ;
      RECT 14.240000  73.910000 65.085000  73.980000 ;
      RECT 14.240000  73.910000 65.085000  73.980000 ;
      RECT 14.240000  73.980000 65.155000  74.050000 ;
      RECT 14.240000  73.980000 65.155000  74.050000 ;
      RECT 14.240000  74.050000 65.225000  74.120000 ;
      RECT 14.240000  74.050000 65.225000  74.120000 ;
      RECT 14.240000  74.120000 65.295000  74.180000 ;
      RECT 14.240000  74.120000 65.295000  74.180000 ;
      RECT 14.240000  74.180000 65.350000  74.250000 ;
      RECT 14.240000  74.180000 65.350000  74.250000 ;
      RECT 14.240000  74.250000 65.425000  74.320000 ;
      RECT 14.240000  74.250000 65.425000  74.320000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.390000 65.565000  74.460000 ;
      RECT 14.240000  74.390000 65.565000  74.460000 ;
      RECT 14.240000  74.390000 65.860000  74.490000 ;
      RECT 14.240000  74.460000 65.635000  74.530000 ;
      RECT 14.240000  74.460000 65.635000  74.530000 ;
      RECT 14.240000  74.490000 65.860000  98.700000 ;
      RECT 14.240000  74.530000 65.705000  74.545000 ;
      RECT 14.240000  74.530000 65.705000  74.545000 ;
      RECT 14.240000  74.545000 65.720000  98.840000 ;
      RECT 14.240000  98.700000 75.000000 129.820000 ;
      RECT 14.240000  98.840000 75.000000 129.820000 ;
      RECT 14.240000 129.820000 75.000000 130.705000 ;
      RECT 14.240000 134.795000 75.000000 139.825000 ;
      RECT 14.240000 134.795000 75.000000 139.825000 ;
      RECT 14.240000 139.825000 75.000000 140.710000 ;
      RECT 14.240000 144.795000 75.000000 149.825000 ;
      RECT 14.240000 144.795000 75.000000 149.825000 ;
      RECT 14.240000 149.825000 75.000000 150.710000 ;
      RECT 14.240000 154.795000 75.000000 159.825000 ;
      RECT 14.240000 154.795000 75.000000 159.825000 ;
      RECT 14.240000 159.825000 75.000000 160.710000 ;
      RECT 14.240000 164.795000 75.000000 169.825000 ;
      RECT 14.240000 164.795000 75.000000 169.825000 ;
      RECT 14.240000 169.825000 75.000000 170.710000 ;
      RECT 14.240000 174.795000 75.000000 179.825000 ;
      RECT 14.240000 174.795000 75.000000 179.825000 ;
      RECT 14.240000 179.825000 75.000000 180.710000 ;
      RECT 14.240000 184.795000 75.000000 189.825000 ;
      RECT 14.240000 184.795000 75.000000 189.825000 ;
      RECT 14.240000 189.825000 75.000000 190.710000 ;
      RECT 14.275000  25.055000 65.220000  25.125000 ;
      RECT 14.275000  25.055000 65.220000  25.125000 ;
      RECT 14.285000 134.750000 75.000000 134.795000 ;
      RECT 14.285000 134.750000 75.000000 134.795000 ;
      RECT 14.285000 144.750000 75.000000 144.795000 ;
      RECT 14.285000 144.750000 75.000000 144.795000 ;
      RECT 14.285000 154.750000 75.000000 154.795000 ;
      RECT 14.285000 154.750000 75.000000 154.795000 ;
      RECT 14.285000 164.750000 75.000000 164.795000 ;
      RECT 14.285000 164.750000 75.000000 164.795000 ;
      RECT 14.285000 174.750000 75.000000 174.795000 ;
      RECT 14.285000 174.750000 75.000000 174.795000 ;
      RECT 14.285000 184.750000 75.000000 184.795000 ;
      RECT 14.285000 184.750000 75.000000 184.795000 ;
      RECT 14.310000 129.820000 75.000000 129.890000 ;
      RECT 14.310000 129.820000 75.000000 129.890000 ;
      RECT 14.310000 139.825000 75.000000 139.895000 ;
      RECT 14.310000 139.825000 75.000000 139.895000 ;
      RECT 14.310000 149.825000 75.000000 149.895000 ;
      RECT 14.310000 149.825000 75.000000 149.895000 ;
      RECT 14.310000 159.825000 75.000000 159.895000 ;
      RECT 14.310000 159.825000 75.000000 159.895000 ;
      RECT 14.310000 169.825000 75.000000 169.895000 ;
      RECT 14.310000 169.825000 75.000000 169.895000 ;
      RECT 14.310000 179.825000 75.000000 179.895000 ;
      RECT 14.310000 179.825000 75.000000 179.895000 ;
      RECT 14.310000 189.825000 75.000000 189.895000 ;
      RECT 14.310000 189.825000 75.000000 189.895000 ;
      RECT 14.345000  24.985000 65.150000  25.055000 ;
      RECT 14.345000  24.985000 65.150000  25.055000 ;
      RECT 14.355000 134.680000 75.000000 134.750000 ;
      RECT 14.355000 134.680000 75.000000 134.750000 ;
      RECT 14.355000 144.680000 75.000000 144.750000 ;
      RECT 14.355000 144.680000 75.000000 144.750000 ;
      RECT 14.355000 154.680000 75.000000 154.750000 ;
      RECT 14.355000 154.680000 75.000000 154.750000 ;
      RECT 14.355000 164.680000 75.000000 164.750000 ;
      RECT 14.355000 164.680000 75.000000 164.750000 ;
      RECT 14.355000 174.680000 75.000000 174.750000 ;
      RECT 14.355000 174.680000 75.000000 174.750000 ;
      RECT 14.355000 184.680000 75.000000 184.750000 ;
      RECT 14.355000 184.680000 75.000000 184.750000 ;
      RECT 14.380000 129.890000 75.000000 129.960000 ;
      RECT 14.380000 129.890000 75.000000 129.960000 ;
      RECT 14.380000 139.895000 75.000000 139.965000 ;
      RECT 14.380000 139.895000 75.000000 139.965000 ;
      RECT 14.380000 149.895000 75.000000 149.965000 ;
      RECT 14.380000 149.895000 75.000000 149.965000 ;
      RECT 14.380000 159.895000 75.000000 159.965000 ;
      RECT 14.380000 159.895000 75.000000 159.965000 ;
      RECT 14.380000 169.895000 75.000000 169.965000 ;
      RECT 14.380000 169.895000 75.000000 169.965000 ;
      RECT 14.380000 179.895000 75.000000 179.965000 ;
      RECT 14.380000 179.895000 75.000000 179.965000 ;
      RECT 14.380000 189.895000 75.000000 189.965000 ;
      RECT 14.380000 189.895000 75.000000 189.965000 ;
      RECT 14.415000  24.915000 65.080000  24.985000 ;
      RECT 14.415000  24.915000 65.080000  24.985000 ;
      RECT 14.425000 134.610000 75.000000 134.680000 ;
      RECT 14.425000 134.610000 75.000000 134.680000 ;
      RECT 14.425000 144.610000 75.000000 144.680000 ;
      RECT 14.425000 144.610000 75.000000 144.680000 ;
      RECT 14.425000 154.610000 75.000000 154.680000 ;
      RECT 14.425000 154.610000 75.000000 154.680000 ;
      RECT 14.425000 164.610000 75.000000 164.680000 ;
      RECT 14.425000 164.610000 75.000000 164.680000 ;
      RECT 14.425000 174.610000 75.000000 174.680000 ;
      RECT 14.425000 174.610000 75.000000 174.680000 ;
      RECT 14.425000 184.610000 75.000000 184.680000 ;
      RECT 14.425000 184.610000 75.000000 184.680000 ;
      RECT 14.450000 129.960000 75.000000 130.030000 ;
      RECT 14.450000 129.960000 75.000000 130.030000 ;
      RECT 14.450000 139.965000 75.000000 140.035000 ;
      RECT 14.450000 139.965000 75.000000 140.035000 ;
      RECT 14.450000 149.965000 75.000000 150.035000 ;
      RECT 14.450000 149.965000 75.000000 150.035000 ;
      RECT 14.450000 159.965000 75.000000 160.035000 ;
      RECT 14.450000 159.965000 75.000000 160.035000 ;
      RECT 14.450000 169.965000 75.000000 170.035000 ;
      RECT 14.450000 169.965000 75.000000 170.035000 ;
      RECT 14.450000 179.965000 75.000000 180.035000 ;
      RECT 14.450000 179.965000 75.000000 180.035000 ;
      RECT 14.450000 189.965000 75.000000 190.035000 ;
      RECT 14.450000 189.965000 75.000000 190.035000 ;
      RECT 14.485000  24.845000 65.010000  24.915000 ;
      RECT 14.485000  24.845000 65.010000  24.915000 ;
      RECT 14.495000 134.540000 75.000000 134.610000 ;
      RECT 14.495000 134.540000 75.000000 134.610000 ;
      RECT 14.495000 144.540000 75.000000 144.610000 ;
      RECT 14.495000 144.540000 75.000000 144.610000 ;
      RECT 14.495000 154.540000 75.000000 154.610000 ;
      RECT 14.495000 154.540000 75.000000 154.610000 ;
      RECT 14.495000 164.540000 75.000000 164.610000 ;
      RECT 14.495000 164.540000 75.000000 164.610000 ;
      RECT 14.495000 174.540000 75.000000 174.610000 ;
      RECT 14.495000 174.540000 75.000000 174.610000 ;
      RECT 14.495000 184.540000 75.000000 184.610000 ;
      RECT 14.495000 184.540000 75.000000 184.610000 ;
      RECT 14.520000 130.030000 75.000000 130.100000 ;
      RECT 14.520000 130.030000 75.000000 130.100000 ;
      RECT 14.520000 140.035000 75.000000 140.105000 ;
      RECT 14.520000 140.035000 75.000000 140.105000 ;
      RECT 14.520000 150.035000 75.000000 150.105000 ;
      RECT 14.520000 150.035000 75.000000 150.105000 ;
      RECT 14.520000 160.035000 75.000000 160.105000 ;
      RECT 14.520000 160.035000 75.000000 160.105000 ;
      RECT 14.520000 170.035000 75.000000 170.105000 ;
      RECT 14.520000 170.035000 75.000000 170.105000 ;
      RECT 14.520000 180.035000 75.000000 180.105000 ;
      RECT 14.520000 180.035000 75.000000 180.105000 ;
      RECT 14.520000 190.035000 75.000000 190.105000 ;
      RECT 14.520000 190.035000 75.000000 190.105000 ;
      RECT 14.555000  24.775000 64.940000  24.845000 ;
      RECT 14.555000  24.775000 64.940000  24.845000 ;
      RECT 14.565000 134.470000 75.000000 134.540000 ;
      RECT 14.565000 134.470000 75.000000 134.540000 ;
      RECT 14.565000 144.470000 75.000000 144.540000 ;
      RECT 14.565000 144.470000 75.000000 144.540000 ;
      RECT 14.565000 154.470000 75.000000 154.540000 ;
      RECT 14.565000 154.470000 75.000000 154.540000 ;
      RECT 14.565000 164.470000 75.000000 164.540000 ;
      RECT 14.565000 164.470000 75.000000 164.540000 ;
      RECT 14.565000 174.470000 75.000000 174.540000 ;
      RECT 14.565000 174.470000 75.000000 174.540000 ;
      RECT 14.565000 184.470000 75.000000 184.540000 ;
      RECT 14.565000 184.470000 75.000000 184.540000 ;
      RECT 14.590000 130.100000 75.000000 130.170000 ;
      RECT 14.590000 130.100000 75.000000 130.170000 ;
      RECT 14.590000 140.105000 75.000000 140.175000 ;
      RECT 14.590000 140.105000 75.000000 140.175000 ;
      RECT 14.590000 150.105000 75.000000 150.175000 ;
      RECT 14.590000 150.105000 75.000000 150.175000 ;
      RECT 14.590000 160.105000 75.000000 160.175000 ;
      RECT 14.590000 160.105000 75.000000 160.175000 ;
      RECT 14.590000 170.105000 75.000000 170.175000 ;
      RECT 14.590000 170.105000 75.000000 170.175000 ;
      RECT 14.590000 180.105000 75.000000 180.175000 ;
      RECT 14.590000 180.105000 75.000000 180.175000 ;
      RECT 14.590000 190.105000 75.000000 190.175000 ;
      RECT 14.590000 190.105000 75.000000 190.175000 ;
      RECT 14.625000  24.705000 64.870000  24.775000 ;
      RECT 14.625000  24.705000 64.870000  24.775000 ;
      RECT 14.635000 134.400000 75.000000 134.470000 ;
      RECT 14.635000 134.400000 75.000000 134.470000 ;
      RECT 14.635000 144.400000 75.000000 144.470000 ;
      RECT 14.635000 144.400000 75.000000 144.470000 ;
      RECT 14.635000 154.400000 75.000000 154.470000 ;
      RECT 14.635000 154.400000 75.000000 154.470000 ;
      RECT 14.635000 164.400000 75.000000 164.470000 ;
      RECT 14.635000 164.400000 75.000000 164.470000 ;
      RECT 14.635000 174.400000 75.000000 174.470000 ;
      RECT 14.635000 174.400000 75.000000 174.470000 ;
      RECT 14.635000 184.400000 75.000000 184.470000 ;
      RECT 14.635000 184.400000 75.000000 184.470000 ;
      RECT 14.660000 130.170000 75.000000 130.240000 ;
      RECT 14.660000 130.170000 75.000000 130.240000 ;
      RECT 14.660000 140.175000 75.000000 140.245000 ;
      RECT 14.660000 140.175000 75.000000 140.245000 ;
      RECT 14.660000 150.175000 75.000000 150.245000 ;
      RECT 14.660000 150.175000 75.000000 150.245000 ;
      RECT 14.660000 160.175000 75.000000 160.245000 ;
      RECT 14.660000 160.175000 75.000000 160.245000 ;
      RECT 14.660000 170.175000 75.000000 170.245000 ;
      RECT 14.660000 170.175000 75.000000 170.245000 ;
      RECT 14.660000 180.175000 75.000000 180.245000 ;
      RECT 14.660000 180.175000 75.000000 180.245000 ;
      RECT 14.660000 190.175000 75.000000 190.245000 ;
      RECT 14.660000 190.175000 75.000000 190.245000 ;
      RECT 14.695000  24.635000 64.800000  24.705000 ;
      RECT 14.695000  24.635000 64.800000  24.705000 ;
      RECT 14.705000 134.330000 75.000000 134.400000 ;
      RECT 14.705000 134.330000 75.000000 134.400000 ;
      RECT 14.705000 144.330000 75.000000 144.400000 ;
      RECT 14.705000 144.330000 75.000000 144.400000 ;
      RECT 14.705000 154.330000 75.000000 154.400000 ;
      RECT 14.705000 154.330000 75.000000 154.400000 ;
      RECT 14.705000 164.330000 75.000000 164.400000 ;
      RECT 14.705000 164.330000 75.000000 164.400000 ;
      RECT 14.705000 174.330000 75.000000 174.400000 ;
      RECT 14.705000 174.330000 75.000000 174.400000 ;
      RECT 14.705000 184.330000 75.000000 184.400000 ;
      RECT 14.705000 184.330000 75.000000 184.400000 ;
      RECT 14.730000 130.240000 75.000000 130.310000 ;
      RECT 14.730000 130.240000 75.000000 130.310000 ;
      RECT 14.730000 140.245000 75.000000 140.315000 ;
      RECT 14.730000 140.245000 75.000000 140.315000 ;
      RECT 14.730000 150.245000 75.000000 150.315000 ;
      RECT 14.730000 150.245000 75.000000 150.315000 ;
      RECT 14.730000 160.245000 75.000000 160.315000 ;
      RECT 14.730000 160.245000 75.000000 160.315000 ;
      RECT 14.730000 170.245000 75.000000 170.315000 ;
      RECT 14.730000 170.245000 75.000000 170.315000 ;
      RECT 14.730000 180.245000 75.000000 180.315000 ;
      RECT 14.730000 180.245000 75.000000 180.315000 ;
      RECT 14.730000 190.245000 75.000000 190.315000 ;
      RECT 14.730000 190.245000 75.000000 190.315000 ;
      RECT 14.765000  24.565000 64.730000  24.635000 ;
      RECT 14.765000  24.565000 64.730000  24.635000 ;
      RECT 14.775000 134.260000 75.000000 134.330000 ;
      RECT 14.775000 134.260000 75.000000 134.330000 ;
      RECT 14.775000 144.260000 75.000000 144.330000 ;
      RECT 14.775000 144.260000 75.000000 144.330000 ;
      RECT 14.775000 154.260000 75.000000 154.330000 ;
      RECT 14.775000 154.260000 75.000000 154.330000 ;
      RECT 14.775000 164.260000 75.000000 164.330000 ;
      RECT 14.775000 164.260000 75.000000 164.330000 ;
      RECT 14.775000 174.260000 75.000000 174.330000 ;
      RECT 14.775000 174.260000 75.000000 174.330000 ;
      RECT 14.775000 184.260000 75.000000 184.330000 ;
      RECT 14.775000 184.260000 75.000000 184.330000 ;
      RECT 14.800000 130.310000 75.000000 130.380000 ;
      RECT 14.800000 130.310000 75.000000 130.380000 ;
      RECT 14.800000 140.315000 75.000000 140.385000 ;
      RECT 14.800000 140.315000 75.000000 140.385000 ;
      RECT 14.800000 150.315000 75.000000 150.385000 ;
      RECT 14.800000 150.315000 75.000000 150.385000 ;
      RECT 14.800000 160.315000 75.000000 160.385000 ;
      RECT 14.800000 160.315000 75.000000 160.385000 ;
      RECT 14.800000 170.315000 75.000000 170.385000 ;
      RECT 14.800000 170.315000 75.000000 170.385000 ;
      RECT 14.800000 180.315000 75.000000 180.385000 ;
      RECT 14.800000 180.315000 75.000000 180.385000 ;
      RECT 14.800000 190.315000 75.000000 190.385000 ;
      RECT 14.800000 190.315000 75.000000 190.385000 ;
      RECT 14.835000  24.495000 64.660000  24.565000 ;
      RECT 14.835000  24.495000 64.660000  24.565000 ;
      RECT 14.845000 134.190000 75.000000 134.260000 ;
      RECT 14.845000 134.190000 75.000000 134.260000 ;
      RECT 14.845000 144.190000 75.000000 144.260000 ;
      RECT 14.845000 144.190000 75.000000 144.260000 ;
      RECT 14.845000 154.190000 75.000000 154.260000 ;
      RECT 14.845000 154.190000 75.000000 154.260000 ;
      RECT 14.845000 164.190000 75.000000 164.260000 ;
      RECT 14.845000 164.190000 75.000000 164.260000 ;
      RECT 14.845000 174.190000 75.000000 174.260000 ;
      RECT 14.845000 174.190000 75.000000 174.260000 ;
      RECT 14.845000 184.190000 75.000000 184.260000 ;
      RECT 14.845000 184.190000 75.000000 184.260000 ;
      RECT 14.870000 130.380000 75.000000 130.450000 ;
      RECT 14.870000 130.380000 75.000000 130.450000 ;
      RECT 14.870000 140.385000 75.000000 140.455000 ;
      RECT 14.870000 140.385000 75.000000 140.455000 ;
      RECT 14.870000 150.385000 75.000000 150.455000 ;
      RECT 14.870000 150.385000 75.000000 150.455000 ;
      RECT 14.870000 160.385000 75.000000 160.455000 ;
      RECT 14.870000 160.385000 75.000000 160.455000 ;
      RECT 14.870000 170.385000 75.000000 170.455000 ;
      RECT 14.870000 170.385000 75.000000 170.455000 ;
      RECT 14.870000 180.385000 75.000000 180.455000 ;
      RECT 14.870000 180.385000 75.000000 180.455000 ;
      RECT 14.870000 190.385000 75.000000 190.455000 ;
      RECT 14.870000 190.385000 75.000000 190.455000 ;
      RECT 14.905000  24.425000 64.590000  24.495000 ;
      RECT 14.905000  24.425000 64.590000  24.495000 ;
      RECT 14.915000 134.120000 75.000000 134.190000 ;
      RECT 14.915000 134.120000 75.000000 134.190000 ;
      RECT 14.915000 144.120000 75.000000 144.190000 ;
      RECT 14.915000 144.120000 75.000000 144.190000 ;
      RECT 14.915000 154.120000 75.000000 154.190000 ;
      RECT 14.915000 154.120000 75.000000 154.190000 ;
      RECT 14.915000 164.120000 75.000000 164.190000 ;
      RECT 14.915000 164.120000 75.000000 164.190000 ;
      RECT 14.915000 174.120000 75.000000 174.190000 ;
      RECT 14.915000 174.120000 75.000000 174.190000 ;
      RECT 14.915000 184.120000 75.000000 184.190000 ;
      RECT 14.915000 184.120000 75.000000 184.190000 ;
      RECT 14.940000 130.450000 75.000000 130.520000 ;
      RECT 14.940000 130.450000 75.000000 130.520000 ;
      RECT 14.940000 140.455000 75.000000 140.525000 ;
      RECT 14.940000 140.455000 75.000000 140.525000 ;
      RECT 14.940000 150.455000 75.000000 150.525000 ;
      RECT 14.940000 150.455000 75.000000 150.525000 ;
      RECT 14.940000 160.455000 75.000000 160.525000 ;
      RECT 14.940000 160.455000 75.000000 160.525000 ;
      RECT 14.940000 170.455000 75.000000 170.525000 ;
      RECT 14.940000 170.455000 75.000000 170.525000 ;
      RECT 14.940000 180.455000 75.000000 180.525000 ;
      RECT 14.940000 180.455000 75.000000 180.525000 ;
      RECT 14.940000 190.455000 75.000000 190.525000 ;
      RECT 14.940000 190.455000 75.000000 190.525000 ;
      RECT 14.975000  24.355000 64.520000  24.425000 ;
      RECT 14.975000  24.355000 64.520000  24.425000 ;
      RECT 14.985000 134.050000 75.000000 134.120000 ;
      RECT 14.985000 134.050000 75.000000 134.120000 ;
      RECT 14.985000 144.050000 75.000000 144.120000 ;
      RECT 14.985000 144.050000 75.000000 144.120000 ;
      RECT 14.985000 154.050000 75.000000 154.120000 ;
      RECT 14.985000 154.050000 75.000000 154.120000 ;
      RECT 14.985000 164.050000 75.000000 164.120000 ;
      RECT 14.985000 164.050000 75.000000 164.120000 ;
      RECT 14.985000 174.050000 75.000000 174.120000 ;
      RECT 14.985000 174.050000 75.000000 174.120000 ;
      RECT 14.985000 184.050000 75.000000 184.120000 ;
      RECT 14.985000 184.050000 75.000000 184.120000 ;
      RECT 15.010000 130.520000 75.000000 130.590000 ;
      RECT 15.010000 130.520000 75.000000 130.590000 ;
      RECT 15.010000 140.525000 75.000000 140.595000 ;
      RECT 15.010000 140.525000 75.000000 140.595000 ;
      RECT 15.010000 150.525000 75.000000 150.595000 ;
      RECT 15.010000 150.525000 75.000000 150.595000 ;
      RECT 15.010000 160.525000 75.000000 160.595000 ;
      RECT 15.010000 160.525000 75.000000 160.595000 ;
      RECT 15.010000 170.525000 75.000000 170.595000 ;
      RECT 15.010000 170.525000 75.000000 170.595000 ;
      RECT 15.010000 180.525000 75.000000 180.595000 ;
      RECT 15.010000 180.525000 75.000000 180.595000 ;
      RECT 15.010000 190.525000 75.000000 190.595000 ;
      RECT 15.010000 190.525000 75.000000 190.595000 ;
      RECT 15.045000  24.285000 64.450000  24.355000 ;
      RECT 15.045000  24.285000 64.450000  24.355000 ;
      RECT 15.055000 133.980000 75.000000 134.050000 ;
      RECT 15.055000 133.980000 75.000000 134.050000 ;
      RECT 15.055000 143.980000 75.000000 144.050000 ;
      RECT 15.055000 143.980000 75.000000 144.050000 ;
      RECT 15.055000 153.980000 75.000000 154.050000 ;
      RECT 15.055000 153.980000 75.000000 154.050000 ;
      RECT 15.055000 163.980000 75.000000 164.050000 ;
      RECT 15.055000 163.980000 75.000000 164.050000 ;
      RECT 15.055000 173.980000 75.000000 174.050000 ;
      RECT 15.055000 173.980000 75.000000 174.050000 ;
      RECT 15.055000 183.980000 75.000000 184.050000 ;
      RECT 15.055000 183.980000 75.000000 184.050000 ;
      RECT 15.080000 130.590000 75.000000 130.660000 ;
      RECT 15.080000 130.590000 75.000000 130.660000 ;
      RECT 15.080000 140.595000 75.000000 140.665000 ;
      RECT 15.080000 140.595000 75.000000 140.665000 ;
      RECT 15.080000 150.595000 75.000000 150.665000 ;
      RECT 15.080000 150.595000 75.000000 150.665000 ;
      RECT 15.080000 160.595000 75.000000 160.665000 ;
      RECT 15.080000 160.595000 75.000000 160.665000 ;
      RECT 15.080000 170.595000 75.000000 170.665000 ;
      RECT 15.080000 170.595000 75.000000 170.665000 ;
      RECT 15.080000 180.595000 75.000000 180.665000 ;
      RECT 15.080000 180.595000 75.000000 180.665000 ;
      RECT 15.080000 190.595000 75.000000 190.665000 ;
      RECT 15.080000 190.595000 75.000000 190.665000 ;
      RECT 15.115000  24.215000 64.380000  24.285000 ;
      RECT 15.115000  24.215000 64.380000  24.285000 ;
      RECT 15.125000 130.660000 75.000000 130.705000 ;
      RECT 15.125000 130.660000 75.000000 130.705000 ;
      RECT 15.125000 133.910000 75.000000 133.980000 ;
      RECT 15.125000 133.910000 75.000000 133.980000 ;
      RECT 15.125000 133.910000 75.000000 134.795000 ;
      RECT 15.125000 140.665000 75.000000 140.710000 ;
      RECT 15.125000 140.665000 75.000000 140.710000 ;
      RECT 15.125000 143.910000 75.000000 143.980000 ;
      RECT 15.125000 143.910000 75.000000 143.980000 ;
      RECT 15.125000 143.910000 75.000000 144.795000 ;
      RECT 15.125000 150.665000 75.000000 150.710000 ;
      RECT 15.125000 150.665000 75.000000 150.710000 ;
      RECT 15.125000 153.910000 75.000000 153.980000 ;
      RECT 15.125000 153.910000 75.000000 153.980000 ;
      RECT 15.125000 153.910000 75.000000 154.795000 ;
      RECT 15.125000 160.665000 75.000000 160.710000 ;
      RECT 15.125000 160.665000 75.000000 160.710000 ;
      RECT 15.125000 163.910000 75.000000 163.980000 ;
      RECT 15.125000 163.910000 75.000000 163.980000 ;
      RECT 15.125000 163.910000 75.000000 164.795000 ;
      RECT 15.125000 170.665000 75.000000 170.710000 ;
      RECT 15.125000 170.665000 75.000000 170.710000 ;
      RECT 15.125000 173.910000 75.000000 173.980000 ;
      RECT 15.125000 173.910000 75.000000 173.980000 ;
      RECT 15.125000 173.910000 75.000000 174.795000 ;
      RECT 15.125000 180.665000 75.000000 180.710000 ;
      RECT 15.125000 180.665000 75.000000 180.710000 ;
      RECT 15.125000 183.910000 75.000000 183.980000 ;
      RECT 15.125000 183.910000 75.000000 183.980000 ;
      RECT 15.125000 183.910000 75.000000 184.795000 ;
      RECT 15.125000 190.665000 75.000000 190.710000 ;
      RECT 15.125000 190.665000 75.000000 190.710000 ;
      RECT 15.185000  24.145000 64.310000  24.215000 ;
      RECT 15.185000  24.145000 64.310000  24.215000 ;
      RECT 15.255000  24.075000 64.240000  24.145000 ;
      RECT 15.255000  24.075000 64.240000  24.145000 ;
      RECT 15.325000  24.005000 64.170000  24.075000 ;
      RECT 15.325000  24.005000 64.170000  24.075000 ;
      RECT 15.395000  23.935000 64.100000  24.005000 ;
      RECT 15.395000  23.935000 64.100000  24.005000 ;
      RECT 15.465000  23.865000 64.030000  23.935000 ;
      RECT 15.465000  23.865000 64.030000  23.935000 ;
      RECT 15.520000 130.705000 75.000000 130.845000 ;
      RECT 15.520000 140.710000 75.000000 140.850000 ;
      RECT 15.520000 150.710000 75.000000 150.850000 ;
      RECT 15.520000 160.710000 75.000000 160.850000 ;
      RECT 15.520000 170.710000 75.000000 170.850000 ;
      RECT 15.520000 180.710000 75.000000 180.850000 ;
      RECT 15.520000 190.710000 75.000000 190.850000 ;
      RECT 15.535000  23.795000 63.960000  23.865000 ;
      RECT 15.535000  23.795000 63.960000  23.865000 ;
      RECT 15.605000  23.725000 63.890000  23.795000 ;
      RECT 15.605000  23.725000 63.890000  23.795000 ;
      RECT 15.660000 133.770000 75.000000 133.910000 ;
      RECT 15.660000 143.770000 75.000000 143.910000 ;
      RECT 15.660000 153.770000 75.000000 153.910000 ;
      RECT 15.660000 163.770000 75.000000 163.910000 ;
      RECT 15.660000 173.770000 75.000000 173.910000 ;
      RECT 15.660000 183.770000 75.000000 183.910000 ;
      RECT 15.675000  23.655000 63.820000  23.725000 ;
      RECT 15.675000  23.655000 63.820000  23.725000 ;
      RECT 15.745000  23.585000 63.750000  23.655000 ;
      RECT 15.745000  23.585000 63.750000  23.655000 ;
      RECT 15.815000  23.515000 63.680000  23.585000 ;
      RECT 15.815000  23.515000 63.680000  23.585000 ;
      RECT 15.885000  23.445000 63.610000  23.515000 ;
      RECT 15.885000  23.445000 63.610000  23.515000 ;
      RECT 15.955000  23.375000 63.540000  23.445000 ;
      RECT 15.955000  23.375000 63.540000  23.445000 ;
      RECT 16.025000  23.305000 63.470000  23.375000 ;
      RECT 16.025000  23.305000 63.470000  23.375000 ;
      RECT 16.095000  23.235000 63.400000  23.305000 ;
      RECT 16.095000  23.235000 63.400000  23.305000 ;
      RECT 16.165000  23.165000 63.330000  23.235000 ;
      RECT 16.165000  23.165000 63.330000  23.235000 ;
      RECT 16.235000  23.095000 63.260000  23.165000 ;
      RECT 16.235000  23.095000 63.260000  23.165000 ;
      RECT 16.305000  23.025000 63.190000  23.095000 ;
      RECT 16.305000  23.025000 63.190000  23.095000 ;
      RECT 16.375000  22.955000 63.120000  23.025000 ;
      RECT 16.375000  22.955000 63.120000  23.025000 ;
      RECT 16.445000  22.885000 63.050000  22.955000 ;
      RECT 16.445000  22.885000 63.050000  22.955000 ;
      RECT 16.515000  22.815000 62.980000  22.885000 ;
      RECT 16.515000  22.815000 62.980000  22.885000 ;
      RECT 16.585000  22.745000 62.910000  22.815000 ;
      RECT 16.585000  22.745000 62.910000  22.815000 ;
      RECT 16.655000  22.675000 62.840000  22.745000 ;
      RECT 16.655000  22.675000 62.840000  22.745000 ;
      RECT 16.725000  22.605000 62.770000  22.675000 ;
      RECT 16.725000  22.605000 62.770000  22.675000 ;
      RECT 16.795000  22.535000 62.700000  22.605000 ;
      RECT 16.795000  22.535000 62.700000  22.605000 ;
      RECT 16.865000  22.465000 62.630000  22.535000 ;
      RECT 16.865000  22.465000 62.630000  22.535000 ;
      RECT 16.935000  22.395000 62.560000  22.465000 ;
      RECT 16.935000  22.395000 62.560000  22.465000 ;
      RECT 17.005000  22.325000 62.490000  22.395000 ;
      RECT 17.005000  22.325000 62.490000  22.395000 ;
      RECT 17.075000  22.255000 62.420000  22.325000 ;
      RECT 17.075000  22.255000 62.420000  22.325000 ;
      RECT 17.140000   5.235000 17.350000   9.250000 ;
      RECT 17.140000   5.235000 17.490000   9.250000 ;
      RECT 17.140000   9.250000 17.490000   9.600000 ;
      RECT 17.145000  22.185000 62.350000  22.255000 ;
      RECT 17.145000  22.185000 62.350000  22.255000 ;
      RECT 17.210000   5.165000 17.350000   5.235000 ;
      RECT 17.210000   9.250000 17.350000   9.320000 ;
      RECT 17.215000  22.115000 62.280000  22.185000 ;
      RECT 17.215000  22.115000 62.280000  22.185000 ;
      RECT 17.280000   5.095000 17.350000   5.165000 ;
      RECT 17.280000   9.320000 17.350000   9.390000 ;
      RECT 17.285000  22.045000 62.210000  22.115000 ;
      RECT 17.285000  22.045000 62.210000  22.115000 ;
      RECT 17.320000   5.055000 17.490000   5.235000 ;
      RECT 17.355000  21.975000 62.140000  22.045000 ;
      RECT 17.355000  21.975000 62.140000  22.045000 ;
      RECT 17.425000  21.905000 53.815000  21.975000 ;
      RECT 17.425000  21.905000 53.815000  21.975000 ;
      RECT 17.495000  21.835000 53.815000  21.905000 ;
      RECT 17.495000  21.835000 53.815000  21.905000 ;
      RECT 17.495000  21.835000 65.660000  25.300000 ;
      RECT 17.565000  21.765000 53.815000  21.835000 ;
      RECT 17.565000  21.765000 53.815000  21.835000 ;
      RECT 17.570000   9.680000 55.880000   9.800000 ;
      RECT 17.635000  21.695000 53.815000  21.765000 ;
      RECT 17.635000  21.695000 53.815000  21.765000 ;
      RECT 17.705000  21.625000 53.815000  21.695000 ;
      RECT 17.705000  21.625000 53.815000  21.695000 ;
      RECT 17.775000  21.555000 53.815000  21.625000 ;
      RECT 17.775000  21.555000 53.815000  21.625000 ;
      RECT 17.845000  21.485000 53.815000  21.555000 ;
      RECT 17.845000  21.485000 53.815000  21.555000 ;
      RECT 17.915000  21.415000 53.815000  21.485000 ;
      RECT 17.915000  21.415000 53.815000  21.485000 ;
      RECT 17.985000  21.345000 53.815000  21.415000 ;
      RECT 17.985000  21.345000 53.815000  21.415000 ;
      RECT 18.055000  21.275000 53.815000  21.345000 ;
      RECT 18.055000  21.275000 53.815000  21.345000 ;
      RECT 18.125000  21.205000 53.815000  21.275000 ;
      RECT 18.125000  21.205000 53.815000  21.275000 ;
      RECT 18.195000  21.135000 53.815000  21.205000 ;
      RECT 18.195000  21.135000 53.815000  21.205000 ;
      RECT 18.265000  21.065000 53.815000  21.135000 ;
      RECT 18.265000  21.065000 53.815000  21.135000 ;
      RECT 18.335000  20.995000 53.815000  21.065000 ;
      RECT 18.335000  20.995000 53.815000  21.065000 ;
      RECT 18.405000  20.925000 53.815000  20.995000 ;
      RECT 18.405000  20.925000 53.815000  20.995000 ;
      RECT 18.475000  20.855000 53.815000  20.925000 ;
      RECT 18.475000  20.855000 53.815000  20.925000 ;
      RECT 18.545000  20.785000 53.815000  20.855000 ;
      RECT 18.545000  20.785000 53.815000  20.855000 ;
      RECT 18.580000 193.770000 75.000000 193.910000 ;
      RECT 18.615000  20.715000 53.815000  20.785000 ;
      RECT 18.615000  20.715000 53.815000  20.785000 ;
      RECT 18.685000  20.645000 53.815000  20.715000 ;
      RECT 18.685000  20.645000 53.815000  20.715000 ;
      RECT 18.755000  20.575000 53.815000  20.645000 ;
      RECT 18.755000  20.575000 53.815000  20.645000 ;
      RECT 18.825000  20.505000 53.815000  20.575000 ;
      RECT 18.825000  20.505000 53.815000  20.575000 ;
      RECT 18.895000  20.435000 53.815000  20.505000 ;
      RECT 18.895000  20.435000 53.815000  20.505000 ;
      RECT 18.965000  20.365000 53.815000  20.435000 ;
      RECT 18.965000  20.365000 53.815000  20.435000 ;
      RECT 19.035000  20.295000 53.815000  20.365000 ;
      RECT 19.035000  20.295000 53.815000  20.365000 ;
      RECT 19.105000  20.225000 53.815000  20.295000 ;
      RECT 19.105000  20.225000 53.815000  20.295000 ;
      RECT 19.175000  20.155000 53.815000  20.225000 ;
      RECT 19.175000  20.155000 53.815000  20.225000 ;
      RECT 19.245000  20.085000 53.815000  20.155000 ;
      RECT 19.245000  20.085000 53.815000  20.155000 ;
      RECT 19.315000  20.015000 53.815000  20.085000 ;
      RECT 19.315000  20.015000 53.815000  20.085000 ;
      RECT 19.385000  19.945000 53.815000  20.015000 ;
      RECT 19.385000  19.945000 53.815000  20.015000 ;
      RECT 19.400000  19.930000 53.955000  21.835000 ;
      RECT 19.455000  19.875000 53.815000  19.945000 ;
      RECT 19.455000  19.875000 53.815000  19.945000 ;
      RECT 19.510000  19.820000 53.815000  19.875000 ;
      RECT 19.510000  19.820000 53.815000  19.875000 ;
      RECT 19.580000  19.750000 53.870000  19.820000 ;
      RECT 19.580000  19.750000 53.870000  19.820000 ;
      RECT 19.650000  19.680000 53.940000  19.750000 ;
      RECT 19.650000  19.680000 53.940000  19.750000 ;
      RECT 19.720000  19.610000 54.010000  19.680000 ;
      RECT 19.720000  19.610000 54.010000  19.680000 ;
      RECT 19.790000  19.540000 54.080000  19.610000 ;
      RECT 19.790000  19.540000 54.080000  19.610000 ;
      RECT 19.860000  19.470000 54.150000  19.540000 ;
      RECT 19.860000  19.470000 54.150000  19.540000 ;
      RECT 19.930000  19.400000 54.220000  19.470000 ;
      RECT 19.930000  19.400000 54.220000  19.470000 ;
      RECT 20.000000  19.330000 54.290000  19.400000 ;
      RECT 20.000000  19.330000 54.290000  19.400000 ;
      RECT 20.070000  19.260000 54.360000  19.330000 ;
      RECT 20.070000  19.260000 54.360000  19.330000 ;
      RECT 20.140000  19.190000 54.430000  19.260000 ;
      RECT 20.140000  19.190000 54.430000  19.260000 ;
      RECT 20.210000  19.120000 54.500000  19.190000 ;
      RECT 20.210000  19.120000 54.500000  19.190000 ;
      RECT 20.280000  19.050000 54.570000  19.120000 ;
      RECT 20.280000  19.050000 54.570000  19.120000 ;
      RECT 20.350000  18.980000 54.640000  19.050000 ;
      RECT 20.350000  18.980000 54.640000  19.050000 ;
      RECT 20.420000  18.910000 54.710000  18.980000 ;
      RECT 20.420000  18.910000 54.710000  18.980000 ;
      RECT 20.490000  18.840000 54.780000  18.910000 ;
      RECT 20.490000  18.840000 54.780000  18.910000 ;
      RECT 20.560000  18.770000 54.850000  18.840000 ;
      RECT 20.560000  18.770000 54.850000  18.840000 ;
      RECT 20.630000  18.700000 54.920000  18.770000 ;
      RECT 20.630000  18.700000 54.920000  18.770000 ;
      RECT 20.700000  18.630000 54.990000  18.700000 ;
      RECT 20.700000  18.630000 54.990000  18.700000 ;
      RECT 20.770000  18.560000 55.060000  18.630000 ;
      RECT 20.770000  18.560000 55.060000  18.630000 ;
      RECT 20.775000   0.000000 20.785000   1.600000 ;
      RECT 20.775000   1.600000 20.785000   1.760000 ;
      RECT 20.840000  18.490000 55.130000  18.560000 ;
      RECT 20.840000  18.490000 55.130000  18.560000 ;
      RECT 20.910000  18.420000 55.200000  18.490000 ;
      RECT 20.910000  18.420000 55.200000  18.490000 ;
      RECT 20.980000  18.350000 55.270000  18.420000 ;
      RECT 20.980000  18.350000 55.270000  18.420000 ;
      RECT 21.050000  18.280000 55.340000  18.350000 ;
      RECT 21.050000  18.280000 55.340000  18.350000 ;
      RECT 21.120000  18.210000 55.410000  18.280000 ;
      RECT 21.120000  18.210000 55.410000  18.280000 ;
      RECT 21.190000  18.140000 55.480000  18.210000 ;
      RECT 21.190000  18.140000 55.480000  18.210000 ;
      RECT 21.260000  18.070000 55.550000  18.140000 ;
      RECT 21.260000  18.070000 55.550000  18.140000 ;
      RECT 21.330000  18.000000 55.620000  18.070000 ;
      RECT 21.330000  18.000000 55.620000  18.070000 ;
      RECT 21.400000  17.930000 55.690000  18.000000 ;
      RECT 21.400000  17.930000 55.690000  18.000000 ;
      RECT 21.470000  17.860000 55.760000  17.930000 ;
      RECT 21.470000  17.860000 55.760000  17.930000 ;
      RECT 21.540000  17.790000 55.830000  17.860000 ;
      RECT 21.540000  17.790000 55.830000  17.860000 ;
      RECT 21.555000  17.775000 53.955000  19.930000 ;
      RECT 21.610000  17.720000 55.900000  17.790000 ;
      RECT 21.610000  17.720000 55.900000  17.790000 ;
      RECT 21.620000  17.710000 55.970000  17.720000 ;
      RECT 21.620000  17.710000 55.970000  17.720000 ;
      RECT 21.690000  17.640000 55.970000  17.710000 ;
      RECT 21.690000  17.640000 55.970000  17.710000 ;
      RECT 21.760000  17.570000 55.970000  17.640000 ;
      RECT 21.760000  17.570000 55.970000  17.640000 ;
      RECT 21.830000  17.500000 55.970000  17.570000 ;
      RECT 21.830000  17.500000 55.970000  17.570000 ;
      RECT 21.900000  17.430000 55.970000  17.500000 ;
      RECT 21.900000  17.430000 55.970000  17.500000 ;
      RECT 21.970000  17.360000 55.970000  17.430000 ;
      RECT 21.970000  17.360000 55.970000  17.430000 ;
      RECT 21.970000  17.360000 56.110000  17.775000 ;
      RECT 53.675000   0.000000 53.955000   7.875000 ;
      RECT 53.675000   7.875000 55.760000   9.680000 ;
      RECT 53.815000   8.000000 53.885000   8.070000 ;
      RECT 53.815000   8.070000 53.955000   8.140000 ;
      RECT 53.815000   8.140000 54.025000   8.210000 ;
      RECT 53.815000   8.210000 54.095000   8.280000 ;
      RECT 53.815000   8.280000 54.165000   8.350000 ;
      RECT 53.815000   8.350000 54.235000   8.420000 ;
      RECT 53.815000   8.420000 54.305000   8.490000 ;
      RECT 53.815000   8.490000 54.375000   8.560000 ;
      RECT 53.815000   8.560000 54.445000   8.630000 ;
      RECT 53.815000   8.630000 54.515000   8.700000 ;
      RECT 53.815000   8.700000 54.585000   8.770000 ;
      RECT 53.815000   8.770000 54.655000   8.840000 ;
      RECT 53.815000   8.840000 54.725000   8.910000 ;
      RECT 53.815000   8.910000 54.795000   8.980000 ;
      RECT 53.815000   8.980000 54.865000   9.050000 ;
      RECT 53.815000   9.050000 54.935000   9.120000 ;
      RECT 53.815000   9.120000 55.005000   9.190000 ;
      RECT 53.815000   9.190000 55.075000   9.260000 ;
      RECT 53.815000   9.260000 55.145000   9.330000 ;
      RECT 53.815000   9.330000 55.215000   9.400000 ;
      RECT 53.815000   9.400000 55.285000   9.470000 ;
      RECT 53.815000   9.470000 55.355000   9.540000 ;
      RECT 53.815000   9.540000 55.425000   9.610000 ;
      RECT 53.815000   9.610000 55.495000   9.680000 ;
      RECT 53.815000   9.680000 55.565000   9.750000 ;
      RECT 53.815000   9.750000 55.635000   9.800000 ;
      RECT 55.875000   9.800000 56.110000  10.030000 ;
      RECT 55.875000  10.030000 56.110000  17.360000 ;
      RECT 68.150000  74.490000 75.000000  98.700000 ;
      RECT 68.150000 130.845000 75.000000 133.770000 ;
      RECT 68.150000 140.850000 75.000000 143.770000 ;
      RECT 68.150000 150.850000 75.000000 153.770000 ;
      RECT 68.150000 160.850000 75.000000 163.770000 ;
      RECT 68.150000 170.850000 75.000000 173.770000 ;
      RECT 68.150000 180.850000 75.000000 183.770000 ;
      RECT 68.150000 190.850000 75.000000 193.770000 ;
      RECT 68.290000  74.545000 75.000000  98.840000 ;
      RECT 68.290000 130.705000 75.000000 133.910000 ;
      RECT 68.290000 140.710000 75.000000 143.910000 ;
      RECT 68.290000 150.710000 75.000000 153.910000 ;
      RECT 68.290000 160.710000 75.000000 163.910000 ;
      RECT 68.290000 170.710000 75.000000 173.910000 ;
      RECT 68.290000 180.710000 75.000000 183.910000 ;
      RECT 68.290000 190.710000 75.000000 193.910000 ;
      RECT 68.295000  74.540000 75.000000  74.545000 ;
      RECT 68.295000  74.540000 75.000000  74.545000 ;
      RECT 68.365000  74.470000 75.000000  74.540000 ;
      RECT 68.365000  74.470000 75.000000  74.540000 ;
      RECT 68.435000  74.400000 75.000000  74.470000 ;
      RECT 68.435000  74.400000 75.000000  74.470000 ;
      RECT 68.505000  74.330000 75.000000  74.400000 ;
      RECT 68.505000  74.330000 75.000000  74.400000 ;
      RECT 68.575000  74.260000 75.000000  74.330000 ;
      RECT 68.575000  74.260000 75.000000  74.330000 ;
      RECT 68.645000  74.190000 75.000000  74.260000 ;
      RECT 68.645000  74.190000 75.000000  74.260000 ;
      RECT 68.715000  74.120000 75.000000  74.190000 ;
      RECT 68.715000  74.120000 75.000000  74.190000 ;
      RECT 68.785000  74.050000 75.000000  74.120000 ;
      RECT 68.785000  74.050000 75.000000  74.120000 ;
      RECT 68.855000  73.980000 75.000000  74.050000 ;
      RECT 68.855000  73.980000 75.000000  74.050000 ;
      RECT 68.865000  73.770000 75.000000  74.490000 ;
      RECT 68.925000  73.910000 75.000000  73.980000 ;
      RECT 68.925000  73.910000 75.000000  73.980000 ;
      RECT 74.840000   0.000000 75.000000  73.770000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.200000 171.495000 ;
      RECT  0.000000 171.495000 15.205000 189.915000 ;
      RECT  0.000000 171.595000 15.205000 189.915000 ;
      RECT  0.000000 171.595000 15.205000 198.000000 ;
      RECT  0.000000 189.915000 75.000000 198.000000 ;
      RECT  0.000000 189.915000 75.000000 198.000000 ;
      RECT 13.200000  94.385000 15.205000 171.495000 ;
      RECT 13.300000  94.425000 15.205000 171.595000 ;
      RECT 13.440000  94.145000 15.205000  94.385000 ;
      RECT 13.440000  94.285000 15.205000  94.425000 ;
      RECT 13.580000  94.145000 15.205000  94.285000 ;
      RECT 13.725000  94.000000 15.205000  94.145000 ;
      RECT 13.875000  93.850000 15.350000  94.000000 ;
      RECT 14.025000  93.700000 15.500000  93.850000 ;
      RECT 14.175000  93.550000 15.650000  93.700000 ;
      RECT 14.325000  93.400000 15.800000  93.550000 ;
      RECT 14.475000  93.250000 15.950000  93.400000 ;
      RECT 14.625000  93.100000 16.100000  93.250000 ;
      RECT 14.775000  92.950000 16.250000  93.100000 ;
      RECT 14.925000  92.800000 16.400000  92.950000 ;
      RECT 15.075000  92.650000 16.550000  92.800000 ;
      RECT 15.225000  92.500000 16.700000  92.650000 ;
      RECT 15.375000  92.350000 16.850000  92.500000 ;
      RECT 15.525000  92.200000 17.000000  92.350000 ;
      RECT 15.675000  92.050000 17.150000  92.200000 ;
      RECT 15.825000  91.900000 17.300000  92.050000 ;
      RECT 15.975000  91.750000 17.450000  91.900000 ;
      RECT 16.125000  91.600000 17.600000  91.750000 ;
      RECT 16.275000  91.450000 17.750000  91.600000 ;
      RECT 16.425000  91.300000 17.900000  91.450000 ;
      RECT 16.575000  91.150000 18.050000  91.300000 ;
      RECT 16.725000  91.000000 18.200000  91.150000 ;
      RECT 16.875000  90.850000 18.350000  91.000000 ;
      RECT 17.025000  90.700000 18.500000  90.850000 ;
      RECT 17.175000  90.550000 18.650000  90.700000 ;
      RECT 17.325000  90.400000 18.800000  90.550000 ;
      RECT 17.475000  90.250000 18.950000  90.400000 ;
      RECT 17.625000  90.100000 19.100000  90.250000 ;
      RECT 17.775000  89.950000 19.250000  90.100000 ;
      RECT 17.925000  89.800000 19.400000  89.950000 ;
      RECT 18.075000  89.650000 19.550000  89.800000 ;
      RECT 18.225000  89.500000 19.700000  89.650000 ;
      RECT 18.375000  89.350000 19.850000  89.500000 ;
      RECT 18.525000  89.200000 20.000000  89.350000 ;
      RECT 18.675000  89.050000 20.150000  89.200000 ;
      RECT 18.825000  88.900000 20.300000  89.050000 ;
      RECT 18.975000  88.750000 20.450000  88.900000 ;
      RECT 19.125000  88.600000 20.600000  88.750000 ;
      RECT 19.275000  88.450000 20.750000  88.600000 ;
      RECT 19.425000  88.300000 20.900000  88.450000 ;
      RECT 19.575000  88.150000 21.050000  88.300000 ;
      RECT 19.725000  88.000000 21.200000  88.150000 ;
      RECT 19.875000  87.850000 21.350000  88.000000 ;
      RECT 20.025000  87.700000 21.500000  87.850000 ;
      RECT 20.175000  87.550000 21.650000  87.700000 ;
      RECT 20.325000  87.400000 21.800000  87.550000 ;
      RECT 20.475000  87.250000 21.950000  87.400000 ;
      RECT 20.625000  87.100000 22.100000  87.250000 ;
      RECT 20.775000  86.950000 22.250000  87.100000 ;
      RECT 20.925000  86.800000 22.400000  86.950000 ;
      RECT 21.075000  86.650000 22.550000  86.800000 ;
      RECT 21.225000  86.500000 22.700000  86.650000 ;
      RECT 21.375000  86.350000 22.850000  86.500000 ;
      RECT 21.525000  86.200000 23.000000  86.350000 ;
      RECT 21.675000  86.050000 23.150000  86.200000 ;
      RECT 21.825000  85.900000 23.300000  86.050000 ;
      RECT 21.950000  85.775000 23.450000  85.900000 ;
      RECT 22.005000  96.955000 25.635000 166.935000 ;
      RECT 22.005000  96.955000 25.635000 166.935000 ;
      RECT 22.005000 166.935000 25.635000 170.445000 ;
      RECT 22.075000  96.885000 25.635000  96.955000 ;
      RECT 22.100000  85.625000 23.450000  85.775000 ;
      RECT 22.155000 166.935000 25.635000 167.085000 ;
      RECT 22.225000  96.735000 25.635000  96.885000 ;
      RECT 22.250000  85.475000 23.450000  85.625000 ;
      RECT 22.305000 167.085000 25.635000 167.235000 ;
      RECT 22.375000  96.585000 25.635000  96.735000 ;
      RECT 22.400000  85.325000 23.450000  85.475000 ;
      RECT 22.455000 167.235000 25.635000 167.385000 ;
      RECT 22.525000  96.435000 25.635000  96.585000 ;
      RECT 22.550000  85.175000 23.450000  85.325000 ;
      RECT 22.605000 167.385000 25.635000 167.535000 ;
      RECT 22.675000  96.285000 25.635000  96.435000 ;
      RECT 22.700000  85.025000 23.450000  85.175000 ;
      RECT 22.755000 167.535000 25.635000 167.685000 ;
      RECT 22.825000  96.135000 25.635000  96.285000 ;
      RECT 22.850000  84.875000 23.450000  85.025000 ;
      RECT 22.905000 167.685000 25.635000 167.835000 ;
      RECT 22.975000  95.985000 25.635000  96.135000 ;
      RECT 23.000000  84.725000 23.450000  84.875000 ;
      RECT 23.055000 167.835000 25.635000 167.985000 ;
      RECT 23.100000  84.485000 23.450000  85.900000 ;
      RECT 23.125000  95.835000 25.635000  95.985000 ;
      RECT 23.150000  84.575000 23.450000  84.725000 ;
      RECT 23.205000 167.985000 25.635000 168.135000 ;
      RECT 23.275000  95.685000 25.635000  95.835000 ;
      RECT 23.300000  84.425000 23.450000  84.575000 ;
      RECT 23.355000 168.135000 25.635000 168.285000 ;
      RECT 23.425000  95.535000 25.635000  95.685000 ;
      RECT 23.505000 168.285000 25.635000 168.435000 ;
      RECT 23.575000  95.385000 25.635000  95.535000 ;
      RECT 23.655000 168.435000 25.635000 168.585000 ;
      RECT 23.725000  95.235000 25.635000  95.385000 ;
      RECT 23.805000 168.585000 25.635000 168.735000 ;
      RECT 23.875000  95.085000 25.635000  95.235000 ;
      RECT 23.955000 168.735000 25.635000 168.885000 ;
      RECT 24.025000  94.935000 25.635000  95.085000 ;
      RECT 24.105000 168.885000 25.635000 169.035000 ;
      RECT 24.175000  94.785000 25.635000  94.935000 ;
      RECT 24.255000 169.035000 25.635000 169.185000 ;
      RECT 24.325000  94.635000 25.635000  94.785000 ;
      RECT 24.405000 169.185000 25.635000 169.335000 ;
      RECT 24.475000  94.485000 25.635000  94.635000 ;
      RECT 24.555000 169.335000 25.635000 169.485000 ;
      RECT 24.625000  94.335000 25.635000  94.485000 ;
      RECT 24.625000  94.335000 25.635000  96.955000 ;
      RECT 24.705000 169.485000 25.635000 169.635000 ;
      RECT 24.745000  94.215000 25.635000  94.335000 ;
      RECT 24.800000   0.000000 25.600000  82.335000 ;
      RECT 24.800000  82.335000 25.150000  82.785000 ;
      RECT 24.855000 169.635000 25.635000 169.785000 ;
      RECT 24.895000  94.065000 25.755000  94.215000 ;
      RECT 24.900000   0.000000 25.600000  82.335000 ;
      RECT 24.900000  82.335000 25.450000  82.485000 ;
      RECT 24.900000  82.485000 25.300000  82.635000 ;
      RECT 24.900000  82.635000 25.150000  82.785000 ;
      RECT 24.900000  82.785000 25.000000  82.935000 ;
      RECT 25.005000 169.785000 25.635000 169.935000 ;
      RECT 25.045000  93.915000 25.905000  94.065000 ;
      RECT 25.155000 169.935000 25.635000 170.085000 ;
      RECT 25.195000  93.765000 26.055000  93.915000 ;
      RECT 25.305000 170.085000 25.635000 170.235000 ;
      RECT 25.345000  93.615000 26.205000  93.765000 ;
      RECT 25.455000 170.235000 25.635000 170.385000 ;
      RECT 25.495000  93.465000 26.355000  93.615000 ;
      RECT 25.515000 170.445000 25.635000 189.915000 ;
      RECT 25.605000 170.385000 25.635000 170.535000 ;
      RECT 25.645000  93.315000 26.505000  93.465000 ;
      RECT 25.795000  93.165000 26.655000  93.315000 ;
      RECT 25.945000  93.015000 26.805000  93.165000 ;
      RECT 26.095000  92.865000 26.955000  93.015000 ;
      RECT 26.245000  92.715000 27.105000  92.865000 ;
      RECT 26.395000  92.565000 27.255000  92.715000 ;
      RECT 26.545000  92.415000 27.405000  92.565000 ;
      RECT 26.695000  92.265000 27.555000  92.415000 ;
      RECT 26.845000  92.115000 27.705000  92.265000 ;
      RECT 26.995000  91.965000 27.855000  92.115000 ;
      RECT 27.145000  91.815000 28.005000  91.965000 ;
      RECT 27.295000  91.665000 28.155000  91.815000 ;
      RECT 27.445000  91.515000 28.305000  91.665000 ;
      RECT 27.595000  91.365000 28.455000  91.515000 ;
      RECT 27.745000  91.215000 28.605000  91.365000 ;
      RECT 27.895000  91.065000 28.755000  91.215000 ;
      RECT 28.045000  90.915000 28.905000  91.065000 ;
      RECT 28.195000  90.765000 29.055000  90.915000 ;
      RECT 28.345000  90.615000 29.205000  90.765000 ;
      RECT 28.495000  90.465000 29.355000  90.615000 ;
      RECT 28.645000  90.315000 29.505000  90.465000 ;
      RECT 28.795000  90.165000 29.655000  90.315000 ;
      RECT 28.945000  90.015000 29.805000  90.165000 ;
      RECT 29.095000  89.865000 29.955000  90.015000 ;
      RECT 29.245000  89.715000 30.105000  89.865000 ;
      RECT 29.395000  89.565000 30.255000  89.715000 ;
      RECT 29.545000  89.415000 30.405000  89.565000 ;
      RECT 29.695000  89.265000 30.555000  89.415000 ;
      RECT 29.845000  89.115000 30.705000  89.265000 ;
      RECT 29.995000  88.965000 30.855000  89.115000 ;
      RECT 30.145000  88.815000 31.005000  88.965000 ;
      RECT 30.295000  88.665000 31.155000  88.815000 ;
      RECT 30.445000  88.515000 31.305000  88.665000 ;
      RECT 30.595000  88.365000 31.455000  88.515000 ;
      RECT 30.745000  88.215000 31.605000  88.365000 ;
      RECT 30.895000  88.065000 31.755000  88.215000 ;
      RECT 31.045000  87.915000 31.905000  88.065000 ;
      RECT 31.195000  87.765000 32.055000  87.915000 ;
      RECT 31.345000  87.615000 32.205000  87.765000 ;
      RECT 31.495000  87.465000 32.355000  87.615000 ;
      RECT 31.645000  87.315000 32.505000  87.465000 ;
      RECT 31.795000  87.165000 32.655000  87.315000 ;
      RECT 31.945000  87.015000 32.805000  87.165000 ;
      RECT 32.095000  86.865000 32.955000  87.015000 ;
      RECT 32.245000  86.715000 33.105000  86.865000 ;
      RECT 32.395000  86.565000 33.255000  86.715000 ;
      RECT 32.435000  93.555000 40.410000  93.705000 ;
      RECT 32.435000  93.555000 42.435000  95.580000 ;
      RECT 32.435000  93.705000 40.560000  93.855000 ;
      RECT 32.435000  93.855000 40.710000  94.005000 ;
      RECT 32.435000  94.005000 40.860000  94.155000 ;
      RECT 32.435000  94.155000 41.010000  94.305000 ;
      RECT 32.435000  94.305000 41.160000  94.455000 ;
      RECT 32.435000  94.455000 41.310000  94.605000 ;
      RECT 32.435000  94.605000 41.460000  94.755000 ;
      RECT 32.435000  94.755000 41.610000  94.905000 ;
      RECT 32.435000  94.905000 41.760000  95.055000 ;
      RECT 32.435000  95.055000 41.910000  95.205000 ;
      RECT 32.435000  95.205000 42.060000  95.355000 ;
      RECT 32.435000  95.355000 42.210000  95.505000 ;
      RECT 32.435000  95.505000 42.360000  95.580000 ;
      RECT 32.435000  95.580000 35.440000 159.400000 ;
      RECT 32.435000  95.580000 42.435000 162.405000 ;
      RECT 32.435000 159.400000 36.680000 162.405000 ;
      RECT 32.435000 162.405000 42.435000 163.970000 ;
      RECT 32.515000  93.475000 40.330000  93.555000 ;
      RECT 32.545000  84.855000 34.105000  85.865000 ;
      RECT 32.545000  84.855000 34.105000  85.865000 ;
      RECT 32.545000  85.865000 33.555000  86.415000 ;
      RECT 32.545000  85.865000 33.955000  86.015000 ;
      RECT 32.545000  86.015000 33.805000  86.165000 ;
      RECT 32.545000  86.165000 33.655000  86.315000 ;
      RECT 32.545000  86.315000 33.555000  86.415000 ;
      RECT 32.545000  86.415000 33.405000  86.565000 ;
      RECT 32.570000  84.830000 34.080000  84.855000 ;
      RECT 32.585000 162.405000 42.435000 162.555000 ;
      RECT 32.665000  93.325000 40.180000  93.475000 ;
      RECT 32.720000  84.680000 33.930000  84.830000 ;
      RECT 32.735000 162.555000 42.435000 162.705000 ;
      RECT 32.815000  93.175000 40.030000  93.325000 ;
      RECT 32.870000  84.530000 33.780000  84.680000 ;
      RECT 32.885000 162.705000 42.435000 162.855000 ;
      RECT 32.965000  93.025000 39.880000  93.175000 ;
      RECT 33.020000  84.380000 33.630000  84.530000 ;
      RECT 33.020000  84.380000 34.105000  84.855000 ;
      RECT 33.035000 162.855000 42.435000 163.005000 ;
      RECT 33.115000  92.875000 39.730000  93.025000 ;
      RECT 33.185000 163.005000 42.435000 163.155000 ;
      RECT 33.265000  92.725000 39.580000  92.875000 ;
      RECT 33.335000 163.155000 42.435000 163.305000 ;
      RECT 33.415000  92.575000 39.430000  92.725000 ;
      RECT 33.485000 163.305000 42.435000 163.455000 ;
      RECT 33.565000  92.425000 39.280000  92.575000 ;
      RECT 33.635000 163.455000 42.435000 163.605000 ;
      RECT 33.715000  92.275000 39.130000  92.425000 ;
      RECT 33.785000 163.605000 42.435000 163.755000 ;
      RECT 33.865000  92.125000 38.980000  92.275000 ;
      RECT 33.935000 163.755000 42.435000 163.905000 ;
      RECT 34.000000 163.905000 42.435000 163.970000 ;
      RECT 34.000000 163.970000 39.110000 167.295000 ;
      RECT 34.015000  91.975000 38.830000  92.125000 ;
      RECT 34.150000 163.970000 42.285000 164.120000 ;
      RECT 34.165000  91.825000 38.680000  91.975000 ;
      RECT 34.300000 164.120000 42.135000 164.270000 ;
      RECT 34.315000  91.675000 38.530000  91.825000 ;
      RECT 34.450000 164.270000 41.985000 164.420000 ;
      RECT 34.465000  91.525000 38.380000  91.675000 ;
      RECT 34.600000 164.420000 41.835000 164.570000 ;
      RECT 34.615000  91.375000 38.230000  91.525000 ;
      RECT 34.750000 164.570000 41.685000 164.720000 ;
      RECT 34.765000  91.225000 38.080000  91.375000 ;
      RECT 34.900000 164.720000 41.535000 164.870000 ;
      RECT 34.915000  91.075000 37.930000  91.225000 ;
      RECT 35.050000 164.870000 41.385000 165.020000 ;
      RECT 35.065000  90.925000 37.780000  91.075000 ;
      RECT 35.200000 165.020000 41.235000 165.170000 ;
      RECT 35.215000  90.775000 37.630000  90.925000 ;
      RECT 35.215000  90.775000 40.410000  93.555000 ;
      RECT 35.350000 165.170000 41.085000 165.320000 ;
      RECT 35.435000  94.800000 37.410000  94.950000 ;
      RECT 35.435000  94.800000 37.410000  94.950000 ;
      RECT 35.435000  94.950000 37.560000  95.100000 ;
      RECT 35.435000  94.950000 37.560000  95.100000 ;
      RECT 35.435000  95.100000 37.710000  95.250000 ;
      RECT 35.435000  95.100000 37.710000  95.250000 ;
      RECT 35.435000  95.250000 37.860000  95.400000 ;
      RECT 35.435000  95.250000 37.860000  95.400000 ;
      RECT 35.435000  95.400000 38.010000  95.550000 ;
      RECT 35.435000  95.400000 38.010000  95.550000 ;
      RECT 35.435000  95.550000 38.160000  95.700000 ;
      RECT 35.435000  95.550000 38.160000  95.700000 ;
      RECT 35.435000  95.700000 38.310000  95.850000 ;
      RECT 35.435000  95.700000 38.310000  95.850000 ;
      RECT 35.435000  95.850000 38.460000  96.000000 ;
      RECT 35.435000  95.850000 38.460000  96.000000 ;
      RECT 35.435000  96.000000 38.610000  96.150000 ;
      RECT 35.435000  96.000000 38.610000  96.150000 ;
      RECT 35.435000  96.150000 38.760000  96.300000 ;
      RECT 35.435000  96.150000 38.760000  96.300000 ;
      RECT 35.435000  96.300000 38.910000  96.450000 ;
      RECT 35.435000  96.300000 38.910000  96.450000 ;
      RECT 35.435000  96.450000 39.060000  96.600000 ;
      RECT 35.435000  96.450000 39.060000  96.600000 ;
      RECT 35.435000  96.600000 39.210000  96.750000 ;
      RECT 35.435000  96.600000 39.210000  96.750000 ;
      RECT 35.435000  96.750000 39.360000  96.825000 ;
      RECT 35.435000  96.750000 39.360000  96.825000 ;
      RECT 35.435000  96.825000 39.435000 161.160000 ;
      RECT 35.500000 165.320000 40.935000 165.470000 ;
      RECT 35.520000  94.715000 37.325000  94.800000 ;
      RECT 35.520000  94.715000 37.325000  94.800000 ;
      RECT 35.585000 161.160000 39.435000 161.310000 ;
      RECT 35.585000 161.160000 39.435000 161.310000 ;
      RECT 35.650000 165.470000 40.785000 165.620000 ;
      RECT 35.670000  94.565000 37.175000  94.715000 ;
      RECT 35.670000  94.565000 37.175000  94.715000 ;
      RECT 35.735000 161.310000 39.435000 161.460000 ;
      RECT 35.735000 161.310000 39.435000 161.460000 ;
      RECT 35.800000 165.620000 40.635000 165.770000 ;
      RECT 35.820000  94.415000 37.025000  94.565000 ;
      RECT 35.820000  94.415000 37.025000  94.565000 ;
      RECT 35.885000 161.460000 39.435000 161.610000 ;
      RECT 35.885000 161.460000 39.435000 161.610000 ;
      RECT 35.950000 165.770000 40.485000 165.920000 ;
      RECT 35.975000  94.265000 36.875000  94.415000 ;
      RECT 35.975000  94.265000 36.875000  94.415000 ;
      RECT 36.035000 161.610000 39.435000 161.760000 ;
      RECT 36.035000 161.610000 39.435000 161.760000 ;
      RECT 36.100000 165.920000 40.335000 166.070000 ;
      RECT 36.125000  94.115000 36.725000  94.265000 ;
      RECT 36.125000  94.115000 36.725000  94.265000 ;
      RECT 36.185000 161.760000 39.435000 161.910000 ;
      RECT 36.185000 161.760000 39.435000 161.910000 ;
      RECT 36.250000 166.070000 40.185000 166.220000 ;
      RECT 36.275000  93.965000 36.575000  94.115000 ;
      RECT 36.275000  93.965000 36.575000  94.115000 ;
      RECT 36.335000 161.910000 39.435000 162.060000 ;
      RECT 36.335000 161.910000 39.435000 162.060000 ;
      RECT 36.400000 166.220000 40.035000 166.370000 ;
      RECT 36.485000 162.060000 39.435000 162.210000 ;
      RECT 36.485000 162.060000 39.435000 162.210000 ;
      RECT 36.550000 166.370000 39.885000 166.520000 ;
      RECT 36.635000 162.210000 39.435000 162.360000 ;
      RECT 36.635000 162.210000 39.435000 162.360000 ;
      RECT 36.700000 166.520000 39.735000 166.670000 ;
      RECT 36.785000 162.360000 39.435000 162.510000 ;
      RECT 36.785000 162.360000 39.435000 162.510000 ;
      RECT 36.850000 166.670000 39.585000 166.820000 ;
      RECT 36.935000 162.510000 39.435000 162.660000 ;
      RECT 36.935000 162.510000 39.435000 162.660000 ;
      RECT 37.000000 162.660000 39.435000 162.725000 ;
      RECT 37.000000 162.660000 39.435000 162.725000 ;
      RECT 37.000000 166.820000 39.435000 166.970000 ;
      RECT 37.150000 162.725000 39.285000 162.875000 ;
      RECT 37.150000 162.725000 39.285000 162.875000 ;
      RECT 37.150000 166.970000 39.285000 167.120000 ;
      RECT 37.280000   0.000000 37.980000  69.890000 ;
      RECT 37.280000   0.000000 37.980000  69.890000 ;
      RECT 37.280000  69.890000 50.355000  70.940000 ;
      RECT 37.280000  69.890000 50.355000  74.340000 ;
      RECT 37.280000  69.890000 50.455000  70.940000 ;
      RECT 37.280000  70.940000 50.455000  74.340000 ;
      RECT 37.300000 162.875000 39.135000 163.025000 ;
      RECT 37.300000 162.875000 39.135000 163.025000 ;
      RECT 37.300000 167.120000 39.135000 167.270000 ;
      RECT 37.325000 167.270000 39.110000 167.295000 ;
      RECT 37.325000 167.295000 37.545000 168.860000 ;
      RECT 37.325000 167.295000 38.960000 167.445000 ;
      RECT 37.325000 167.445000 38.810000 167.595000 ;
      RECT 37.325000 167.595000 38.660000 167.745000 ;
      RECT 37.325000 167.745000 38.510000 167.895000 ;
      RECT 37.325000 167.895000 38.360000 168.045000 ;
      RECT 37.325000 168.045000 38.210000 168.195000 ;
      RECT 37.325000 168.195000 38.060000 168.345000 ;
      RECT 37.325000 168.345000 37.910000 168.495000 ;
      RECT 37.325000 168.495000 37.760000 168.645000 ;
      RECT 37.325000 168.645000 37.610000 168.795000 ;
      RECT 37.325000 168.795000 37.460000 168.945000 ;
      RECT 37.325000 168.860000 37.545000 189.915000 ;
      RECT 37.430000  70.940000 50.355000  71.090000 ;
      RECT 37.430000  70.940000 50.355000  71.090000 ;
      RECT 37.450000 163.025000 38.985000 163.175000 ;
      RECT 37.450000 163.025000 38.985000 163.175000 ;
      RECT 37.580000  71.090000 50.355000  71.240000 ;
      RECT 37.580000  71.090000 50.355000  71.240000 ;
      RECT 37.600000 163.175000 38.835000 163.325000 ;
      RECT 37.600000 163.175000 38.835000 163.325000 ;
      RECT 37.730000  71.240000 50.355000  71.390000 ;
      RECT 37.730000  71.240000 50.355000  71.390000 ;
      RECT 37.750000 163.325000 38.685000 163.475000 ;
      RECT 37.750000 163.325000 38.685000 163.475000 ;
      RECT 37.880000  71.390000 50.355000  71.540000 ;
      RECT 37.880000  71.390000 50.355000  71.540000 ;
      RECT 37.900000 163.475000 38.535000 163.625000 ;
      RECT 37.900000 163.475000 38.535000 163.625000 ;
      RECT 38.030000  71.540000 50.355000  71.690000 ;
      RECT 38.030000  71.540000 50.355000  71.690000 ;
      RECT 38.050000 163.625000 38.385000 163.775000 ;
      RECT 38.050000 163.625000 38.385000 163.775000 ;
      RECT 38.180000  71.690000 50.355000  71.840000 ;
      RECT 38.180000  71.690000 50.355000  71.840000 ;
      RECT 38.190000  95.580000 42.435000  98.585000 ;
      RECT 38.200000 163.775000 38.235000 163.925000 ;
      RECT 38.200000 163.775000 38.235000 163.925000 ;
      RECT 38.215000 163.925000 38.220000 163.940000 ;
      RECT 38.215000 163.925000 38.220000 163.940000 ;
      RECT 38.330000  71.840000 50.355000  71.990000 ;
      RECT 38.330000  71.840000 50.355000  71.990000 ;
      RECT 38.480000  71.990000 50.355000  72.140000 ;
      RECT 38.480000  71.990000 50.355000  72.140000 ;
      RECT 38.630000  72.140000 50.355000  72.290000 ;
      RECT 38.630000  72.140000 50.355000  72.290000 ;
      RECT 38.780000  72.290000 50.355000  72.440000 ;
      RECT 38.780000  72.290000 50.355000  72.440000 ;
      RECT 38.930000  72.440000 50.355000  72.590000 ;
      RECT 38.930000  72.440000 50.355000  72.590000 ;
      RECT 39.080000  72.590000 50.355000  72.740000 ;
      RECT 39.080000  72.590000 50.355000  72.740000 ;
      RECT 39.230000  72.740000 50.355000  72.890000 ;
      RECT 39.230000  72.740000 50.355000  72.890000 ;
      RECT 39.380000  72.890000 50.355000  73.040000 ;
      RECT 39.380000  72.890000 50.355000  73.040000 ;
      RECT 39.430000  98.585000 42.435000 162.405000 ;
      RECT 39.530000  73.040000 50.355000  73.190000 ;
      RECT 39.530000  73.040000 50.355000  73.190000 ;
      RECT 39.680000  73.190000 50.355000  73.340000 ;
      RECT 39.680000  73.190000 50.355000  73.340000 ;
      RECT 39.785000  84.855000 41.210000  87.195000 ;
      RECT 39.785000  84.855000 41.210000  87.195000 ;
      RECT 39.785000  87.195000 41.210000  87.610000 ;
      RECT 39.810000  84.830000 41.185000  84.855000 ;
      RECT 39.830000  73.340000 50.355000  73.490000 ;
      RECT 39.830000  73.340000 50.355000  73.490000 ;
      RECT 39.935000  87.195000 41.210000  87.345000 ;
      RECT 39.960000  84.680000 41.035000  84.830000 ;
      RECT 39.980000  73.490000 50.355000  73.640000 ;
      RECT 39.980000  73.490000 50.355000  73.640000 ;
      RECT 40.085000  87.345000 41.210000  87.495000 ;
      RECT 40.110000  84.530000 40.885000  84.680000 ;
      RECT 40.130000  73.640000 50.355000  73.790000 ;
      RECT 40.130000  73.640000 50.355000  73.790000 ;
      RECT 40.200000  87.495000 41.210000  87.610000 ;
      RECT 40.200000  87.610000 50.245000  96.645000 ;
      RECT 40.260000  84.380000 40.735000  84.530000 ;
      RECT 40.260000  84.380000 41.210000  84.855000 ;
      RECT 40.280000  73.790000 50.355000  73.940000 ;
      RECT 40.280000  73.790000 50.355000  73.940000 ;
      RECT 40.350000  87.610000 41.210000  87.760000 ;
      RECT 40.430000  73.940000 50.355000  74.090000 ;
      RECT 40.430000  73.940000 50.355000  74.090000 ;
      RECT 40.500000  87.760000 41.360000  87.910000 ;
      RECT 40.580000  74.090000 50.355000  74.240000 ;
      RECT 40.580000  74.090000 50.355000  74.240000 ;
      RECT 40.650000  87.910000 41.510000  88.060000 ;
      RECT 40.680000  74.240000 50.355000  74.340000 ;
      RECT 40.680000  74.240000 50.355000  74.340000 ;
      RECT 40.800000  88.060000 41.660000  88.210000 ;
      RECT 40.950000  88.210000 41.810000  88.360000 ;
      RECT 41.100000  88.360000 41.960000  88.510000 ;
      RECT 41.250000  88.510000 42.110000  88.660000 ;
      RECT 41.400000  88.660000 42.260000  88.810000 ;
      RECT 41.550000  88.810000 42.410000  88.960000 ;
      RECT 41.700000  88.960000 42.560000  89.110000 ;
      RECT 41.850000  89.110000 42.710000  89.260000 ;
      RECT 42.000000  89.260000 42.860000  89.410000 ;
      RECT 42.150000  89.410000 43.010000  89.560000 ;
      RECT 42.300000  89.560000 43.160000  89.710000 ;
      RECT 42.450000  89.710000 43.310000  89.860000 ;
      RECT 42.600000  89.860000 43.460000  90.010000 ;
      RECT 42.750000  90.010000 43.610000  90.160000 ;
      RECT 42.900000  90.160000 43.760000  90.310000 ;
      RECT 43.050000  90.310000 43.910000  90.460000 ;
      RECT 43.200000  90.460000 44.060000  90.610000 ;
      RECT 43.350000  90.610000 44.210000  90.760000 ;
      RECT 43.500000  90.760000 44.360000  90.910000 ;
      RECT 43.650000  90.910000 44.510000  91.060000 ;
      RECT 43.800000  91.060000 44.660000  91.210000 ;
      RECT 43.950000  91.210000 44.810000  91.360000 ;
      RECT 44.100000  91.360000 44.960000  91.510000 ;
      RECT 44.250000  91.510000 45.110000  91.660000 ;
      RECT 44.400000  91.660000 45.260000  91.810000 ;
      RECT 44.550000  91.810000 45.410000  91.960000 ;
      RECT 44.700000  91.960000 45.560000  92.110000 ;
      RECT 44.850000  92.110000 45.710000  92.260000 ;
      RECT 45.000000  92.260000 45.860000  92.410000 ;
      RECT 45.150000  92.410000 46.010000  92.560000 ;
      RECT 45.300000  92.560000 46.160000  92.710000 ;
      RECT 45.450000  92.710000 46.310000  92.860000 ;
      RECT 45.600000  92.860000 46.460000  93.010000 ;
      RECT 45.750000  93.010000 46.610000  93.160000 ;
      RECT 45.900000  93.160000 46.760000  93.310000 ;
      RECT 46.050000  93.310000 46.910000  93.460000 ;
      RECT 46.200000  93.460000 47.060000  93.610000 ;
      RECT 46.350000  93.610000 47.210000  93.760000 ;
      RECT 46.500000  93.760000 47.360000  93.910000 ;
      RECT 46.650000  93.910000 47.510000  94.060000 ;
      RECT 46.800000  94.060000 47.660000  94.210000 ;
      RECT 46.950000  94.210000 47.810000  94.360000 ;
      RECT 46.960000  74.340000 50.455000  76.650000 ;
      RECT 47.100000  94.360000 47.960000  94.510000 ;
      RECT 47.110000  74.340000 50.355000  74.490000 ;
      RECT 47.110000  74.340000 50.355000  74.490000 ;
      RECT 47.250000  94.510000 48.110000  94.660000 ;
      RECT 47.260000  74.490000 50.355000  74.640000 ;
      RECT 47.260000  74.490000 50.355000  74.640000 ;
      RECT 47.400000  94.660000 48.260000  94.810000 ;
      RECT 47.410000  74.640000 50.355000  74.790000 ;
      RECT 47.410000  74.640000 50.355000  74.790000 ;
      RECT 47.550000  94.810000 48.410000  94.960000 ;
      RECT 47.560000  74.790000 50.355000  74.940000 ;
      RECT 47.560000  74.790000 50.355000  74.940000 ;
      RECT 47.700000  94.960000 48.560000  95.110000 ;
      RECT 47.710000  74.940000 50.355000  75.090000 ;
      RECT 47.710000  74.940000 50.355000  75.090000 ;
      RECT 47.850000  95.110000 48.710000  95.260000 ;
      RECT 47.860000  75.090000 50.355000  75.240000 ;
      RECT 47.860000  75.090000 50.355000  75.240000 ;
      RECT 48.000000  95.260000 48.860000  95.410000 ;
      RECT 48.010000  75.240000 50.355000  75.390000 ;
      RECT 48.010000  75.240000 50.355000  75.390000 ;
      RECT 48.150000  95.410000 49.010000  95.560000 ;
      RECT 48.160000  75.390000 50.355000  75.540000 ;
      RECT 48.160000  75.390000 50.355000  75.540000 ;
      RECT 48.300000  95.560000 49.160000  95.710000 ;
      RECT 48.310000  75.540000 50.355000  75.690000 ;
      RECT 48.310000  75.540000 50.355000  75.690000 ;
      RECT 48.450000  95.710000 49.310000  95.860000 ;
      RECT 48.460000  75.690000 50.355000  75.840000 ;
      RECT 48.460000  75.690000 50.355000  75.840000 ;
      RECT 48.600000  95.860000 49.460000  96.010000 ;
      RECT 48.610000  75.840000 50.355000  75.990000 ;
      RECT 48.610000  75.840000 50.355000  75.990000 ;
      RECT 48.750000  96.010000 49.610000  96.160000 ;
      RECT 48.760000  75.990000 50.355000  76.140000 ;
      RECT 48.760000  75.990000 50.355000  76.140000 ;
      RECT 48.900000  96.160000 49.760000  96.310000 ;
      RECT 48.910000  76.140000 50.355000  76.290000 ;
      RECT 48.910000  76.140000 50.355000  76.290000 ;
      RECT 49.050000  96.310000 49.910000  96.460000 ;
      RECT 49.060000  76.290000 50.355000  76.440000 ;
      RECT 49.060000  76.290000 50.355000  76.440000 ;
      RECT 49.200000  96.460000 50.060000  96.610000 ;
      RECT 49.210000  76.440000 50.355000  76.590000 ;
      RECT 49.210000  76.440000 50.355000  76.590000 ;
      RECT 49.235000  96.610000 50.210000  96.645000 ;
      RECT 49.235000  96.645000 50.245000  96.795000 ;
      RECT 49.235000  96.645000 53.930000 100.330000 ;
      RECT 49.235000  96.795000 50.395000  96.945000 ;
      RECT 49.235000  96.945000 50.545000  97.095000 ;
      RECT 49.235000  97.095000 50.695000  97.245000 ;
      RECT 49.235000  97.245000 50.845000  97.395000 ;
      RECT 49.235000  97.395000 50.995000  97.545000 ;
      RECT 49.235000  97.545000 51.145000  97.695000 ;
      RECT 49.235000  97.695000 51.295000  97.845000 ;
      RECT 49.235000  97.845000 51.445000  97.995000 ;
      RECT 49.235000  97.995000 51.595000  98.145000 ;
      RECT 49.235000  98.145000 51.745000  98.295000 ;
      RECT 49.235000  98.295000 51.895000  98.445000 ;
      RECT 49.235000  98.445000 52.045000  98.595000 ;
      RECT 49.235000  98.595000 52.195000  98.745000 ;
      RECT 49.235000  98.745000 52.345000  98.895000 ;
      RECT 49.235000  98.895000 52.495000  99.045000 ;
      RECT 49.235000  99.045000 52.645000  99.195000 ;
      RECT 49.235000  99.195000 52.795000  99.345000 ;
      RECT 49.235000  99.345000 52.945000  99.495000 ;
      RECT 49.235000  99.495000 53.095000  99.645000 ;
      RECT 49.235000  99.645000 53.245000  99.795000 ;
      RECT 49.235000  99.795000 53.395000  99.945000 ;
      RECT 49.235000  99.945000 53.545000 100.095000 ;
      RECT 49.235000 100.095000 53.695000 100.245000 ;
      RECT 49.235000 100.245000 53.845000 100.330000 ;
      RECT 49.235000 100.330000 53.930000 164.295000 ;
      RECT 49.235000 100.330000 53.930000 164.295000 ;
      RECT 49.235000 164.295000 49.470000 168.755000 ;
      RECT 49.235000 164.295000 53.780000 164.445000 ;
      RECT 49.235000 164.445000 53.630000 164.595000 ;
      RECT 49.235000 164.595000 53.480000 164.745000 ;
      RECT 49.235000 164.745000 53.330000 164.895000 ;
      RECT 49.235000 164.895000 53.180000 165.045000 ;
      RECT 49.235000 165.045000 53.030000 165.195000 ;
      RECT 49.235000 165.195000 52.880000 165.345000 ;
      RECT 49.235000 165.345000 52.730000 165.495000 ;
      RECT 49.235000 165.495000 52.580000 165.645000 ;
      RECT 49.235000 165.645000 52.430000 165.795000 ;
      RECT 49.235000 165.795000 52.280000 165.945000 ;
      RECT 49.235000 165.945000 52.130000 166.095000 ;
      RECT 49.235000 166.095000 51.980000 166.245000 ;
      RECT 49.235000 166.245000 51.830000 166.395000 ;
      RECT 49.235000 166.395000 51.680000 166.545000 ;
      RECT 49.235000 166.545000 51.530000 166.695000 ;
      RECT 49.235000 166.695000 51.380000 166.845000 ;
      RECT 49.235000 166.845000 51.230000 166.995000 ;
      RECT 49.235000 166.995000 51.080000 167.145000 ;
      RECT 49.235000 167.145000 50.930000 167.295000 ;
      RECT 49.235000 167.295000 50.780000 167.445000 ;
      RECT 49.235000 167.445000 50.630000 167.595000 ;
      RECT 49.235000 167.595000 50.480000 167.745000 ;
      RECT 49.235000 167.745000 50.330000 167.895000 ;
      RECT 49.235000 167.895000 50.180000 168.045000 ;
      RECT 49.235000 168.045000 50.030000 168.195000 ;
      RECT 49.235000 168.195000 49.880000 168.345000 ;
      RECT 49.235000 168.345000 49.730000 168.495000 ;
      RECT 49.235000 168.495000 49.580000 168.645000 ;
      RECT 49.235000 168.645000 49.430000 168.795000 ;
      RECT 49.235000 168.755000 49.470000 189.915000 ;
      RECT 49.235000 168.795000 49.280000 168.945000 ;
      RECT 49.270000  76.590000 50.355000  76.650000 ;
      RECT 49.270000  76.590000 50.355000  76.650000 ;
      RECT 49.270000  76.650000 50.455000  84.590000 ;
      RECT 49.270000  77.735000 50.355000  84.630000 ;
      RECT 49.270000  84.590000 50.510000  84.645000 ;
      RECT 49.270000  84.630000 50.355000  84.635000 ;
      RECT 49.270000  84.635000 50.360000  84.640000 ;
      RECT 49.270000  84.640000 50.365000  84.645000 ;
      RECT 49.270000  84.645000 52.660000  86.795000 ;
      RECT 49.420000  76.650000 50.355000  76.800000 ;
      RECT 49.420000  76.650000 50.355000  76.800000 ;
      RECT 49.420000  84.645000 50.370000  84.795000 ;
      RECT 49.570000  76.800000 50.355000  76.950000 ;
      RECT 49.570000  76.800000 50.355000  76.950000 ;
      RECT 49.570000  84.795000 50.520000  84.945000 ;
      RECT 49.655000   0.000000 50.355000  69.890000 ;
      RECT 49.655000   0.000000 50.455000  69.890000 ;
      RECT 49.720000  76.950000 50.355000  77.100000 ;
      RECT 49.720000  76.950000 50.355000  77.100000 ;
      RECT 49.720000  84.945000 50.670000  85.095000 ;
      RECT 49.870000  77.100000 50.355000  77.250000 ;
      RECT 49.870000  77.100000 50.355000  77.250000 ;
      RECT 49.870000  85.095000 50.820000  85.245000 ;
      RECT 50.020000  77.250000 50.355000  77.400000 ;
      RECT 50.020000  77.250000 50.355000  77.400000 ;
      RECT 50.020000  85.245000 50.970000  85.395000 ;
      RECT 50.170000  77.400000 50.355000  77.550000 ;
      RECT 50.170000  77.400000 50.355000  77.550000 ;
      RECT 50.170000  85.395000 51.120000  85.545000 ;
      RECT 50.320000  77.550000 50.355000  77.700000 ;
      RECT 50.320000  77.550000 50.355000  77.700000 ;
      RECT 50.320000  85.545000 51.270000  85.695000 ;
      RECT 50.470000  85.695000 51.420000  85.845000 ;
      RECT 50.620000  85.845000 51.570000  85.995000 ;
      RECT 50.770000  85.995000 51.720000  86.145000 ;
      RECT 50.920000  86.145000 51.870000  86.295000 ;
      RECT 51.070000  86.295000 52.020000  86.445000 ;
      RECT 51.220000  86.445000 52.170000  86.595000 ;
      RECT 51.370000  86.595000 52.320000  86.745000 ;
      RECT 51.420000  86.745000 52.470000  86.795000 ;
      RECT 51.420000  86.795000 52.520000  86.945000 ;
      RECT 51.420000  86.795000 54.075000  88.210000 ;
      RECT 51.420000  86.945000 52.670000  87.095000 ;
      RECT 51.420000  87.095000 52.820000  87.245000 ;
      RECT 51.420000  87.245000 52.970000  87.395000 ;
      RECT 51.420000  87.395000 53.120000  87.545000 ;
      RECT 51.420000  87.545000 53.270000  87.695000 ;
      RECT 51.420000  87.695000 53.420000  87.845000 ;
      RECT 51.420000  87.845000 53.570000  87.995000 ;
      RECT 51.420000  87.995000 53.720000  88.145000 ;
      RECT 51.420000  88.145000 53.870000  88.210000 ;
      RECT 51.420000  88.210000 61.745000  95.880000 ;
      RECT 51.570000  88.210000 53.935000  88.360000 ;
      RECT 51.720000  88.360000 54.085000  88.510000 ;
      RECT 51.870000  88.510000 54.235000  88.660000 ;
      RECT 52.020000  88.660000 54.385000  88.810000 ;
      RECT 52.170000  88.810000 54.535000  88.960000 ;
      RECT 52.320000  88.960000 54.685000  89.110000 ;
      RECT 52.470000  89.110000 54.835000  89.260000 ;
      RECT 52.620000  89.260000 54.985000  89.410000 ;
      RECT 52.770000  89.410000 55.135000  89.560000 ;
      RECT 52.920000  89.560000 55.285000  89.710000 ;
      RECT 53.070000  89.710000 55.435000  89.860000 ;
      RECT 53.220000  89.860000 55.585000  90.010000 ;
      RECT 53.370000  90.010000 55.735000  90.160000 ;
      RECT 53.520000  90.160000 55.885000  90.310000 ;
      RECT 53.670000  90.310000 56.035000  90.460000 ;
      RECT 53.820000  90.460000 56.185000  90.610000 ;
      RECT 53.970000  90.610000 56.335000  90.760000 ;
      RECT 54.120000  90.760000 56.485000  90.910000 ;
      RECT 54.270000  90.910000 56.635000  91.060000 ;
      RECT 54.420000  91.060000 56.785000  91.210000 ;
      RECT 54.570000  91.210000 56.935000  91.360000 ;
      RECT 54.720000  91.360000 57.085000  91.510000 ;
      RECT 54.870000  91.510000 57.235000  91.660000 ;
      RECT 55.020000  91.660000 57.385000  91.810000 ;
      RECT 55.170000  91.810000 57.535000  91.960000 ;
      RECT 55.320000  91.960000 57.685000  92.110000 ;
      RECT 55.470000  92.110000 57.835000  92.260000 ;
      RECT 55.620000  92.260000 57.985000  92.410000 ;
      RECT 55.770000  92.410000 58.135000  92.560000 ;
      RECT 55.920000  92.560000 58.285000  92.710000 ;
      RECT 56.070000  92.710000 58.435000  92.860000 ;
      RECT 56.220000  92.860000 58.585000  93.010000 ;
      RECT 56.370000  93.010000 58.735000  93.160000 ;
      RECT 56.520000  93.160000 58.885000  93.310000 ;
      RECT 56.670000  93.310000 59.035000  93.460000 ;
      RECT 56.820000  93.460000 59.185000  93.610000 ;
      RECT 56.970000  93.610000 59.335000  93.760000 ;
      RECT 57.120000  93.760000 59.485000  93.910000 ;
      RECT 57.270000  93.910000 59.635000  94.060000 ;
      RECT 57.420000  94.060000 59.785000  94.210000 ;
      RECT 57.570000  94.210000 59.935000  94.360000 ;
      RECT 57.720000  94.360000 60.085000  94.510000 ;
      RECT 57.870000  94.510000 60.235000  94.660000 ;
      RECT 58.020000  94.660000 60.385000  94.810000 ;
      RECT 58.170000  94.810000 60.535000  94.960000 ;
      RECT 58.320000  94.960000 60.685000  95.110000 ;
      RECT 58.470000  95.110000 60.835000  95.260000 ;
      RECT 58.620000  95.260000 60.985000  95.410000 ;
      RECT 58.770000  95.410000 61.135000  95.560000 ;
      RECT 58.920000  95.560000 61.285000  95.710000 ;
      RECT 59.070000  95.710000 61.435000  95.860000 ;
      RECT 59.090000  95.880000 61.745000  97.520000 ;
      RECT 59.130000  95.860000 61.585000  95.920000 ;
      RECT 59.280000  95.920000 61.645000  96.070000 ;
      RECT 59.430000  96.070000 61.645000  96.220000 ;
      RECT 59.580000  96.220000 61.645000  96.370000 ;
      RECT 59.730000  96.370000 61.645000  96.520000 ;
      RECT 59.880000  96.520000 61.645000  96.670000 ;
      RECT 60.030000  96.670000 61.645000  96.820000 ;
      RECT 60.180000  96.820000 61.645000  96.970000 ;
      RECT 60.330000  96.970000 61.645000  97.120000 ;
      RECT 60.480000  97.120000 61.645000  97.270000 ;
      RECT 60.630000  97.270000 61.645000  97.420000 ;
      RECT 60.730000  97.420000 61.645000  97.520000 ;
      RECT 60.730000  97.520000 61.645000 172.635000 ;
      RECT 60.730000  97.520000 61.745000 172.535000 ;
      RECT 60.730000 172.535000 75.000000 189.915000 ;
      RECT 60.730000 172.635000 75.000000 189.915000 ;
      RECT 60.730000 172.635000 75.000000 198.000000 ;
    LAYER met4 ;
      RECT  4.820000 102.300000  7.470000 164.545000 ;
      RECT  5.440000 101.650000  5.945000 102.180000 ;
      RECT  5.440000 164.605000  5.945000 165.135000 ;
      RECT  6.070000 101.090000  8.445000 102.160000 ;
      RECT  6.070000 164.625000  8.445000 165.695000 ;
      RECT  6.555000 100.535000  7.060000 101.065000 ;
      RECT  6.555000 165.720000  7.060000 166.250000 ;
      RECT  7.350000  99.950000  9.725000 101.020000 ;
      RECT  7.350000 165.765000  9.725000 166.835000 ;
      RECT  7.535000 102.245000  8.040000 102.775000 ;
      RECT  7.535000 164.010000  8.040000 164.540000 ;
      RECT  7.750000  99.340000  8.255000  99.870000 ;
      RECT  7.750000 166.915000  8.255000 167.445000 ;
      RECT  8.340000  98.810000 10.715000  99.880000 ;
      RECT  8.415000 166.915000 10.700000 167.865000 ;
      RECT  8.650000 101.130000  9.155000 101.660000 ;
      RECT  8.650000 165.125000  9.155000 165.655000 ;
      RECT  8.825000  98.265000  9.330000  98.795000 ;
      RECT  8.825000 167.990000  9.330000 168.520000 ;
      RECT  9.460000  97.645000 11.835000  98.715000 ;
      RECT  9.460000 168.025000 11.835000 169.095000 ;
      RECT  9.845000  99.935000 10.350000 100.465000 ;
      RECT  9.845000 166.320000 10.350000 166.850000 ;
      RECT  9.985000  97.070000 10.490000  97.600000 ;
      RECT  9.985000 169.150000 10.490000 169.680000 ;
      RECT 10.595000  96.475000 11.850000  96.480000 ;
      RECT 10.595000  96.480000 11.835000  97.545000 ;
      RECT 10.610000 169.340000 11.745000 170.260000 ;
      RECT 10.920000  98.860000 11.425000  99.390000 ;
      RECT 10.920000 167.395000 11.425000 167.925000 ;
      RECT 11.095000  95.950000 11.850000  96.475000 ;
      RECT 11.095000 170.260000 11.850000 170.790000 ;
      RECT 11.965000  95.795000 12.835000  98.295000 ;
      RECT 11.965000 168.490000 12.835000 170.990000 ;
      RECT 25.035000  17.815000 25.465000  22.250000 ;
      RECT 25.035000  39.785000 25.365000  41.435000 ;
      RECT 62.225000  95.795000 63.095000  98.295000 ;
      RECT 62.225000 168.490000 63.095000 170.990000 ;
      RECT 63.225000  96.475000 64.465000  97.545000 ;
      RECT 63.225000  97.645000 65.600000  98.715000 ;
      RECT 63.225000 169.160000 64.465000 170.230000 ;
      RECT 63.235000 168.165000 65.495000 169.005000 ;
      RECT 63.635000  98.860000 64.140000  99.390000 ;
      RECT 63.635000 167.395000 64.140000 167.925000 ;
      RECT 64.345000  98.810000 66.720000  99.880000 ;
      RECT 64.345000 166.905000 66.720000 167.975000 ;
      RECT 64.570000  97.070000 65.075000  97.600000 ;
      RECT 64.570000 169.150000 65.075000 169.680000 ;
      RECT 64.710000  99.935000 65.215000 100.465000 ;
      RECT 64.710000 166.320000 65.215000 166.850000 ;
      RECT 65.335000  99.950000 67.710000 101.020000 ;
      RECT 65.335000 165.765000 67.710000 166.835000 ;
      RECT 65.730000  98.265000 66.235000  98.795000 ;
      RECT 65.730000 167.990000 66.235000 168.520000 ;
      RECT 65.905000 101.130000 66.410000 101.660000 ;
      RECT 65.905000 165.125000 66.410000 165.655000 ;
      RECT 66.615000 101.090000 68.990000 102.160000 ;
      RECT 66.615000 164.625000 68.990000 165.695000 ;
      RECT 66.805000  99.340000 67.310000  99.870000 ;
      RECT 66.805000 166.915000 67.310000 167.445000 ;
      RECT 67.020000 102.245000 70.110000 102.775000 ;
      RECT 67.020000 164.010000 70.165000 164.350000 ;
      RECT 67.020000 164.350000 67.525000 164.540000 ;
      RECT 67.515000 103.000000 70.165000 164.010000 ;
      RECT 68.000000 100.535000 68.505000 101.065000 ;
      RECT 68.000000 165.720000 68.505000 166.250000 ;
      RECT 69.115000 101.650000 69.620000 102.180000 ;
      RECT 69.115000 164.605000 69.620000 165.135000 ;
  END
END sky130_fd_io__top_ground_lvc_wpad


MACRO sky130_fd_io__top_gpio_ovtv2
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 140 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  215.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 53.125000 140.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  215.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 48.365000 140.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN ANALOG_EN
    ANTENNAPARTIALCUTAREA  0.320000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 7.930000 14.070000 8.710000 14.390000 ;
        RECT 7.935000 14.065000 8.705000 14.070000 ;
        RECT 8.025000 13.975000 8.615000 14.065000 ;
        RECT 8.115000  0.000000 8.445000 13.805000 ;
        RECT 8.115000 13.805000 8.445000 13.845000 ;
        RECT 8.115000 13.845000 8.485000 13.885000 ;
        RECT 8.115000 13.885000 8.525000 13.975000 ;
    END
  END ANALOG_EN
  PIN ANALOG_POL
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.785000 1.165000 65.565000 1.485000 ;
        RECT 65.110000 1.040000 65.565000 1.165000 ;
        RECT 65.235000 0.000000 65.565000 0.915000 ;
        RECT 65.235000 0.915000 65.565000 1.040000 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 51.655000 0.000000 51.985000 7.760000 ;
        RECT 51.655000 7.760000 51.985000 7.910000 ;
        RECT 51.655000 7.910000 52.135000 8.060000 ;
        RECT 51.655000 8.060000 52.435000 8.380000 ;
    END
  END ANALOG_SEL
  PIN DM[0]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.105000 20.955000 129.435000 21.685000 ;
        RECT 129.125000  0.000000 129.455000 20.955000 ;
    END
  END DM[0]
  PIN DM[1]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.275000  0.000000 128.605000 19.875000 ;
        RECT 128.275000 19.875000 128.605000 19.885000 ;
        RECT 128.275000 19.885000 128.615000 19.895000 ;
        RECT 128.275000 19.895000 128.625000 20.180000 ;
        RECT 128.285000 20.180000 128.625000 20.190000 ;
        RECT 128.295000 20.190000 128.625000 20.200000 ;
        RECT 128.295000 20.200000 128.625000 21.685000 ;
    END
  END DM[1]
  PIN DM[2]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.375000 20.280000 108.725000 20.640000 ;
        RECT 108.375000 20.640000 108.705000 21.685000 ;
        RECT 108.395000  0.000000 108.725000 20.280000 ;
    END
  END DM[2]
  PIN ENABLE_H
    ANTENNAGATEAREA  8.880000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.135000  0.000000 22.465000 31.675000 ;
        RECT 22.135000 31.675000 22.465000 31.810000 ;
        RECT 22.135000 31.810000 22.600000 31.945000 ;
        RECT 22.135000 31.945000 22.875000 32.275000 ;
    END
  END ENABLE_H
  PIN ENABLE_INP_H
    ANTENNAGATEAREA  3.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 7.110000 0.000000 7.440000 19.735000 ;
    END
  END ENABLE_INP_H
  PIN ENABLE_VDDA_H
    ANTENNAGATEAREA  3.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.770000 0.000000 9.100000 8.620000 ;
    END
  END ENABLE_VDDA_H
  PIN ENABLE_VDDIO
    ANTENNAGATEAREA  6.620000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 95.845000 0.000000 96.215000 1.740000 ;
    END
  END ENABLE_VDDIO
  PIN ENABLE_VSWITCH_H
    ANTENNAGATEAREA  3.120000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.765000 0.000000 6.365000 13.205000 ;
    END
  END ENABLE_VSWITCH_H
  PIN HLD_H_N
    ANTENNAGATEAREA  1.620000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 19.635000  0.000000 19.965000 17.750000 ;
        RECT 19.635000 17.750000 19.965000 17.865000 ;
        RECT 19.635000 17.865000 20.080000 17.980000 ;
        RECT 19.635000 17.980000 20.195000 17.985000 ;
        RECT 19.675000 17.985000 20.200000 18.025000 ;
        RECT 19.715000 18.025000 20.240000 18.065000 ;
        RECT 19.830000 18.065000 20.280000 18.180000 ;
        RECT 19.945000 18.180000 20.280000 18.295000 ;
        RECT 19.950000 18.295000 20.280000 18.300000 ;
        RECT 19.950000 18.300000 20.280000 22.865000 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.900000 14.055000 27.680000 14.375000 ;
        RECT 26.905000 14.050000 27.685000 14.055000 ;
        RECT 27.055000 13.900000 27.685000 14.050000 ;
        RECT 27.205000 13.750000 27.685000 13.900000 ;
        RECT 27.355000  0.000000 27.685000 13.600000 ;
        RECT 27.355000 13.600000 27.685000 13.750000 ;
    END
  END HLD_OVR
  PIN HYS_TRIM
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.905000 8.060000 45.685000 8.380000 ;
        RECT 45.055000 7.910000 45.685000 8.060000 ;
        RECT 45.205000 7.760000 45.685000 7.910000 ;
        RECT 45.355000 0.000000 45.685000 7.610000 ;
        RECT 45.355000 7.610000 45.685000 7.760000 ;
    END
  END HYS_TRIM
  PIN IB_MODE_SEL[0]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.815000 0.000000 87.145000 21.685000 ;
    END
  END IB_MODE_SEL[0]
  PIN IB_MODE_SEL[1]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.935000 0.000000 67.265000 21.685000 ;
    END
  END IB_MODE_SEL[1]
  PIN IN
    ANTENNAPARTIALMETALSIDEAREA  23.36800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.380000 0.000000 20.710000 15.275000 ;
    END
  END IN
  PIN INP_DIS
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.095000 8.060000 107.875000 8.380000 ;
        RECT 107.285000 8.055000 107.875000 8.060000 ;
        RECT 107.415000 7.925000 107.875000 8.055000 ;
        RECT 107.545000 0.000000 107.875000 7.795000 ;
        RECT 107.545000 7.795000 107.875000 7.925000 ;
    END
  END INP_DIS
  PIN IN_H
    ANTENNAPARTIALMETALSIDEAREA  1.722440 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 23.490000 0.610000 24.710000 0.940000 ;
        RECT 24.100000 0.605000 24.710000 0.610000 ;
        RECT 24.240000 0.465000 24.710000 0.605000 ;
        RECT 24.380000 0.000000 24.710000 0.325000 ;
        RECT 24.380000 0.325000 24.710000 0.465000 ;
    END
  END IN_H
  PIN OE_N
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 123.995000 8.060000 124.775000 8.380000 ;
        RECT 124.325000 7.940000 124.775000 8.060000 ;
        RECT 124.445000 0.000000 124.775000 7.820000 ;
        RECT 124.445000 7.820000 124.775000 7.940000 ;
    END
  END OE_N
  PIN OUT
    ANTENNAGATEAREA  1.529000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.125000  0.000000 74.455000 14.140000 ;
        RECT 74.125000 14.140000 74.455000 14.290000 ;
        RECT 74.125000 14.290000 74.605000 14.440000 ;
        RECT 74.125000 14.440000 74.755000 14.535000 ;
        RECT 74.125000 14.535000 78.505000 14.865000 ;
        RECT 77.870000 51.155000 78.600000 51.485000 ;
        RECT 77.930000 14.865000 78.505000 15.015000 ;
        RECT 77.950000 31.465000 78.355000 31.535000 ;
        RECT 77.950000 31.535000 78.285000 31.605000 ;
        RECT 77.950000 31.605000 78.280000 31.610000 ;
        RECT 77.950000 31.610000 78.280000 33.835000 ;
        RECT 77.950000 33.835000 78.280000 33.905000 ;
        RECT 77.950000 33.905000 78.350000 33.975000 ;
        RECT 77.950000 33.975000 78.420000 33.980000 ;
        RECT 77.990000 31.425000 78.425000 31.465000 ;
        RECT 77.990000 33.980000 78.425000 34.020000 ;
        RECT 78.030000 31.385000 78.465000 31.425000 ;
        RECT 78.030000 34.020000 78.465000 34.060000 ;
        RECT 78.035000 31.380000 78.505000 31.385000 ;
        RECT 78.080000 15.015000 78.505000 15.165000 ;
        RECT 78.100000 34.060000 78.505000 34.130000 ;
        RECT 78.105000 31.310000 78.505000 31.380000 ;
        RECT 78.170000 34.130000 78.505000 34.200000 ;
        RECT 78.175000 15.165000 78.505000 15.260000 ;
        RECT 78.175000 15.260000 78.505000 31.240000 ;
        RECT 78.175000 31.240000 78.505000 31.310000 ;
        RECT 78.175000 34.200000 78.505000 34.205000 ;
        RECT 78.175000 34.205000 78.505000 51.155000 ;
    END
  END OUT
  PIN PAD
    ANTENNAPARTIALMETALSIDEAREA  228.2030 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 40.095000 132.705000 63.135000 147.730000 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    ANTENNAPARTIALMETALSIDEAREA  256.0560 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.240000  5.465000 2.200000   5.470000 ;
        RECT 1.240000  5.470000 2.050000   5.620000 ;
        RECT 1.240000  5.620000 1.900000   5.770000 ;
        RECT 1.240000  5.770000 1.840000   5.830000 ;
        RECT 1.240000  5.830000 1.840000  70.535000 ;
        RECT 1.240000 70.535000 1.840000  70.680000 ;
        RECT 1.240000 70.680000 1.985000  70.825000 ;
        RECT 1.300000  5.405000 2.200000   5.465000 ;
        RECT 1.390000 70.825000 2.130000  70.975000 ;
        RECT 1.450000  5.255000 2.200000   5.405000 ;
        RECT 1.540000 70.975000 2.280000  71.125000 ;
        RECT 1.600000  0.000000 2.200000   5.105000 ;
        RECT 1.600000  5.105000 2.200000   5.255000 ;
        RECT 1.690000 71.125000 2.430000  71.275000 ;
        RECT 1.840000 71.275000 2.580000  71.425000 ;
        RECT 1.990000 71.425000 2.730000  71.575000 ;
        RECT 2.140000 71.575000 2.880000  71.725000 ;
        RECT 2.290000 71.725000 3.030000  71.875000 ;
        RECT 2.440000 71.875000 3.180000  72.025000 ;
        RECT 2.590000 72.025000 3.330000  72.175000 ;
        RECT 2.740000 72.175000 3.480000  72.325000 ;
        RECT 2.890000 72.325000 3.630000  72.475000 ;
        RECT 3.040000 72.475000 3.780000  72.625000 ;
        RECT 3.190000 72.625000 3.930000  72.775000 ;
        RECT 3.340000 72.775000 4.080000  72.925000 ;
        RECT 3.490000 72.925000 4.230000  73.075000 ;
        RECT 3.640000 73.075000 4.380000  73.225000 ;
        RECT 3.725000 73.225000 4.530000  73.310000 ;
        RECT 3.865000 73.310000 4.615000  73.450000 ;
        RECT 4.005000 73.450000 4.615000  73.590000 ;
        RECT 4.010000 73.590000 4.615000  73.595000 ;
        RECT 4.010000 73.595000 4.615000 159.560000 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    ANTENNAPARTIALMETALSIDEAREA  257.9440 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.330000  0.000000 0.930000  71.100000 ;
        RECT 0.330000 71.100000 0.930000  71.240000 ;
        RECT 0.330000 71.240000 1.070000  71.380000 ;
        RECT 0.480000 71.380000 1.210000  71.530000 ;
        RECT 0.630000 71.530000 1.360000  71.680000 ;
        RECT 0.780000 71.680000 1.510000  71.830000 ;
        RECT 0.930000 71.830000 1.660000  71.980000 ;
        RECT 1.080000 71.980000 1.810000  72.130000 ;
        RECT 1.230000 72.130000 1.960000  72.280000 ;
        RECT 1.380000 72.280000 2.110000  72.430000 ;
        RECT 1.530000 72.430000 2.260000  72.580000 ;
        RECT 1.680000 72.580000 2.410000  72.730000 ;
        RECT 1.830000 72.730000 2.560000  72.880000 ;
        RECT 1.980000 72.880000 2.710000  73.030000 ;
        RECT 2.130000 73.030000 2.860000  73.180000 ;
        RECT 2.280000 73.180000 3.010000  73.330000 ;
        RECT 2.430000 73.330000 3.160000  73.480000 ;
        RECT 2.580000 73.480000 3.310000  73.630000 ;
        RECT 2.705000 73.630000 3.460000  73.755000 ;
        RECT 2.845000 73.755000 3.585000  73.895000 ;
        RECT 2.985000 73.895000 3.585000  74.035000 ;
        RECT 2.985000 74.035000 3.585000 160.945000 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    ANTENNAPARTIALCUTAREA  0.120000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2.150000  6.260000 2.975000   6.410000 ;
        RECT 2.150000  6.410000 2.825000   6.560000 ;
        RECT 2.150000  6.560000 2.750000   6.635000 ;
        RECT 2.150000  6.635000 2.750000  70.075000 ;
        RECT 2.150000 70.075000 2.750000  70.220000 ;
        RECT 2.150000 70.220000 2.895000  70.365000 ;
        RECT 2.210000  6.200000 3.125000   6.260000 ;
        RECT 2.300000 70.365000 3.040000  70.515000 ;
        RECT 2.360000  6.050000 3.185000   6.200000 ;
        RECT 2.450000 70.515000 3.190000  70.665000 ;
        RECT 2.510000  5.900000 3.335000   6.050000 ;
        RECT 2.585000  5.825000 3.485000   5.900000 ;
        RECT 2.600000 70.665000 3.340000  70.815000 ;
        RECT 2.735000  5.675000 3.485000   5.825000 ;
        RECT 2.750000 70.815000 3.490000  70.965000 ;
        RECT 2.885000  0.000000 3.485000   5.525000 ;
        RECT 2.885000  5.525000 3.485000   5.675000 ;
        RECT 2.900000 70.965000 3.640000  71.115000 ;
        RECT 3.050000 71.115000 3.790000  71.265000 ;
        RECT 3.200000 71.265000 3.940000  71.415000 ;
        RECT 3.350000 71.415000 4.090000  71.565000 ;
        RECT 3.500000 71.565000 4.240000  71.715000 ;
        RECT 3.650000 71.715000 4.390000  71.865000 ;
        RECT 3.800000 71.865000 4.540000  72.015000 ;
        RECT 3.950000 72.015000 4.690000  72.165000 ;
        RECT 4.100000 72.165000 4.840000  72.315000 ;
        RECT 4.250000 72.315000 4.990000  72.465000 ;
        RECT 4.400000 72.465000 5.140000  72.615000 ;
        RECT 4.550000 72.615000 5.290000  72.765000 ;
        RECT 4.675000 72.765000 5.440000  72.890000 ;
        RECT 4.820000 72.890000 5.565000  73.035000 ;
        RECT 4.965000 73.035000 5.565000  73.180000 ;
        RECT 4.965000 73.180000 5.565000 122.920000 ;
    END
  END PAD_A_NOESD_H
  PIN SLEW_CTL[0]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.085000 0.000000 66.415000 21.685000 ;
    END
  END SLEW_CTL[0]
  PIN SLEW_CTL[1]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.205000 0.000000 46.535000 21.685000 ;
    END
  END SLEW_CTL[1]
  PIN SLOW
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 124.580000 12.150000 125.135000 12.300000 ;
        RECT 124.580000 12.300000 124.985000 12.450000 ;
        RECT 124.580000 12.450000 124.910000 12.525000 ;
        RECT 124.580000 12.525000 124.910000 18.470000 ;
        RECT 124.580000 18.470000 124.910000 18.615000 ;
        RECT 124.580000 18.615000 125.055000 18.760000 ;
        RECT 124.580000 18.760000 125.200000 18.765000 ;
        RECT 124.585000 12.145000 125.285000 12.150000 ;
        RECT 124.675000 12.055000 125.290000 12.145000 ;
        RECT 124.710000 18.765000 125.205000 18.895000 ;
        RECT 124.765000 11.965000 125.380000 12.055000 ;
        RECT 124.840000 11.890000 125.470000 11.965000 ;
        RECT 124.840000 18.895000 125.335000 19.025000 ;
        RECT 124.845000 19.025000 125.465000 19.030000 ;
        RECT 124.990000 11.740000 125.470000 11.890000 ;
        RECT 124.990000 19.030000 125.470000 19.175000 ;
        RECT 125.135000 19.175000 125.470000 19.320000 ;
        RECT 125.140000  0.000000 125.470000 11.590000 ;
        RECT 125.140000 11.590000 125.470000 11.740000 ;
        RECT 125.140000 19.320000 125.470000 19.325000 ;
        RECT 125.140000 19.325000 125.470000 31.390000 ;
    END
  END SLOW
  PIN TIE_HI_ESD
    ANTENNAGATEAREA 21 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.975000   0.000000 130.305000  61.465000 ;
        RECT 129.975000  61.465000 130.305000  61.560000 ;
        RECT 129.975000  61.560000 130.400000  61.655000 ;
        RECT 130.125000  61.655000 130.495000  61.805000 ;
        RECT 130.275000  61.805000 130.645000  61.955000 ;
        RECT 130.425000  61.955000 130.795000  62.105000 ;
        RECT 130.460000 110.205000 131.140000 110.935000 ;
        RECT 130.575000  62.105000 130.945000  62.255000 ;
        RECT 130.620000  62.255000 131.095000  62.300000 ;
        RECT 130.715000  62.300000 131.140000  62.395000 ;
        RECT 130.730000 110.125000 131.140000 110.205000 ;
        RECT 130.810000  62.395000 131.140000  62.490000 ;
        RECT 130.810000  62.490000 131.140000 110.045000 ;
        RECT 130.810000 110.045000 131.140000 110.125000 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    ANTENNAGATEAREA  2.400000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 114.650000 111.180000 115.485000 111.265000 ;
        RECT 114.650000 111.265000 115.400000 111.350000 ;
        RECT 114.670000 111.160000 115.570000 111.180000 ;
        RECT 114.820000 111.010000 115.590000 111.160000 ;
        RECT 114.970000 110.860000 115.740000 111.010000 ;
        RECT 114.990000 110.840000 115.890000 110.860000 ;
        RECT 115.140000 110.690000 115.890000 110.840000 ;
        RECT 115.290000   0.000000 115.890000 110.540000 ;
        RECT 115.290000 110.540000 115.890000 110.690000 ;
    END
  END TIE_LO_ESD
  PIN VINREF
    ANTENNAGATEAREA 54 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.035000 0.000000 44.365000 4.460000 ;
        RECT 44.035000 4.460000 44.365000 4.610000 ;
        RECT 44.035000 4.610000 44.515000 4.760000 ;
        RECT 44.035000 4.760000 44.665000 4.860000 ;
        RECT 44.035000 4.860000 44.765000 5.190000 ;
    END
  END VINREF
  PIN VTRIP_SEL
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 87.665000 0.000000 87.995000 21.685000 ;
    END
  END VTRIP_SEL
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.255000  8.930000 140.000000 13.465000 ;
        RECT 138.730000  8.885000 140.000000  8.930000 ;
        RECT 138.730000 13.465000 140.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 8.985000 140.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 2.035000 140.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 2.135000 140.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 139.035000 14.935000 140.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 139.035000 15.035000 140.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 19.785000 140.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 70.035000 140.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 19.885000 140.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 70.035000 140.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 64.085000 140.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 64.185000 140.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 36.735000 140.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 47.735000 140.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 51.645000 140.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 56.405000 140.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 36.840000 140.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 47.735000 140.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 41.585000 140.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 41.685000 140.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 175.785000 140.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 25.835000 140.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 175.785000 140.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 25.935000 140.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 58.235000 140.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 58.335000 140.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 31.885000 140.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 31.985000 140.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  10.485000 187.010000  10.715000 187.105000 ;
      RECT  10.485000 187.105000  10.830000 187.335000 ;
      RECT  11.220000 170.660000  15.760000 172.700000 ;
      RECT  11.395000 162.715000  13.005000 163.245000 ;
      RECT  11.600000  17.150000  16.580000  18.770000 ;
      RECT  11.600000  18.770000 140.000000  20.300000 ;
      RECT  11.600000  20.300000  22.570000  20.755000 ;
      RECT  13.915000 162.715000  15.525000 163.245000 ;
      RECT  18.005000  10.045000  18.175000  10.575000 ;
      RECT  32.245000  17.150000 140.000000  18.770000 ;
      RECT  69.500000  59.375000  69.820000  59.965000 ;
      RECT  84.135000  47.800000  88.065000  47.970000 ;
      RECT 118.305000 114.495000 140.145000 116.765000 ;
      RECT 120.645000  82.020000 123.195000  96.125000 ;
      RECT 120.725000  81.690000 123.195000  82.020000 ;
      RECT 129.625000  57.445000 131.645000  58.925000 ;
      RECT 131.375000 110.400000 140.145000 114.495000 ;
      RECT 135.060000  74.915000 135.565000 104.150000 ;
      RECT 135.140000  74.890000 135.565000  74.915000 ;
      RECT 135.140000 104.150000 135.565000 104.230000 ;
      RECT 136.065000 186.065000 138.125000 186.295000 ;
      RECT 136.065000 186.295000 136.295000 186.895000 ;
      RECT 136.065000 187.570000 136.295000 187.870000 ;
      RECT 136.065000 187.870000 138.125000 188.100000 ;
      RECT 136.815000 187.175000 137.345000 187.345000 ;
      RECT 137.895000 186.295000 138.125000 187.870000 ;
    LAYER met1 ;
      RECT   0.000000  0.000000 140.000000 200.000000 ;
      RECT 140.000000 53.225000 140.350000  53.955000 ;
      RECT 140.000000 63.715000 140.160000  64.685000 ;
    LAYER met2 ;
      RECT 0.000000  0.000000 140.000000  63.715000 ;
      RECT 0.000000 63.715000 140.325000  68.140000 ;
      RECT 0.000000 68.140000 140.000000 200.000000 ;
    LAYER met3 ;
      RECT   0.000000   0.000000   0.030000  71.505000 ;
      RECT   0.000000  71.505000   2.685000  74.160000 ;
      RECT   0.000000  71.765000   0.150000  71.915000 ;
      RECT   0.000000  71.915000   0.300000  72.065000 ;
      RECT   0.000000  72.065000   0.450000  72.215000 ;
      RECT   0.000000  72.215000   0.600000  72.365000 ;
      RECT   0.000000  72.365000   0.750000  72.515000 ;
      RECT   0.000000  72.515000   0.900000  72.665000 ;
      RECT   0.000000  72.665000   1.050000  72.815000 ;
      RECT   0.000000  72.815000   1.200000  72.965000 ;
      RECT   0.000000  72.965000   1.350000  73.115000 ;
      RECT   0.000000  73.115000   1.500000  73.265000 ;
      RECT   0.000000  73.265000   1.650000  73.415000 ;
      RECT   0.000000  73.415000   1.800000  73.565000 ;
      RECT   0.000000  73.565000   1.950000  73.715000 ;
      RECT   0.000000  73.715000   2.100000  73.865000 ;
      RECT   0.000000  73.865000   2.250000  74.015000 ;
      RECT   0.000000  74.015000   2.400000  74.165000 ;
      RECT   0.000000  74.160000   2.685000 161.245000 ;
      RECT   0.000000  74.165000   2.550000  74.200000 ;
      RECT   0.000000  74.200000   2.585000 161.345000 ;
      RECT   0.000000 161.245000 140.000000 200.000000 ;
      RECT   0.000000 161.345000 140.000000 200.000000 ;
      RECT   1.230000   0.000000   1.300000   4.980000 ;
      RECT   2.500000   0.000000   2.585000   5.400000 ;
      RECT   3.050000   6.760000   5.465000  13.505000 ;
      RECT   3.050000  13.505000   6.810000  20.035000 ;
      RECT   3.050000  20.035000  19.650000  23.165000 ;
      RECT   3.050000  23.165000  21.835000  32.575000 ;
      RECT   3.050000  32.575000  77.650000  34.105000 ;
      RECT   3.050000  34.105000  77.875000  34.330000 ;
      RECT   3.050000  34.330000  77.875000  50.855000 ;
      RECT   3.050000  50.855000  77.570000  51.785000 ;
      RECT   3.050000  51.785000 114.990000  69.950000 ;
      RECT   3.050000  69.950000 114.990000  72.765000 ;
      RECT   3.150000   6.800000   5.365000  13.605000 ;
      RECT   3.150000  13.605000   6.710000  20.135000 ;
      RECT   3.150000  13.605000   6.710000  23.265000 ;
      RECT   3.150000  20.135000  19.550000  23.265000 ;
      RECT   3.150000  20.135000  19.550000  32.675000 ;
      RECT   3.150000  23.265000  21.735000  32.675000 ;
      RECT   3.150000  23.265000  21.735000  34.145000 ;
      RECT   3.150000  23.265000  21.735000  34.145000 ;
      RECT   3.150000  23.265000  21.735000  34.145000 ;
      RECT   3.150000  32.675000  77.550000  34.145000 ;
      RECT   3.150000  32.675000  77.550000  50.755000 ;
      RECT   3.150000  32.675000  77.550000  50.755000 ;
      RECT   3.150000  32.675000  77.550000  50.755000 ;
      RECT   3.150000  32.675000  77.550000  50.755000 ;
      RECT   3.150000  34.145000  77.550000  34.260000 ;
      RECT   3.150000  34.145000  77.550000  34.260000 ;
      RECT   3.150000  34.260000  77.665000  34.370000 ;
      RECT   3.150000  34.260000  77.665000  34.370000 ;
      RECT   3.150000  34.370000  77.470000  51.885000 ;
      RECT   3.150000  34.370000  77.470000  69.910000 ;
      RECT   3.150000  34.370000  77.775000  50.755000 ;
      RECT   3.150000  50.755000  77.470000  51.885000 ;
      RECT   3.150000  51.885000 114.890000  69.910000 ;
      RECT   3.285000   6.665000   5.365000   6.800000 ;
      RECT   3.300000  69.910000 114.890000  70.060000 ;
      RECT   3.300000  69.910000 114.890000  70.060000 ;
      RECT   3.435000   6.515000   5.365000   6.665000 ;
      RECT   3.450000  70.060000 114.890000  70.210000 ;
      RECT   3.450000  70.060000 114.890000  70.210000 ;
      RECT   3.585000   6.365000   5.365000   6.515000 ;
      RECT   3.600000  70.210000 114.890000  70.360000 ;
      RECT   3.600000  70.210000 114.890000  70.360000 ;
      RECT   3.735000   6.215000   5.365000   6.365000 ;
      RECT   3.750000  70.360000 114.890000  70.510000 ;
      RECT   3.750000  70.360000 114.890000  70.510000 ;
      RECT   3.785000   0.000000   5.465000   6.025000 ;
      RECT   3.785000   6.025000   5.465000   6.760000 ;
      RECT   3.885000   0.000000   5.365000   6.065000 ;
      RECT   3.885000   6.065000   5.365000   6.215000 ;
      RECT   3.885000 159.860000 140.000000 161.245000 ;
      RECT   3.900000  70.510000 114.890000  70.660000 ;
      RECT   3.900000  70.510000 114.890000  70.660000 ;
      RECT   3.985000 159.960000 140.000000 161.345000 ;
      RECT   3.985000 159.960000 140.000000 200.000000 ;
      RECT   4.050000  70.660000 114.890000  70.810000 ;
      RECT   4.050000  70.660000 114.890000  70.810000 ;
      RECT   4.200000  70.810000 114.890000  70.960000 ;
      RECT   4.200000  70.810000 114.890000  70.960000 ;
      RECT   4.350000  70.960000 114.890000  71.110000 ;
      RECT   4.350000  70.960000 114.890000  71.110000 ;
      RECT   4.500000  71.110000 114.890000  71.260000 ;
      RECT   4.500000  71.110000 114.890000  71.260000 ;
      RECT   4.650000  71.260000 114.890000  71.410000 ;
      RECT   4.650000  71.260000 114.890000  71.410000 ;
      RECT   4.800000  71.410000 114.890000  71.560000 ;
      RECT   4.800000  71.410000 114.890000  71.560000 ;
      RECT   4.915000 123.220000 140.000000 159.860000 ;
      RECT   4.950000  71.560000 114.890000  71.710000 ;
      RECT   4.950000  71.560000 114.890000  71.710000 ;
      RECT   5.015000 123.320000 140.000000 159.960000 ;
      RECT   5.015000 123.320000 140.000000 200.000000 ;
      RECT   5.100000  71.710000 114.890000  71.860000 ;
      RECT   5.100000  71.710000 114.890000  71.860000 ;
      RECT   5.250000  71.860000 114.890000  72.010000 ;
      RECT   5.250000  71.860000 114.890000  72.010000 ;
      RECT   5.400000  72.010000 114.890000  72.160000 ;
      RECT   5.400000  72.010000 114.890000  72.160000 ;
      RECT   5.550000  72.160000 114.890000  72.310000 ;
      RECT   5.550000  72.160000 114.890000  72.310000 ;
      RECT   5.700000  72.310000 114.890000  72.460000 ;
      RECT   5.700000  72.310000 114.890000  72.460000 ;
      RECT   5.850000  72.460000 114.890000  72.610000 ;
      RECT   5.850000  72.460000 114.890000  72.610000 ;
      RECT   5.865000  72.765000 114.990000 110.415000 ;
      RECT   5.865000 110.415000 114.350000 111.055000 ;
      RECT   5.865000 111.055000 114.350000 111.650000 ;
      RECT   5.865000 111.650000 114.965000 112.210000 ;
      RECT   5.865000 112.210000 140.000000 123.220000 ;
      RECT   5.965000  72.610000 114.890000  72.725000 ;
      RECT   5.965000  72.610000 114.890000  72.725000 ;
      RECT   5.965000  72.725000 114.890000 110.375000 ;
      RECT   5.965000 110.375000 114.250000 123.320000 ;
      RECT   5.965000 110.375000 114.250000 123.320000 ;
      RECT   5.965000 110.375000 114.250000 123.320000 ;
      RECT   5.965000 110.375000 114.740000 110.525000 ;
      RECT   5.965000 110.375000 114.740000 110.525000 ;
      RECT   5.965000 110.525000 114.590000 110.675000 ;
      RECT   5.965000 110.525000 114.590000 110.675000 ;
      RECT   5.965000 110.675000 114.440000 110.825000 ;
      RECT   5.965000 110.675000 114.440000 110.825000 ;
      RECT   5.965000 110.825000 114.290000 110.975000 ;
      RECT   5.965000 110.825000 114.290000 110.975000 ;
      RECT   5.965000 110.975000 114.250000 111.015000 ;
      RECT   5.965000 110.975000 114.250000 111.015000 ;
      RECT   5.965000 111.015000 114.250000 111.750000 ;
      RECT   5.965000 111.750000 114.865000 112.450000 ;
      RECT   5.965000 111.750000 114.865000 123.320000 ;
      RECT   5.965000 111.750000 114.865000 123.320000 ;
      RECT   5.965000 111.750000 114.865000 123.320000 ;
      RECT   5.965000 112.450000 140.000000 123.320000 ;
      RECT   6.665000   0.000000   6.810000  13.505000 ;
      RECT   7.740000   0.000000   7.815000  13.760000 ;
      RECT   7.740000  14.690000  19.335000  18.110000 ;
      RECT   7.740000  18.110000  19.650000  18.425000 ;
      RECT   7.740000  18.425000  19.650000  20.035000 ;
      RECT   7.840000  14.790000  19.235000  18.150000 ;
      RECT   7.840000  14.790000  19.235000  18.465000 ;
      RECT   7.840000  18.150000  19.235000  18.300000 ;
      RECT   7.840000  18.150000  19.235000  18.300000 ;
      RECT   7.840000  18.300000  19.385000  18.450000 ;
      RECT   7.840000  18.300000  19.385000  18.450000 ;
      RECT   7.840000  18.450000  19.535000  18.465000 ;
      RECT   7.840000  18.450000  19.535000  18.465000 ;
      RECT   7.840000  18.465000  19.550000  20.135000 ;
      RECT   7.840000  18.465000  19.550000  32.675000 ;
      RECT   8.745000   8.920000  19.335000  13.680000 ;
      RECT   8.745000  13.680000  19.335000  13.945000 ;
      RECT   8.845000   9.020000  19.235000  13.640000 ;
      RECT   8.975000  13.640000  19.235000  13.770000 ;
      RECT   8.975000  13.640000  19.235000  13.770000 ;
      RECT   9.010000  13.945000  19.335000  14.690000 ;
      RECT   9.105000  13.770000  19.235000  13.900000 ;
      RECT   9.105000  13.770000  19.235000  13.900000 ;
      RECT   9.110000   9.020000  19.235000  18.150000 ;
      RECT   9.110000  13.900000  19.235000  13.905000 ;
      RECT   9.110000  13.900000  19.235000  13.905000 ;
      RECT   9.110000  13.905000  19.235000  14.790000 ;
      RECT   9.400000   0.000000  19.335000   8.920000 ;
      RECT   9.500000   0.000000  19.235000   9.020000 ;
      RECT  20.265000  15.575000  21.835000  17.625000 ;
      RECT  20.265000  17.625000  21.835000  17.940000 ;
      RECT  20.365000  15.675000  21.735000  17.585000 ;
      RECT  20.515000  17.585000  21.735000  17.735000 ;
      RECT  20.580000  17.940000  21.835000  23.165000 ;
      RECT  20.665000  17.735000  21.735000  17.885000 ;
      RECT  20.680000  17.885000  21.735000  17.900000 ;
      RECT  20.680000  17.900000  21.735000  23.265000 ;
      RECT  21.010000   0.000000  21.835000  15.575000 ;
      RECT  21.110000   0.000000  21.735000  15.675000 ;
      RECT  22.765000   0.000000  24.080000   0.200000 ;
      RECT  22.765000   0.200000  23.970000   0.310000 ;
      RECT  22.765000   0.310000  23.190000   1.240000 ;
      RECT  22.765000   1.240000  27.055000  13.475000 ;
      RECT  22.765000  13.475000  26.600000  13.930000 ;
      RECT  22.765000  13.930000  26.600000  14.675000 ;
      RECT  22.765000  14.675000  45.905000  21.985000 ;
      RECT  22.765000  21.985000  77.875000  31.115000 ;
      RECT  22.765000  31.115000  77.650000  31.340000 ;
      RECT  22.765000  31.340000  77.650000  31.550000 ;
      RECT  22.765000  31.550000  77.650000  31.645000 ;
      RECT  22.865000   1.340000  26.955000  13.435000 ;
      RECT  22.865000  13.435000  26.500000  22.085000 ;
      RECT  22.865000  13.435000  26.500000  22.085000 ;
      RECT  22.865000  13.435000  26.805000  13.585000 ;
      RECT  22.865000  13.435000  26.805000  13.585000 ;
      RECT  22.865000  13.585000  26.655000  13.735000 ;
      RECT  22.865000  13.585000  26.655000  13.735000 ;
      RECT  22.865000  13.735000  26.505000  13.885000 ;
      RECT  22.865000  13.735000  26.505000  13.885000 ;
      RECT  22.865000  13.885000  26.500000  13.890000 ;
      RECT  22.865000  13.885000  26.500000  13.890000 ;
      RECT  22.865000  13.890000  26.500000  14.775000 ;
      RECT  22.865000  14.775000  45.805000  22.085000 ;
      RECT  22.865000  22.085000  77.550000  31.545000 ;
      RECT  22.865000  22.085000  77.550000  31.545000 ;
      RECT  22.865000  22.085000  77.550000  31.545000 ;
      RECT  22.865000  22.085000  77.550000  31.545000 ;
      RECT  22.865000  22.085000  77.775000  31.075000 ;
      RECT  22.865000  31.075000  77.665000  31.185000 ;
      RECT  22.865000  31.075000  77.665000  31.185000 ;
      RECT  22.865000  31.185000  77.555000  31.295000 ;
      RECT  22.865000  31.185000  77.555000  31.295000 ;
      RECT  22.865000  31.295000  77.550000  31.300000 ;
      RECT  22.865000  31.295000  77.550000  31.300000 ;
      RECT  22.865000  31.300000  77.550000  31.545000 ;
      RECT  23.175000  31.645000  77.650000  32.575000 ;
      RECT  23.275000  22.085000  77.550000  50.755000 ;
      RECT  23.275000  22.085000  77.550000  50.755000 ;
      RECT  23.275000  22.085000  77.550000  50.755000 ;
      RECT  23.275000  22.085000  77.550000  50.755000 ;
      RECT  23.275000  31.545000  77.550000  32.675000 ;
      RECT  25.010000   0.000000  27.055000   1.240000 ;
      RECT  25.110000   0.000000  26.955000   1.340000 ;
      RECT  27.980000  14.355000  45.905000  14.675000 ;
      RECT  27.985000   0.000000  43.735000   5.490000 ;
      RECT  27.985000   5.490000  45.055000   7.485000 ;
      RECT  27.985000   7.485000  44.605000   7.935000 ;
      RECT  27.985000   7.935000  44.605000   8.680000 ;
      RECT  27.985000   8.680000  45.905000  14.355000 ;
      RECT  28.080000  14.455000  45.805000  14.775000 ;
      RECT  28.080000  14.455000  45.805000  22.085000 ;
      RECT  28.085000   0.000000  43.635000   5.590000 ;
      RECT  28.085000   0.000000  43.635000  14.455000 ;
      RECT  28.085000   0.000000  43.635000  14.455000 ;
      RECT  28.085000   5.590000  44.505000  14.455000 ;
      RECT  28.085000   5.590000  44.505000  14.455000 ;
      RECT  28.085000   5.590000  44.955000   7.445000 ;
      RECT  28.085000   7.445000  44.805000   7.595000 ;
      RECT  28.085000   7.445000  44.805000   7.595000 ;
      RECT  28.085000   7.595000  44.655000   7.745000 ;
      RECT  28.085000   7.595000  44.655000   7.745000 ;
      RECT  28.085000   7.745000  44.505000   7.895000 ;
      RECT  28.085000   7.745000  44.505000   7.895000 ;
      RECT  28.085000   7.895000  44.505000   8.780000 ;
      RECT  28.085000   8.780000  45.805000  14.455000 ;
      RECT  28.085000   8.780000  45.805000  14.775000 ;
      RECT  28.085000   8.780000  45.805000  22.085000 ;
      RECT  44.665000   0.000000  45.055000   4.335000 ;
      RECT  44.665000   4.335000  45.055000   4.725000 ;
      RECT  46.835000   0.000000  51.355000   8.680000 ;
      RECT  46.835000   8.680000  65.785000  21.985000 ;
      RECT  46.935000   0.000000  51.255000   8.780000 ;
      RECT  46.935000   0.000000  51.255000  22.085000 ;
      RECT  46.935000   0.000000  51.255000  22.085000 ;
      RECT  46.935000   0.000000  51.255000  22.085000 ;
      RECT  46.935000   8.780000  65.685000  22.085000 ;
      RECT  52.285000   0.000000  64.935000   0.790000 ;
      RECT  52.285000   0.790000  64.860000   0.865000 ;
      RECT  52.285000   0.865000  64.485000   1.785000 ;
      RECT  52.285000   1.785000  65.785000   7.635000 ;
      RECT  52.285000   7.635000  65.785000   7.760000 ;
      RECT  52.385000   0.000000  64.835000   0.765000 ;
      RECT  52.385000   0.765000  64.385000   3.005000 ;
      RECT  52.385000   1.885000  65.685000   7.660000 ;
      RECT  52.735000   7.760000  65.785000   8.680000 ;
      RECT  52.835000   1.885000  65.685000  22.085000 ;
      RECT  52.835000   7.660000  65.685000   8.780000 ;
      RECT  67.565000   0.000000  73.825000  15.165000 ;
      RECT  67.565000  15.165000  77.875000  15.385000 ;
      RECT  67.565000  15.385000  77.875000  21.985000 ;
      RECT  67.665000   0.000000  73.725000  15.265000 ;
      RECT  67.665000  15.265000  77.615000  15.345000 ;
      RECT  67.665000  15.265000  77.615000  15.345000 ;
      RECT  67.665000  15.345000  77.695000  15.425000 ;
      RECT  67.665000  15.345000  77.695000  15.425000 ;
      RECT  67.665000  15.425000  77.775000  22.085000 ;
      RECT  74.755000   0.000000  86.515000  14.015000 ;
      RECT  74.755000  14.015000  86.515000  14.235000 ;
      RECT  74.855000   0.000000  86.510000  13.975000 ;
      RECT  74.935000  13.975000  86.510000  14.055000 ;
      RECT  74.935000  13.975000  86.510000  14.055000 ;
      RECT  75.015000  14.055000  86.510000  14.135000 ;
      RECT  75.015000  14.055000  86.510000  14.135000 ;
      RECT  78.580000  31.735000 114.990000  33.710000 ;
      RECT  78.580000  33.710000 114.990000  33.935000 ;
      RECT  78.680000  31.775000 114.890000  33.670000 ;
      RECT  78.790000  31.665000 114.890000  31.775000 ;
      RECT  78.790000  31.665000 114.890000  31.775000 ;
      RECT  78.790000  33.670000 114.890000  33.780000 ;
      RECT  78.790000  33.670000 114.890000  33.780000 ;
      RECT  78.805000  14.235000  86.515000  21.985000 ;
      RECT  78.805000  21.985000 114.990000  31.510000 ;
      RECT  78.805000  31.510000 114.990000  31.735000 ;
      RECT  78.805000  33.935000 114.990000  50.855000 ;
      RECT  78.900000  33.780000 114.890000  33.890000 ;
      RECT  78.900000  33.780000 114.890000  33.890000 ;
      RECT  78.900000  50.855000 114.990000  51.785000 ;
      RECT  78.905000  14.135000  86.510000  22.085000 ;
      RECT  78.905000  14.135000  86.510000  31.550000 ;
      RECT  78.905000  22.085000 114.890000  31.550000 ;
      RECT  78.905000  22.085000 114.890000  33.895000 ;
      RECT  78.905000  22.085000 114.890000  33.895000 ;
      RECT  78.905000  22.085000 114.890000  33.895000 ;
      RECT  78.905000  22.085000 114.890000  33.895000 ;
      RECT  78.905000  31.550000 114.890000  31.665000 ;
      RECT  78.905000  31.550000 114.890000  31.665000 ;
      RECT  78.905000  33.670000 114.890000  50.755000 ;
      RECT  78.905000  33.670000 114.890000  50.755000 ;
      RECT  78.905000  33.670000 114.890000  50.755000 ;
      RECT  78.905000  33.670000 114.890000  50.755000 ;
      RECT  78.905000  33.890000 114.890000  33.895000 ;
      RECT  78.905000  33.890000 114.890000  33.895000 ;
      RECT  78.905000  33.895000 114.890000  50.755000 ;
      RECT  79.000000  33.895000 114.890000  69.910000 ;
      RECT  79.000000  33.895000 114.890000  69.910000 ;
      RECT  79.000000  50.755000 114.890000  51.885000 ;
      RECT  88.295000   0.000000  95.545000   2.040000 ;
      RECT  88.295000   2.040000 107.245000   7.670000 ;
      RECT  88.295000   7.670000 107.155000   7.760000 ;
      RECT  88.295000   7.760000 106.795000   8.680000 ;
      RECT  88.295000   8.680000 108.095000  19.980000 ;
      RECT  88.295000  19.980000 108.075000  21.985000 ;
      RECT  88.395000   0.000000  95.445000   2.140000 ;
      RECT  88.395000   0.000000  95.445000   7.660000 ;
      RECT  88.395000   0.000000  95.445000   7.660000 ;
      RECT  88.395000   2.140000 106.695000  19.880000 ;
      RECT  88.395000   2.140000 107.145000   7.660000 ;
      RECT  88.395000   7.660000 106.695000   8.780000 ;
      RECT  88.395000   8.780000 107.975000  22.085000 ;
      RECT  88.395000   8.780000 107.975000  22.085000 ;
      RECT  88.395000   8.780000 107.995000  19.880000 ;
      RECT  88.395000  19.880000 107.975000  22.085000 ;
      RECT  96.515000   0.000000 107.245000   2.040000 ;
      RECT  96.615000   0.000000 107.145000   2.140000 ;
      RECT  96.615000   0.000000 107.145000   7.660000 ;
      RECT  96.615000   0.000000 107.145000   7.660000 ;
      RECT 109.005000  20.940000 114.990000  21.985000 ;
      RECT 109.025000   0.000000 114.990000  20.940000 ;
      RECT 109.105000  21.040000 114.890000  22.085000 ;
      RECT 109.125000   0.000000 114.890000  21.040000 ;
      RECT 109.125000   0.000000 114.890000  22.085000 ;
      RECT 109.125000   0.000000 114.890000  22.085000 ;
      RECT 114.930000 112.385000 140.000000 112.450000 ;
      RECT 114.930000 112.385000 140.000000 112.450000 ;
      RECT 115.080000 112.235000 140.000000 112.385000 ;
      RECT 115.080000 112.235000 140.000000 112.385000 ;
      RECT 115.230000 112.085000 140.000000 112.235000 ;
      RECT 115.230000 112.085000 140.000000 112.235000 ;
      RECT 115.380000 111.935000 140.000000 112.085000 ;
      RECT 115.380000 111.935000 140.000000 112.085000 ;
      RECT 115.530000 111.785000 140.000000 111.935000 ;
      RECT 115.530000 111.785000 140.000000 111.935000 ;
      RECT 115.680000 111.635000 140.000000 111.785000 ;
      RECT 115.680000 111.635000 140.000000 111.785000 ;
      RECT 115.830000 111.485000 140.000000 111.635000 ;
      RECT 115.830000 111.485000 140.000000 111.635000 ;
      RECT 115.940000 111.235000 140.000000 112.210000 ;
      RECT 115.980000 111.335000 140.000000 111.485000 ;
      RECT 115.980000 111.335000 140.000000 111.485000 ;
      RECT 115.990000 111.325000 130.060000 111.335000 ;
      RECT 115.990000 111.325000 130.060000 111.335000 ;
      RECT 116.140000 111.175000 130.060000 111.325000 ;
      RECT 116.140000 111.175000 130.060000 111.325000 ;
      RECT 116.190000   0.000000 124.145000   7.695000 ;
      RECT 116.190000   7.695000 124.080000   7.760000 ;
      RECT 116.190000   7.760000 123.695000   8.680000 ;
      RECT 116.190000   8.680000 124.840000  11.465000 ;
      RECT 116.190000  11.465000 124.280000  12.025000 ;
      RECT 116.190000  12.025000 124.280000  18.890000 ;
      RECT 116.190000  18.890000 124.840000  19.450000 ;
      RECT 116.190000  19.450000 124.840000  31.690000 ;
      RECT 116.190000  31.690000 129.675000  61.780000 ;
      RECT 116.190000  61.780000 130.510000  62.615000 ;
      RECT 116.190000  62.615000 130.510000 109.905000 ;
      RECT 116.190000 109.905000 130.160000 110.985000 ;
      RECT 116.190000 110.985000 130.160000 111.235000 ;
      RECT 116.290000   0.000000 123.595000  11.985000 ;
      RECT 116.290000   0.000000 123.595000  18.930000 ;
      RECT 116.290000   0.000000 124.045000   7.660000 ;
      RECT 116.290000   7.660000 123.595000   8.780000 ;
      RECT 116.290000   8.780000 124.180000  18.930000 ;
      RECT 116.290000   8.780000 124.740000  11.425000 ;
      RECT 116.290000  11.425000 124.590000  11.575000 ;
      RECT 116.290000  11.425000 124.590000  11.575000 ;
      RECT 116.290000  11.575000 124.440000  11.725000 ;
      RECT 116.290000  11.575000 124.440000  11.725000 ;
      RECT 116.290000  11.725000 124.290000  11.875000 ;
      RECT 116.290000  11.725000 124.290000  11.875000 ;
      RECT 116.290000  11.875000 124.180000  11.985000 ;
      RECT 116.290000  11.875000 124.180000  11.985000 ;
      RECT 116.290000  11.985000 124.180000  18.930000 ;
      RECT 116.290000  11.985000 124.180000  19.490000 ;
      RECT 116.290000  18.930000 124.180000  19.080000 ;
      RECT 116.290000  18.930000 124.180000  19.080000 ;
      RECT 116.290000  19.080000 124.330000  19.230000 ;
      RECT 116.290000  19.080000 124.330000  19.230000 ;
      RECT 116.290000  19.230000 124.480000  19.380000 ;
      RECT 116.290000  19.230000 124.480000  19.380000 ;
      RECT 116.290000  19.380000 124.630000  19.490000 ;
      RECT 116.290000  19.380000 124.630000  19.490000 ;
      RECT 116.290000  19.490000 124.740000  31.790000 ;
      RECT 116.290000  19.490000 124.740000  61.820000 ;
      RECT 116.290000  31.790000 129.575000  61.820000 ;
      RECT 116.290000  61.820000 129.575000  61.970000 ;
      RECT 116.290000  61.820000 129.575000  61.970000 ;
      RECT 116.290000  61.970000 129.725000  62.120000 ;
      RECT 116.290000  61.970000 129.725000  62.120000 ;
      RECT 116.290000  62.120000 129.875000  62.270000 ;
      RECT 116.290000  62.120000 129.875000  62.270000 ;
      RECT 116.290000  62.270000 130.025000  62.420000 ;
      RECT 116.290000  62.270000 130.025000  62.420000 ;
      RECT 116.290000  62.420000 130.175000  62.570000 ;
      RECT 116.290000  62.420000 130.175000  62.570000 ;
      RECT 116.290000  62.570000 130.325000  62.655000 ;
      RECT 116.290000  62.570000 130.325000  62.655000 ;
      RECT 116.290000  62.655000 130.410000 109.805000 ;
      RECT 116.290000 109.805000 130.060000 111.025000 ;
      RECT 116.290000 111.025000 130.060000 111.175000 ;
      RECT 116.290000 111.025000 130.060000 111.175000 ;
      RECT 125.210000  12.650000 127.975000  18.345000 ;
      RECT 125.210000  18.345000 127.975000  18.905000 ;
      RECT 125.310000  12.690000 127.875000  18.305000 ;
      RECT 125.420000  12.580000 127.875000  12.690000 ;
      RECT 125.460000  18.305000 127.875000  18.455000 ;
      RECT 125.570000  12.430000 127.875000  12.580000 ;
      RECT 125.610000  18.455000 127.875000  18.605000 ;
      RECT 125.720000  12.280000 127.875000  12.430000 ;
      RECT 125.760000  18.605000 127.875000  18.755000 ;
      RECT 125.770000   0.000000 127.975000  12.090000 ;
      RECT 125.770000  12.090000 127.975000  12.650000 ;
      RECT 125.770000  18.905000 127.975000  20.305000 ;
      RECT 125.770000  20.305000 127.995000  20.325000 ;
      RECT 125.770000  20.325000 127.995000  21.985000 ;
      RECT 125.770000  21.985000 129.675000  31.690000 ;
      RECT 125.870000   0.000000 127.875000  12.130000 ;
      RECT 125.870000  12.130000 127.875000  12.280000 ;
      RECT 125.870000  18.755000 127.875000  18.865000 ;
      RECT 125.870000  18.865000 127.875000  20.345000 ;
      RECT 125.870000  20.345000 127.875000  20.355000 ;
      RECT 125.870000  20.355000 127.885000  20.365000 ;
      RECT 125.870000  20.365000 127.895000  22.085000 ;
      RECT 125.870000  22.085000 129.575000  31.790000 ;
      RECT 130.605000   0.000000 140.000000  61.340000 ;
      RECT 130.605000  61.340000 140.000000  62.175000 ;
      RECT 130.705000   0.000000 140.000000  61.300000 ;
      RECT 130.855000  61.300000 140.000000  61.450000 ;
      RECT 130.855000  61.300000 140.000000  61.450000 ;
      RECT 131.005000  61.450000 140.000000  61.600000 ;
      RECT 131.005000  61.450000 140.000000  61.600000 ;
      RECT 131.155000  61.600000 140.000000  61.750000 ;
      RECT 131.155000  61.600000 140.000000  61.750000 ;
      RECT 131.305000  61.750000 140.000000  61.900000 ;
      RECT 131.305000  61.750000 140.000000  61.900000 ;
      RECT 131.440000  62.175000 140.000000 111.235000 ;
      RECT 131.455000  61.900000 140.000000  62.050000 ;
      RECT 131.455000  61.900000 140.000000  62.050000 ;
      RECT 131.540000  62.050000 140.000000  62.135000 ;
      RECT 131.540000  62.050000 140.000000  62.135000 ;
      RECT 131.540000  62.135000 140.000000 111.335000 ;
      RECT 131.540000  62.135000 140.000000 112.450000 ;
    LAYER met4 ;
      RECT   0.000000   0.000000   1.670000   1.635000 ;
      RECT   0.000000   0.000000 140.000000   1.635000 ;
      RECT   0.000000   7.885000   1.670000   8.485000 ;
      RECT   0.000000   7.885000 140.000000   8.485000 ;
      RECT   0.000000  13.935000   1.365000  14.535000 ;
      RECT   0.000000  13.935000 140.000000  14.535000 ;
      RECT   0.000000  18.785000   1.365000  19.385000 ;
      RECT   0.000000  18.785000 140.000000  19.385000 ;
      RECT   0.000000  24.835000   1.670000  25.435000 ;
      RECT   0.000000  24.835000 140.000000  25.435000 ;
      RECT   0.000000  30.885000   1.670000  31.485000 ;
      RECT   0.000000  30.885000 140.000000  31.485000 ;
      RECT   0.000000  35.735000   1.670000  36.335000 ;
      RECT   0.000000  35.735000 140.000000  36.335000 ;
      RECT   0.000000  40.585000   1.670000  41.185000 ;
      RECT   0.000000  40.585000 140.000000  41.185000 ;
      RECT   0.000000  46.635000   1.670000  47.335000 ;
      RECT   0.000000  46.635000 140.000000  47.435000 ;
      RECT   0.000000  57.035000 140.000000  57.835000 ;
      RECT   0.000000  57.135000   1.670000  57.835000 ;
      RECT   0.000000  63.085000   1.670000  63.685000 ;
      RECT   0.000000  63.085000 140.000000  63.685000 ;
      RECT   0.000000  68.935000   1.670000  69.635000 ;
      RECT   0.000000  68.935000 140.000000  69.635000 ;
      RECT   0.000000  95.400000 140.000000 175.385000 ;
      RECT   1.365000  13.935000 138.635000  19.385000 ;
      RECT   1.365000  13.935000 138.635000  19.385000 ;
      RECT   1.570000  47.435000 138.430000  57.035000 ;
      RECT   1.670000   0.000000 137.855000 200.000000 ;
      RECT   1.670000   0.000000 138.330000   8.530000 ;
      RECT   1.670000   0.000000 138.330000   8.530000 ;
      RECT   1.670000   0.000000 138.330000   8.530000 ;
      RECT   1.670000   8.485000 140.000000   8.585000 ;
      RECT   1.670000   8.530000 137.855000  13.865000 ;
      RECT   1.670000   8.585000 138.430000   8.630000 ;
      RECT   1.670000   8.630000 137.955000  13.765000 ;
      RECT   1.670000  13.765000 138.430000  13.835000 ;
      RECT   1.670000  13.835000 140.000000  13.935000 ;
      RECT   1.670000  13.865000 138.330000  13.935000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  19.385000 138.330000  95.400000 ;
      RECT   1.670000 175.385000 138.330000 200.000000 ;
      RECT 138.330000   0.000000 140.000000   1.635000 ;
      RECT 138.330000   7.885000 140.000000   8.485000 ;
      RECT 138.330000  24.835000 140.000000  25.435000 ;
      RECT 138.330000  30.885000 140.000000  31.485000 ;
      RECT 138.330000  35.735000 140.000000  36.335000 ;
      RECT 138.330000  40.585000 140.000000  41.185000 ;
      RECT 138.330000  46.635000 140.000000  47.335000 ;
      RECT 138.330000  57.135000 140.000000  57.835000 ;
      RECT 138.330000  63.085000 140.000000  63.685000 ;
      RECT 138.330000  68.935000 140.000000  69.635000 ;
      RECT 138.635000  13.935000 140.000000  14.535000 ;
      RECT 138.635000  18.785000 140.000000  19.385000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000 140.000000   1.335000 ;
      RECT  0.000000  36.035000 140.000000  36.040000 ;
      RECT  0.000000  95.785000 140.000000 131.905000 ;
      RECT  0.000000 131.905000  39.295000 148.530000 ;
      RECT  0.000000 148.530000 140.000000 174.985000 ;
      RECT  1.765000  14.235000 138.235000  19.085000 ;
      RECT  2.070000   1.335000 137.930000  14.235000 ;
      RECT  2.070000  19.085000 137.930000  95.785000 ;
      RECT  2.070000 174.985000 137.930000 200.000000 ;
      RECT  9.605000  96.585000 126.350000 103.180000 ;
      RECT 11.565000 171.780000  99.610000 174.185000 ;
      RECT 63.935000 131.905000 140.000000 148.530000 ;
  END
END sky130_fd_io__top_gpio_ovtv2


MACRO sky130_fd_io__top_ground_hvc_wpad
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN G_PAD
    ANTENNAPARTIALMETALSIDEAREA  284.1730 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 36.645000 139.325000 37.970000 145.935000 ;
    END
  END G_PAD
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 15.620000 185.295000 74.290000 190.015000 ;
        RECT 16.805000  47.455000 74.290000  54.765000 ;
        RECT 16.805000 139.455000 74.290000 146.710000 ;
        RECT 16.805000 162.455000 74.290000 171.155000 ;
        RECT 16.875000 146.710000 74.290000 146.780000 ;
        RECT 16.945000 146.780000 74.290000 146.850000 ;
        RECT 17.015000 146.850000 74.290000 146.920000 ;
        RECT 17.085000 146.920000 74.290000 146.990000 ;
        RECT 17.155000 146.990000 74.290000 147.060000 ;
        RECT 17.225000 147.060000 74.290000 147.130000 ;
        RECT 17.295000 147.130000 74.290000 147.200000 ;
        RECT 17.365000 147.200000 74.290000 147.270000 ;
        RECT 17.435000 147.270000 74.290000 147.340000 ;
        RECT 17.505000 147.340000 74.290000 147.410000 ;
        RECT 17.530000  54.765000 74.290000  54.835000 ;
        RECT 17.575000 147.410000 74.290000 147.480000 ;
        RECT 17.600000  54.835000 74.290000  54.905000 ;
        RECT 17.645000 147.480000 74.290000 147.550000 ;
        RECT 17.670000  54.905000 74.290000  54.975000 ;
        RECT 17.715000 147.550000 74.290000 147.620000 ;
        RECT 17.740000  54.975000 74.290000  55.045000 ;
        RECT 17.785000 147.620000 74.290000 147.690000 ;
        RECT 17.810000  55.045000 74.290000  55.115000 ;
        RECT 17.855000 147.690000 74.290000 147.760000 ;
        RECT 17.880000  55.115000 74.290000  55.185000 ;
        RECT 17.925000 147.760000 74.290000 147.830000 ;
        RECT 17.950000  55.185000 74.290000  55.255000 ;
        RECT 17.995000 147.830000 74.290000 147.900000 ;
        RECT 18.020000  55.255000 74.290000  55.325000 ;
        RECT 18.065000 147.900000 74.290000 147.970000 ;
        RECT 18.090000  55.325000 74.290000  55.395000 ;
        RECT 18.135000 147.970000 74.290000 148.040000 ;
        RECT 18.160000  55.395000 74.290000  55.465000 ;
        RECT 18.205000 148.040000 74.290000 148.110000 ;
        RECT 18.230000  55.465000 74.290000  55.535000 ;
        RECT 18.250000 148.110000 74.290000 148.155000 ;
        RECT 18.300000  55.535000 74.290000  55.605000 ;
        RECT 18.370000  55.605000 74.290000  55.675000 ;
        RECT 18.410000  74.155000 74.290000  74.415000 ;
        RECT 18.440000  55.675000 74.290000  55.745000 ;
        RECT 18.510000  55.745000 74.290000  55.815000 ;
        RECT 18.580000  55.815000 74.290000  55.885000 ;
        RECT 18.650000  55.885000 74.290000  55.955000 ;
        RECT 18.720000  55.955000 74.290000  56.025000 ;
        RECT 18.790000  56.025000 74.290000  56.095000 ;
        RECT 18.850000  56.095000 74.290000  56.155000 ;
        RECT 23.690000  74.415000 74.290000  74.485000 ;
        RECT 23.700000  74.105000 74.290000  74.155000 ;
        RECT 23.760000  74.485000 74.290000  74.555000 ;
        RECT 23.770000  74.035000 74.290000  74.105000 ;
        RECT 23.830000  74.555000 74.290000  74.625000 ;
        RECT 23.840000  73.965000 74.290000  74.035000 ;
        RECT 23.900000  74.625000 74.290000  74.695000 ;
        RECT 23.910000  73.895000 74.290000  73.965000 ;
        RECT 23.970000  74.695000 74.290000  74.765000 ;
        RECT 23.980000  73.825000 74.290000  73.895000 ;
        RECT 24.040000  74.765000 74.290000  74.835000 ;
        RECT 24.050000  73.755000 74.290000  73.825000 ;
        RECT 24.110000  74.835000 74.290000  74.905000 ;
        RECT 24.120000  73.685000 74.290000  73.755000 ;
        RECT 24.180000  74.905000 74.290000  74.975000 ;
        RECT 24.190000  73.615000 74.290000  73.685000 ;
        RECT 24.250000  74.975000 74.290000  75.045000 ;
        RECT 24.260000  73.545000 74.290000  73.615000 ;
        RECT 24.320000  75.045000 74.290000  75.115000 ;
        RECT 24.330000  73.475000 74.290000  73.545000 ;
        RECT 24.390000  75.115000 74.290000  75.185000 ;
        RECT 24.400000  73.405000 74.290000  73.475000 ;
        RECT 24.460000  75.185000 74.290000  75.255000 ;
        RECT 24.470000  73.335000 74.290000  73.405000 ;
        RECT 24.530000  75.255000 74.290000  75.325000 ;
        RECT 24.540000  73.265000 74.290000  73.335000 ;
        RECT 24.600000  75.325000 74.290000  75.395000 ;
        RECT 24.610000  73.195000 74.290000  73.265000 ;
        RECT 24.670000  75.395000 74.290000  75.465000 ;
        RECT 24.680000  73.125000 74.290000  73.195000 ;
        RECT 24.740000  75.465000 74.290000  75.535000 ;
        RECT 24.750000  73.055000 74.290000  73.125000 ;
        RECT 24.810000  75.535000 74.290000  75.605000 ;
        RECT 24.820000  70.455000 74.290000  72.985000 ;
        RECT 24.820000  72.985000 74.290000  73.055000 ;
        RECT 24.820000  75.605000 74.290000  75.615000 ;
        RECT 24.820000  75.615000 74.290000  79.155000 ;
        RECT 24.820000  93.455000 74.290000 102.155000 ;
        RECT 24.820000 116.455000 74.290000 125.155000 ;
        RECT 37.890000  12.295000 74.290000  25.660000 ;
        RECT 46.750000  12.265000 74.290000  12.295000 ;
        RECT 46.820000  12.195000 74.290000  12.265000 ;
        RECT 46.890000  12.125000 74.290000  12.195000 ;
        RECT 46.960000  12.055000 74.290000  12.125000 ;
        RECT 47.030000  11.985000 74.290000  12.055000 ;
        RECT 47.100000  11.915000 74.290000  11.985000 ;
        RECT 47.170000  11.845000 74.290000  11.915000 ;
        RECT 47.240000  11.775000 74.290000  11.845000 ;
        RECT 47.310000  11.705000 74.290000  11.775000 ;
        RECT 47.380000  11.635000 74.290000  11.705000 ;
        RECT 47.450000  11.565000 74.290000  11.635000 ;
        RECT 47.520000  11.495000 74.290000  11.565000 ;
        RECT 47.590000  11.425000 74.290000  11.495000 ;
        RECT 47.660000  11.355000 74.290000  11.425000 ;
        RECT 47.730000  11.285000 74.290000  11.355000 ;
        RECT 47.800000  11.215000 74.290000  11.285000 ;
        RECT 47.870000  11.145000 74.290000  11.215000 ;
        RECT 47.940000  11.075000 74.290000  11.145000 ;
        RECT 48.010000  11.005000 74.290000  11.075000 ;
        RECT 48.080000  10.935000 74.290000  11.005000 ;
        RECT 48.150000  10.865000 74.290000  10.935000 ;
        RECT 48.220000  10.795000 74.290000  10.865000 ;
        RECT 48.290000  10.725000 74.290000  10.795000 ;
        RECT 48.360000  10.655000 74.290000  10.725000 ;
        RECT 48.430000  10.585000 74.290000  10.655000 ;
        RECT 48.500000  10.515000 74.290000  10.585000 ;
        RECT 48.570000  10.445000 74.290000  10.515000 ;
        RECT 48.640000  10.375000 74.290000  10.445000 ;
        RECT 48.710000  10.305000 74.290000  10.375000 ;
        RECT 48.780000  10.235000 74.290000  10.305000 ;
        RECT 48.850000  10.165000 74.290000  10.235000 ;
        RECT 48.920000  10.095000 74.290000  10.165000 ;
        RECT 48.990000  10.025000 74.290000  10.095000 ;
        RECT 49.060000   9.955000 74.290000  10.025000 ;
        RECT 49.130000   9.885000 74.290000   9.955000 ;
        RECT 49.200000   9.815000 74.290000   9.885000 ;
        RECT 49.270000   9.745000 74.290000   9.815000 ;
        RECT 49.340000   9.675000 74.290000   9.745000 ;
        RECT 49.410000   9.605000 74.290000   9.675000 ;
        RECT 49.480000   9.535000 74.290000   9.605000 ;
        RECT 49.550000   9.465000 74.290000   9.535000 ;
        RECT 49.620000   9.395000 74.290000   9.465000 ;
        RECT 49.690000   9.325000 74.290000   9.395000 ;
        RECT 49.760000   9.255000 74.290000   9.325000 ;
        RECT 49.830000   9.185000 74.290000   9.255000 ;
        RECT 49.900000   9.115000 74.290000   9.185000 ;
        RECT 49.970000   9.045000 74.290000   9.115000 ;
        RECT 50.040000   8.975000 74.290000   9.045000 ;
        RECT 50.110000   8.905000 74.290000   8.975000 ;
        RECT 50.180000   8.835000 74.290000   8.905000 ;
        RECT 50.250000   8.765000 74.290000   8.835000 ;
        RECT 50.320000   8.695000 74.290000   8.765000 ;
        RECT 50.390000   0.000000 74.290000   8.625000 ;
        RECT 50.390000   8.625000 74.290000   8.695000 ;
        RECT 55.885000  25.660000 74.290000  25.730000 ;
        RECT 55.955000  25.730000 74.290000  25.800000 ;
        RECT 56.025000  25.800000 74.290000  25.870000 ;
        RECT 56.095000  25.870000 74.290000  25.940000 ;
        RECT 56.165000  25.940000 74.290000  26.010000 ;
        RECT 56.235000  26.010000 74.290000  26.080000 ;
        RECT 56.305000  26.080000 74.290000  26.150000 ;
        RECT 56.375000  26.150000 74.290000  26.220000 ;
        RECT 56.445000  26.220000 74.290000  26.290000 ;
        RECT 56.515000  26.290000 74.290000  26.360000 ;
        RECT 56.585000  26.360000 74.290000  26.430000 ;
        RECT 56.655000  26.430000 74.290000  26.500000 ;
        RECT 56.725000  26.500000 74.290000  26.570000 ;
        RECT 56.795000  26.570000 74.290000  26.640000 ;
        RECT 56.865000  26.640000 74.290000  26.710000 ;
        RECT 56.935000  26.710000 74.290000  26.780000 ;
        RECT 57.005000  26.780000 74.290000  26.850000 ;
        RECT 57.075000  26.850000 74.290000  26.920000 ;
        RECT 57.145000  26.920000 74.290000  26.990000 ;
        RECT 57.215000  26.990000 74.290000  27.060000 ;
        RECT 57.285000  27.060000 74.290000  27.130000 ;
        RECT 57.355000  27.130000 74.290000  27.200000 ;
        RECT 57.425000  27.200000 74.290000  27.270000 ;
        RECT 57.495000  27.270000 74.290000  27.340000 ;
        RECT 57.540000  47.390000 74.290000  47.455000 ;
        RECT 57.540000  70.420000 74.290000  70.455000 ;
        RECT 57.540000 116.390000 74.290000 116.455000 ;
        RECT 57.540000 139.425000 74.290000 139.455000 ;
        RECT 57.540000 162.440000 74.290000 162.455000 ;
        RECT 57.555000 148.155000 74.290000 148.225000 ;
        RECT 57.565000  27.340000 74.290000  27.410000 ;
        RECT 57.595000  56.155000 74.290000  56.225000 ;
        RECT 57.610000  47.320000 74.290000  47.390000 ;
        RECT 57.610000  70.350000 74.290000  70.420000 ;
        RECT 57.610000  93.410000 74.290000  93.455000 ;
        RECT 57.610000 116.320000 74.290000 116.390000 ;
        RECT 57.610000 139.355000 74.290000 139.425000 ;
        RECT 57.610000 162.370000 74.290000 162.440000 ;
        RECT 57.625000  79.155000 74.290000  79.225000 ;
        RECT 57.625000 102.155000 74.290000 102.225000 ;
        RECT 57.625000 125.155000 74.290000 125.225000 ;
        RECT 57.625000 148.225000 74.290000 148.295000 ;
        RECT 57.635000  27.410000 74.290000  27.480000 ;
        RECT 57.635000 171.155000 74.290000 171.225000 ;
        RECT 57.665000  56.225000 74.290000  56.295000 ;
        RECT 57.680000  47.250000 74.290000  47.320000 ;
        RECT 57.680000  70.280000 74.290000  70.350000 ;
        RECT 57.680000  93.340000 74.290000  93.410000 ;
        RECT 57.680000 116.250000 74.290000 116.320000 ;
        RECT 57.680000 139.285000 74.290000 139.355000 ;
        RECT 57.680000 162.300000 74.290000 162.370000 ;
        RECT 57.695000  79.225000 74.290000  79.295000 ;
        RECT 57.695000 102.225000 74.290000 102.295000 ;
        RECT 57.695000 125.225000 74.290000 125.295000 ;
        RECT 57.695000 148.295000 74.290000 148.365000 ;
        RECT 57.705000  27.480000 74.290000  27.550000 ;
        RECT 57.705000 171.225000 74.290000 171.295000 ;
        RECT 57.735000  56.295000 74.290000  56.365000 ;
        RECT 57.750000  47.180000 74.290000  47.250000 ;
        RECT 57.750000  70.210000 74.290000  70.280000 ;
        RECT 57.750000  93.270000 74.290000  93.340000 ;
        RECT 57.750000 116.180000 74.290000 116.250000 ;
        RECT 57.750000 139.215000 74.290000 139.285000 ;
        RECT 57.750000 162.230000 74.290000 162.300000 ;
        RECT 57.765000  79.295000 74.290000  79.365000 ;
        RECT 57.765000 102.295000 74.290000 102.365000 ;
        RECT 57.765000 125.295000 74.290000 125.365000 ;
        RECT 57.765000 148.365000 74.290000 148.435000 ;
        RECT 57.775000  27.550000 74.290000  27.620000 ;
        RECT 57.775000 171.295000 74.290000 171.365000 ;
        RECT 57.805000  56.365000 74.290000  56.435000 ;
        RECT 57.820000  47.110000 74.290000  47.180000 ;
        RECT 57.820000  70.140000 74.290000  70.210000 ;
        RECT 57.820000  93.200000 74.290000  93.270000 ;
        RECT 57.820000 116.110000 74.290000 116.180000 ;
        RECT 57.820000 139.145000 74.290000 139.215000 ;
        RECT 57.820000 162.160000 74.290000 162.230000 ;
        RECT 57.835000  79.365000 74.290000  79.435000 ;
        RECT 57.835000 102.365000 74.290000 102.435000 ;
        RECT 57.835000 125.365000 74.290000 125.435000 ;
        RECT 57.835000 148.435000 74.290000 148.505000 ;
        RECT 57.845000  27.620000 74.290000  27.690000 ;
        RECT 57.845000 171.365000 74.290000 171.435000 ;
        RECT 57.875000  56.435000 74.290000  56.505000 ;
        RECT 57.890000  47.040000 74.290000  47.110000 ;
        RECT 57.890000  70.070000 74.290000  70.140000 ;
        RECT 57.890000  93.130000 74.290000  93.200000 ;
        RECT 57.890000 116.040000 74.290000 116.110000 ;
        RECT 57.890000 139.075000 74.290000 139.145000 ;
        RECT 57.890000 162.090000 74.290000 162.160000 ;
        RECT 57.905000  79.435000 74.290000  79.505000 ;
        RECT 57.905000 102.435000 74.290000 102.505000 ;
        RECT 57.905000 125.435000 74.290000 125.505000 ;
        RECT 57.905000 148.505000 74.290000 148.575000 ;
        RECT 57.915000  27.690000 74.290000  27.760000 ;
        RECT 57.915000 171.435000 74.290000 171.505000 ;
        RECT 57.945000  56.505000 74.290000  56.575000 ;
        RECT 57.960000  46.970000 74.290000  47.040000 ;
        RECT 57.960000  70.000000 74.290000  70.070000 ;
        RECT 57.960000  93.060000 74.290000  93.130000 ;
        RECT 57.960000 115.970000 74.290000 116.040000 ;
        RECT 57.960000 139.005000 74.290000 139.075000 ;
        RECT 57.960000 162.020000 74.290000 162.090000 ;
        RECT 57.975000  79.505000 74.290000  79.575000 ;
        RECT 57.975000 102.505000 74.290000 102.575000 ;
        RECT 57.975000 125.505000 74.290000 125.575000 ;
        RECT 57.975000 148.575000 74.290000 148.645000 ;
        RECT 57.985000  27.760000 74.290000  27.830000 ;
        RECT 57.985000 171.505000 74.290000 171.575000 ;
        RECT 58.015000  56.575000 74.290000  56.645000 ;
        RECT 58.030000  46.900000 74.290000  46.970000 ;
        RECT 58.030000  69.930000 74.290000  70.000000 ;
        RECT 58.030000  92.990000 74.290000  93.060000 ;
        RECT 58.030000 115.900000 74.290000 115.970000 ;
        RECT 58.030000 138.935000 74.290000 139.005000 ;
        RECT 58.030000 161.950000 74.290000 162.020000 ;
        RECT 58.045000  79.575000 74.290000  79.645000 ;
        RECT 58.045000 102.575000 74.290000 102.645000 ;
        RECT 58.045000 125.575000 74.290000 125.645000 ;
        RECT 58.045000 148.645000 74.290000 148.715000 ;
        RECT 58.055000  27.830000 74.290000  27.900000 ;
        RECT 58.055000 171.575000 74.290000 171.645000 ;
        RECT 58.085000  56.645000 74.290000  56.715000 ;
        RECT 58.100000  46.830000 74.290000  46.900000 ;
        RECT 58.100000  69.860000 74.290000  69.930000 ;
        RECT 58.100000  92.920000 74.290000  92.990000 ;
        RECT 58.100000 115.830000 74.290000 115.900000 ;
        RECT 58.100000 138.865000 74.290000 138.935000 ;
        RECT 58.100000 161.880000 74.290000 161.950000 ;
        RECT 58.115000  79.645000 74.290000  79.715000 ;
        RECT 58.115000 102.645000 74.290000 102.715000 ;
        RECT 58.115000 125.645000 74.290000 125.715000 ;
        RECT 58.115000 148.715000 74.290000 148.785000 ;
        RECT 58.125000  27.900000 74.290000  27.970000 ;
        RECT 58.125000 171.645000 74.290000 171.715000 ;
        RECT 58.155000  56.715000 74.290000  56.785000 ;
        RECT 58.170000  46.760000 74.290000  46.830000 ;
        RECT 58.170000  69.790000 74.290000  69.860000 ;
        RECT 58.170000  92.850000 74.290000  92.920000 ;
        RECT 58.170000 115.760000 74.290000 115.830000 ;
        RECT 58.170000 138.795000 74.290000 138.865000 ;
        RECT 58.170000 161.810000 74.290000 161.880000 ;
        RECT 58.185000  79.715000 74.290000  79.785000 ;
        RECT 58.185000 102.715000 74.290000 102.785000 ;
        RECT 58.185000 125.715000 74.290000 125.785000 ;
        RECT 58.185000 148.785000 74.290000 148.855000 ;
        RECT 58.195000  27.970000 74.290000  28.040000 ;
        RECT 58.195000 171.715000 74.290000 171.785000 ;
        RECT 58.225000  56.785000 74.290000  56.855000 ;
        RECT 58.240000  46.690000 74.290000  46.760000 ;
        RECT 58.240000  69.720000 74.290000  69.790000 ;
        RECT 58.240000  92.780000 74.290000  92.850000 ;
        RECT 58.240000 115.690000 74.290000 115.760000 ;
        RECT 58.240000 138.725000 74.290000 138.795000 ;
        RECT 58.240000 161.740000 74.290000 161.810000 ;
        RECT 58.255000  79.785000 74.290000  79.855000 ;
        RECT 58.255000 102.785000 74.290000 102.855000 ;
        RECT 58.255000 125.785000 74.290000 125.855000 ;
        RECT 58.255000 148.855000 74.290000 148.925000 ;
        RECT 58.265000  28.040000 74.290000  28.110000 ;
        RECT 58.265000 171.785000 74.290000 171.855000 ;
        RECT 58.295000  56.855000 74.290000  56.925000 ;
        RECT 58.310000  46.620000 74.290000  46.690000 ;
        RECT 58.310000  69.650000 74.290000  69.720000 ;
        RECT 58.310000  92.710000 74.290000  92.780000 ;
        RECT 58.310000 115.620000 74.290000 115.690000 ;
        RECT 58.310000 138.655000 74.290000 138.725000 ;
        RECT 58.310000 161.670000 74.290000 161.740000 ;
        RECT 58.325000  79.855000 74.290000  79.925000 ;
        RECT 58.325000 102.855000 74.290000 102.925000 ;
        RECT 58.325000 125.855000 74.290000 125.925000 ;
        RECT 58.325000 148.925000 74.290000 148.995000 ;
        RECT 58.335000  28.110000 74.290000  28.180000 ;
        RECT 58.335000 171.855000 74.290000 171.925000 ;
        RECT 58.365000  56.925000 74.290000  56.995000 ;
        RECT 58.380000  46.550000 74.290000  46.620000 ;
        RECT 58.380000  69.580000 74.290000  69.650000 ;
        RECT 58.380000  92.640000 74.290000  92.710000 ;
        RECT 58.380000 115.550000 74.290000 115.620000 ;
        RECT 58.380000 138.585000 74.290000 138.655000 ;
        RECT 58.380000 161.600000 74.290000 161.670000 ;
        RECT 58.395000  79.925000 74.290000  79.995000 ;
        RECT 58.395000 102.925000 74.290000 102.995000 ;
        RECT 58.395000 125.925000 74.290000 125.995000 ;
        RECT 58.395000 148.995000 74.290000 149.065000 ;
        RECT 58.405000  28.180000 74.290000  28.250000 ;
        RECT 58.405000 171.925000 74.290000 171.995000 ;
        RECT 58.435000  56.995000 74.290000  57.065000 ;
        RECT 58.450000  46.480000 74.290000  46.550000 ;
        RECT 58.450000  69.510000 74.290000  69.580000 ;
        RECT 58.450000  92.570000 74.290000  92.640000 ;
        RECT 58.450000 115.480000 74.290000 115.550000 ;
        RECT 58.450000 138.515000 74.290000 138.585000 ;
        RECT 58.450000 161.530000 74.290000 161.600000 ;
        RECT 58.465000  79.995000 74.290000  80.065000 ;
        RECT 58.465000 102.995000 74.290000 103.065000 ;
        RECT 58.465000 125.995000 74.290000 126.065000 ;
        RECT 58.465000 149.065000 74.290000 149.135000 ;
        RECT 58.475000  28.250000 74.290000  28.320000 ;
        RECT 58.475000 171.995000 74.290000 172.065000 ;
        RECT 58.505000  57.065000 74.290000  57.135000 ;
        RECT 58.520000  46.410000 74.290000  46.480000 ;
        RECT 58.520000  69.440000 74.290000  69.510000 ;
        RECT 58.520000  92.500000 74.290000  92.570000 ;
        RECT 58.520000 115.410000 74.290000 115.480000 ;
        RECT 58.520000 138.445000 74.290000 138.515000 ;
        RECT 58.520000 161.460000 74.290000 161.530000 ;
        RECT 58.535000  80.065000 74.290000  80.135000 ;
        RECT 58.535000 103.065000 74.290000 103.135000 ;
        RECT 58.535000 126.065000 74.290000 126.135000 ;
        RECT 58.535000 149.135000 74.290000 149.205000 ;
        RECT 58.545000  28.320000 74.290000  28.390000 ;
        RECT 58.545000 172.065000 74.290000 172.135000 ;
        RECT 58.575000  57.135000 74.290000  57.205000 ;
        RECT 58.590000  46.340000 74.290000  46.410000 ;
        RECT 58.590000  69.370000 74.290000  69.440000 ;
        RECT 58.590000  92.430000 74.290000  92.500000 ;
        RECT 58.590000 115.340000 74.290000 115.410000 ;
        RECT 58.590000 138.375000 74.290000 138.445000 ;
        RECT 58.590000 161.390000 74.290000 161.460000 ;
        RECT 58.605000  80.135000 74.290000  80.205000 ;
        RECT 58.605000 103.135000 74.290000 103.205000 ;
        RECT 58.605000 126.135000 74.290000 126.205000 ;
        RECT 58.605000 149.205000 74.290000 149.275000 ;
        RECT 58.615000  28.390000 74.290000  28.460000 ;
        RECT 58.615000 172.135000 74.290000 172.205000 ;
        RECT 58.645000  57.205000 74.290000  57.275000 ;
        RECT 58.660000  46.270000 74.290000  46.340000 ;
        RECT 58.660000  69.300000 74.290000  69.370000 ;
        RECT 58.660000  92.360000 74.290000  92.430000 ;
        RECT 58.660000 115.270000 74.290000 115.340000 ;
        RECT 58.660000 138.305000 74.290000 138.375000 ;
        RECT 58.660000 161.320000 74.290000 161.390000 ;
        RECT 58.675000  80.205000 74.290000  80.275000 ;
        RECT 58.675000 103.205000 74.290000 103.275000 ;
        RECT 58.675000 126.205000 74.290000 126.275000 ;
        RECT 58.675000 149.275000 74.290000 149.345000 ;
        RECT 58.685000  28.460000 74.290000  28.530000 ;
        RECT 58.685000 172.205000 74.290000 172.275000 ;
        RECT 58.715000  57.275000 74.290000  57.345000 ;
        RECT 58.730000  46.200000 74.290000  46.270000 ;
        RECT 58.730000  69.230000 74.290000  69.300000 ;
        RECT 58.730000  92.290000 74.290000  92.360000 ;
        RECT 58.730000 115.200000 74.290000 115.270000 ;
        RECT 58.730000 138.235000 74.290000 138.305000 ;
        RECT 58.730000 161.250000 74.290000 161.320000 ;
        RECT 58.730000 185.260000 74.290000 185.295000 ;
        RECT 58.745000  80.275000 74.290000  80.345000 ;
        RECT 58.745000 103.275000 74.290000 103.345000 ;
        RECT 58.745000 126.275000 74.290000 126.345000 ;
        RECT 58.745000 149.345000 74.290000 149.415000 ;
        RECT 58.755000  28.530000 74.290000  28.600000 ;
        RECT 58.755000 172.275000 74.290000 172.345000 ;
        RECT 58.785000  57.345000 74.290000  57.415000 ;
        RECT 58.800000  46.130000 74.290000  46.200000 ;
        RECT 58.800000  69.160000 74.290000  69.230000 ;
        RECT 58.800000  92.220000 74.290000  92.290000 ;
        RECT 58.800000 115.130000 74.290000 115.200000 ;
        RECT 58.800000 138.165000 74.290000 138.235000 ;
        RECT 58.800000 161.180000 74.290000 161.250000 ;
        RECT 58.800000 185.190000 74.290000 185.260000 ;
        RECT 58.815000  80.345000 74.290000  80.415000 ;
        RECT 58.815000 103.345000 74.290000 103.415000 ;
        RECT 58.815000 126.345000 74.290000 126.415000 ;
        RECT 58.815000 149.415000 74.290000 149.485000 ;
        RECT 58.825000  28.600000 74.290000  28.670000 ;
        RECT 58.825000 172.345000 74.290000 172.415000 ;
        RECT 58.855000  57.415000 74.290000  57.485000 ;
        RECT 58.870000  46.060000 74.290000  46.130000 ;
        RECT 58.870000  69.090000 74.290000  69.160000 ;
        RECT 58.870000  92.150000 74.290000  92.220000 ;
        RECT 58.870000 115.060000 74.290000 115.130000 ;
        RECT 58.870000 138.095000 74.290000 138.165000 ;
        RECT 58.870000 161.110000 74.290000 161.180000 ;
        RECT 58.870000 185.120000 74.290000 185.190000 ;
        RECT 58.885000  80.415000 74.290000  80.485000 ;
        RECT 58.885000 103.415000 74.290000 103.485000 ;
        RECT 58.885000 126.415000 74.290000 126.485000 ;
        RECT 58.885000 149.485000 74.290000 149.555000 ;
        RECT 58.895000  28.670000 74.290000  28.740000 ;
        RECT 58.895000 172.415000 74.290000 172.485000 ;
        RECT 58.925000  57.485000 74.290000  57.555000 ;
        RECT 58.940000  45.990000 74.290000  46.060000 ;
        RECT 58.940000  69.020000 74.290000  69.090000 ;
        RECT 58.940000  92.080000 74.290000  92.150000 ;
        RECT 58.940000 114.990000 74.290000 115.060000 ;
        RECT 58.940000 138.025000 74.290000 138.095000 ;
        RECT 58.940000 161.040000 74.290000 161.110000 ;
        RECT 58.940000 185.050000 74.290000 185.120000 ;
        RECT 58.955000  80.485000 74.290000  80.555000 ;
        RECT 58.955000 103.485000 74.290000 103.555000 ;
        RECT 58.955000 126.485000 74.290000 126.555000 ;
        RECT 58.955000 149.555000 74.290000 149.625000 ;
        RECT 58.965000  28.740000 74.290000  28.810000 ;
        RECT 58.965000 172.485000 74.290000 172.555000 ;
        RECT 58.995000  57.555000 74.290000  57.625000 ;
        RECT 59.010000  45.920000 74.290000  45.990000 ;
        RECT 59.010000  68.950000 74.290000  69.020000 ;
        RECT 59.010000  92.010000 74.290000  92.080000 ;
        RECT 59.010000 114.920000 74.290000 114.990000 ;
        RECT 59.010000 137.955000 74.290000 138.025000 ;
        RECT 59.010000 160.970000 74.290000 161.040000 ;
        RECT 59.010000 184.980000 74.290000 185.050000 ;
        RECT 59.025000  80.555000 74.290000  80.625000 ;
        RECT 59.025000 103.555000 74.290000 103.625000 ;
        RECT 59.025000 126.555000 74.290000 126.625000 ;
        RECT 59.025000 149.625000 74.290000 149.695000 ;
        RECT 59.035000  28.810000 74.290000  28.880000 ;
        RECT 59.035000 172.555000 74.290000 172.625000 ;
        RECT 59.065000  57.625000 74.290000  57.695000 ;
        RECT 59.080000  45.850000 74.290000  45.920000 ;
        RECT 59.080000  68.880000 74.290000  68.950000 ;
        RECT 59.080000  91.940000 74.290000  92.010000 ;
        RECT 59.080000 114.850000 74.290000 114.920000 ;
        RECT 59.080000 137.885000 74.290000 137.955000 ;
        RECT 59.080000 160.900000 74.290000 160.970000 ;
        RECT 59.080000 184.910000 74.290000 184.980000 ;
        RECT 59.095000  80.625000 74.290000  80.695000 ;
        RECT 59.095000 103.625000 74.290000 103.695000 ;
        RECT 59.095000 126.625000 74.290000 126.695000 ;
        RECT 59.095000 149.695000 74.290000 149.765000 ;
        RECT 59.105000  28.880000 74.290000  28.950000 ;
        RECT 59.105000 172.625000 74.290000 172.695000 ;
        RECT 59.135000  57.695000 74.290000  57.765000 ;
        RECT 59.150000  45.780000 74.290000  45.850000 ;
        RECT 59.150000  68.810000 74.290000  68.880000 ;
        RECT 59.150000  91.870000 74.290000  91.940000 ;
        RECT 59.150000 114.780000 74.290000 114.850000 ;
        RECT 59.150000 137.815000 74.290000 137.885000 ;
        RECT 59.150000 160.830000 74.290000 160.900000 ;
        RECT 59.150000 184.840000 74.290000 184.910000 ;
        RECT 59.165000  80.695000 74.290000  80.765000 ;
        RECT 59.165000 103.695000 74.290000 103.765000 ;
        RECT 59.165000 126.695000 74.290000 126.765000 ;
        RECT 59.165000 149.765000 74.290000 149.835000 ;
        RECT 59.175000  28.950000 74.290000  29.020000 ;
        RECT 59.175000 172.695000 74.290000 172.765000 ;
        RECT 59.205000  57.765000 74.290000  57.835000 ;
        RECT 59.220000  45.710000 74.290000  45.780000 ;
        RECT 59.220000  68.740000 74.290000  68.810000 ;
        RECT 59.220000  91.800000 74.290000  91.870000 ;
        RECT 59.220000 114.710000 74.290000 114.780000 ;
        RECT 59.220000 137.745000 74.290000 137.815000 ;
        RECT 59.220000 160.760000 74.290000 160.830000 ;
        RECT 59.220000 184.770000 74.290000 184.840000 ;
        RECT 59.235000  80.765000 74.290000  80.835000 ;
        RECT 59.235000 103.765000 74.290000 103.835000 ;
        RECT 59.235000 126.765000 74.290000 126.835000 ;
        RECT 59.235000 149.835000 74.290000 149.905000 ;
        RECT 59.245000  29.020000 74.290000  29.090000 ;
        RECT 59.245000 172.765000 74.290000 172.835000 ;
        RECT 59.275000  57.835000 74.290000  57.905000 ;
        RECT 59.290000  45.640000 74.290000  45.710000 ;
        RECT 59.290000  68.670000 74.290000  68.740000 ;
        RECT 59.290000  91.730000 74.290000  91.800000 ;
        RECT 59.290000 114.640000 74.290000 114.710000 ;
        RECT 59.290000 137.675000 74.290000 137.745000 ;
        RECT 59.290000 160.690000 74.290000 160.760000 ;
        RECT 59.290000 184.700000 74.290000 184.770000 ;
        RECT 59.305000  80.835000 74.290000  80.905000 ;
        RECT 59.305000 103.835000 74.290000 103.905000 ;
        RECT 59.305000 126.835000 74.290000 126.905000 ;
        RECT 59.305000 149.905000 74.290000 149.975000 ;
        RECT 59.315000  29.090000 74.290000  29.160000 ;
        RECT 59.315000 172.835000 74.290000 172.905000 ;
        RECT 59.345000  57.905000 74.290000  57.975000 ;
        RECT 59.360000  45.570000 74.290000  45.640000 ;
        RECT 59.360000  68.600000 74.290000  68.670000 ;
        RECT 59.360000  91.660000 74.290000  91.730000 ;
        RECT 59.360000 114.570000 74.290000 114.640000 ;
        RECT 59.360000 137.605000 74.290000 137.675000 ;
        RECT 59.360000 160.620000 74.290000 160.690000 ;
        RECT 59.360000 184.630000 74.290000 184.700000 ;
        RECT 59.375000  80.905000 74.290000  80.975000 ;
        RECT 59.375000 103.905000 74.290000 103.975000 ;
        RECT 59.375000 126.905000 74.290000 126.975000 ;
        RECT 59.375000 149.975000 74.290000 150.045000 ;
        RECT 59.385000  29.160000 74.290000  29.230000 ;
        RECT 59.385000 172.905000 74.290000 172.975000 ;
        RECT 59.415000  57.975000 74.290000  58.045000 ;
        RECT 59.430000  45.500000 74.290000  45.570000 ;
        RECT 59.430000  68.530000 74.290000  68.600000 ;
        RECT 59.430000  91.590000 74.290000  91.660000 ;
        RECT 59.430000 114.500000 74.290000 114.570000 ;
        RECT 59.430000 137.535000 74.290000 137.605000 ;
        RECT 59.430000 160.550000 74.290000 160.620000 ;
        RECT 59.430000 184.560000 74.290000 184.630000 ;
        RECT 59.445000  80.975000 74.290000  81.045000 ;
        RECT 59.445000 103.975000 74.290000 104.045000 ;
        RECT 59.445000 126.975000 74.290000 127.045000 ;
        RECT 59.445000 150.045000 74.290000 150.115000 ;
        RECT 59.455000  29.230000 74.290000  29.300000 ;
        RECT 59.455000 172.975000 74.290000 173.045000 ;
        RECT 59.485000  58.045000 74.290000  58.115000 ;
        RECT 59.500000  45.430000 74.290000  45.500000 ;
        RECT 59.500000  68.460000 74.290000  68.530000 ;
        RECT 59.500000  91.520000 74.290000  91.590000 ;
        RECT 59.500000 114.430000 74.290000 114.500000 ;
        RECT 59.500000 137.465000 74.290000 137.535000 ;
        RECT 59.500000 160.480000 74.290000 160.550000 ;
        RECT 59.500000 184.490000 74.290000 184.560000 ;
        RECT 59.515000  81.045000 74.290000  81.115000 ;
        RECT 59.515000 104.045000 74.290000 104.115000 ;
        RECT 59.515000 127.045000 74.290000 127.115000 ;
        RECT 59.515000 150.115000 74.290000 150.185000 ;
        RECT 59.525000  29.300000 74.290000  29.370000 ;
        RECT 59.525000 173.045000 74.290000 173.115000 ;
        RECT 59.555000  58.115000 74.290000  58.185000 ;
        RECT 59.570000  45.360000 74.290000  45.430000 ;
        RECT 59.570000  68.390000 74.290000  68.460000 ;
        RECT 59.570000  91.450000 74.290000  91.520000 ;
        RECT 59.570000 114.360000 74.290000 114.430000 ;
        RECT 59.570000 137.395000 74.290000 137.465000 ;
        RECT 59.570000 160.410000 74.290000 160.480000 ;
        RECT 59.570000 184.420000 74.290000 184.490000 ;
        RECT 59.585000  81.115000 74.290000  81.185000 ;
        RECT 59.585000 104.115000 74.290000 104.185000 ;
        RECT 59.585000 127.115000 74.290000 127.185000 ;
        RECT 59.585000 150.185000 74.290000 150.255000 ;
        RECT 59.595000  29.370000 74.290000  29.440000 ;
        RECT 59.595000 173.115000 74.290000 173.185000 ;
        RECT 59.625000  58.185000 74.290000  58.255000 ;
        RECT 59.640000  45.290000 74.290000  45.360000 ;
        RECT 59.640000  68.320000 74.290000  68.390000 ;
        RECT 59.640000  91.380000 74.290000  91.450000 ;
        RECT 59.640000 114.290000 74.290000 114.360000 ;
        RECT 59.640000 137.325000 74.290000 137.395000 ;
        RECT 59.640000 160.340000 74.290000 160.410000 ;
        RECT 59.640000 184.350000 74.290000 184.420000 ;
        RECT 59.655000  81.185000 74.290000  81.255000 ;
        RECT 59.655000 104.185000 74.290000 104.255000 ;
        RECT 59.655000 127.185000 74.290000 127.255000 ;
        RECT 59.655000 150.255000 74.290000 150.325000 ;
        RECT 59.665000  29.440000 74.290000  29.510000 ;
        RECT 59.665000 173.185000 74.290000 173.255000 ;
        RECT 59.695000  58.255000 74.290000  58.325000 ;
        RECT 59.710000  45.220000 74.290000  45.290000 ;
        RECT 59.710000  68.250000 74.290000  68.320000 ;
        RECT 59.710000  91.310000 74.290000  91.380000 ;
        RECT 59.710000 114.220000 74.290000 114.290000 ;
        RECT 59.710000 137.255000 74.290000 137.325000 ;
        RECT 59.710000 160.270000 74.290000 160.340000 ;
        RECT 59.710000 184.280000 74.290000 184.350000 ;
        RECT 59.725000  81.255000 74.290000  81.325000 ;
        RECT 59.725000 104.255000 74.290000 104.325000 ;
        RECT 59.725000 127.255000 74.290000 127.325000 ;
        RECT 59.725000 150.325000 74.290000 150.395000 ;
        RECT 59.735000  29.510000 74.290000  29.580000 ;
        RECT 59.735000 173.255000 74.290000 173.325000 ;
        RECT 59.765000  58.325000 74.290000  58.395000 ;
        RECT 59.780000  45.150000 74.290000  45.220000 ;
        RECT 59.780000  68.180000 74.290000  68.250000 ;
        RECT 59.780000  91.240000 74.290000  91.310000 ;
        RECT 59.780000 114.150000 74.290000 114.220000 ;
        RECT 59.780000 137.185000 74.290000 137.255000 ;
        RECT 59.780000 160.200000 74.290000 160.270000 ;
        RECT 59.780000 184.210000 74.290000 184.280000 ;
        RECT 59.795000  81.325000 74.290000  81.395000 ;
        RECT 59.795000 104.325000 74.290000 104.395000 ;
        RECT 59.795000 127.325000 74.290000 127.395000 ;
        RECT 59.795000 150.395000 74.290000 150.465000 ;
        RECT 59.805000  29.580000 74.290000  29.650000 ;
        RECT 59.805000 173.325000 74.290000 173.395000 ;
        RECT 59.835000  58.395000 74.290000  58.465000 ;
        RECT 59.850000  45.080000 74.290000  45.150000 ;
        RECT 59.850000  68.110000 74.290000  68.180000 ;
        RECT 59.850000  91.170000 74.290000  91.240000 ;
        RECT 59.850000 114.080000 74.290000 114.150000 ;
        RECT 59.850000 137.115000 74.290000 137.185000 ;
        RECT 59.850000 160.130000 74.290000 160.200000 ;
        RECT 59.850000 184.140000 74.290000 184.210000 ;
        RECT 59.865000  81.395000 74.290000  81.465000 ;
        RECT 59.865000 104.395000 74.290000 104.465000 ;
        RECT 59.865000 127.395000 74.290000 127.465000 ;
        RECT 59.865000 150.465000 74.290000 150.535000 ;
        RECT 59.875000  29.650000 74.290000  29.720000 ;
        RECT 59.875000 173.395000 74.290000 173.465000 ;
        RECT 59.905000  58.465000 74.290000  58.535000 ;
        RECT 59.920000  45.010000 74.290000  45.080000 ;
        RECT 59.920000  68.040000 74.290000  68.110000 ;
        RECT 59.920000  91.100000 74.290000  91.170000 ;
        RECT 59.920000 114.010000 74.290000 114.080000 ;
        RECT 59.920000 137.045000 74.290000 137.115000 ;
        RECT 59.920000 160.060000 74.290000 160.130000 ;
        RECT 59.920000 184.070000 74.290000 184.140000 ;
        RECT 59.935000  81.465000 74.290000  81.535000 ;
        RECT 59.935000 104.465000 74.290000 104.535000 ;
        RECT 59.935000 127.465000 74.290000 127.535000 ;
        RECT 59.935000 150.535000 74.290000 150.605000 ;
        RECT 59.945000  29.720000 74.290000  29.790000 ;
        RECT 59.945000 173.465000 74.290000 173.535000 ;
        RECT 59.975000  58.535000 74.290000  58.605000 ;
        RECT 59.990000  44.940000 74.290000  45.010000 ;
        RECT 59.990000  67.970000 74.290000  68.040000 ;
        RECT 59.990000  91.030000 74.290000  91.100000 ;
        RECT 59.990000 113.940000 74.290000 114.010000 ;
        RECT 59.990000 136.975000 74.290000 137.045000 ;
        RECT 59.990000 159.990000 74.290000 160.060000 ;
        RECT 59.990000 184.000000 74.290000 184.070000 ;
        RECT 60.005000  81.535000 74.290000  81.605000 ;
        RECT 60.005000 104.535000 74.290000 104.605000 ;
        RECT 60.005000 127.535000 74.290000 127.605000 ;
        RECT 60.005000 150.605000 74.290000 150.675000 ;
        RECT 60.015000  29.790000 74.290000  29.860000 ;
        RECT 60.015000 173.535000 74.290000 173.605000 ;
        RECT 60.045000  58.605000 74.290000  58.675000 ;
        RECT 60.060000  44.870000 74.290000  44.940000 ;
        RECT 60.060000  67.900000 74.290000  67.970000 ;
        RECT 60.060000  90.960000 74.290000  91.030000 ;
        RECT 60.060000 113.870000 74.290000 113.940000 ;
        RECT 60.060000 136.905000 74.290000 136.975000 ;
        RECT 60.060000 159.920000 74.290000 159.990000 ;
        RECT 60.060000 183.930000 74.290000 184.000000 ;
        RECT 60.075000  81.605000 74.290000  81.675000 ;
        RECT 60.075000 104.605000 74.290000 104.675000 ;
        RECT 60.075000 127.605000 74.290000 127.675000 ;
        RECT 60.075000 150.675000 74.290000 150.745000 ;
        RECT 60.085000  29.860000 74.290000  29.930000 ;
        RECT 60.085000 173.605000 74.290000 173.675000 ;
        RECT 60.115000  58.675000 74.290000  58.745000 ;
        RECT 60.130000  44.800000 74.290000  44.870000 ;
        RECT 60.130000  67.830000 74.290000  67.900000 ;
        RECT 60.130000  90.890000 74.290000  90.960000 ;
        RECT 60.130000 113.800000 74.290000 113.870000 ;
        RECT 60.130000 136.835000 74.290000 136.905000 ;
        RECT 60.130000 159.850000 74.290000 159.920000 ;
        RECT 60.130000 183.860000 74.290000 183.930000 ;
        RECT 60.145000  81.675000 74.290000  81.745000 ;
        RECT 60.145000 104.675000 74.290000 104.745000 ;
        RECT 60.145000 127.675000 74.290000 127.745000 ;
        RECT 60.145000 150.745000 74.290000 150.815000 ;
        RECT 60.155000  29.930000 74.290000  30.000000 ;
        RECT 60.155000 173.675000 74.290000 173.745000 ;
        RECT 60.185000  58.745000 74.290000  58.815000 ;
        RECT 60.200000  44.730000 74.290000  44.800000 ;
        RECT 60.200000  67.760000 74.290000  67.830000 ;
        RECT 60.200000  90.820000 74.290000  90.890000 ;
        RECT 60.200000 113.730000 74.290000 113.800000 ;
        RECT 60.200000 136.765000 74.290000 136.835000 ;
        RECT 60.200000 159.780000 74.290000 159.850000 ;
        RECT 60.200000 183.790000 74.290000 183.860000 ;
        RECT 60.215000  81.745000 74.290000  81.815000 ;
        RECT 60.215000 104.745000 74.290000 104.815000 ;
        RECT 60.215000 127.745000 74.290000 127.815000 ;
        RECT 60.215000 150.815000 74.290000 150.885000 ;
        RECT 60.225000  30.000000 74.290000  30.070000 ;
        RECT 60.225000 173.745000 74.290000 173.815000 ;
        RECT 60.255000  58.815000 74.290000  58.885000 ;
        RECT 60.270000  44.660000 74.290000  44.730000 ;
        RECT 60.270000  67.690000 74.290000  67.760000 ;
        RECT 60.270000  90.750000 74.290000  90.820000 ;
        RECT 60.270000 113.660000 74.290000 113.730000 ;
        RECT 60.270000 136.695000 74.290000 136.765000 ;
        RECT 60.270000 159.710000 74.290000 159.780000 ;
        RECT 60.270000 183.720000 74.290000 183.790000 ;
        RECT 60.285000  81.815000 74.290000  81.885000 ;
        RECT 60.285000 104.815000 74.290000 104.885000 ;
        RECT 60.285000 127.815000 74.290000 127.885000 ;
        RECT 60.285000 150.885000 74.290000 150.955000 ;
        RECT 60.295000  30.070000 74.290000  30.140000 ;
        RECT 60.295000 173.815000 74.290000 173.885000 ;
        RECT 60.325000  58.885000 74.290000  58.955000 ;
        RECT 60.340000  44.590000 74.290000  44.660000 ;
        RECT 60.340000  67.620000 74.290000  67.690000 ;
        RECT 60.340000  90.680000 74.290000  90.750000 ;
        RECT 60.340000 113.590000 74.290000 113.660000 ;
        RECT 60.340000 136.625000 74.290000 136.695000 ;
        RECT 60.340000 159.640000 74.290000 159.710000 ;
        RECT 60.340000 183.650000 74.290000 183.720000 ;
        RECT 60.355000  81.885000 74.290000  81.955000 ;
        RECT 60.355000 104.885000 74.290000 104.955000 ;
        RECT 60.355000 127.885000 74.290000 127.955000 ;
        RECT 60.355000 150.955000 74.290000 151.025000 ;
        RECT 60.365000  30.140000 74.290000  30.210000 ;
        RECT 60.365000 173.885000 74.290000 173.955000 ;
        RECT 60.395000  58.955000 74.290000  59.025000 ;
        RECT 60.410000  44.520000 74.290000  44.590000 ;
        RECT 60.410000  67.550000 74.290000  67.620000 ;
        RECT 60.410000  90.610000 74.290000  90.680000 ;
        RECT 60.410000 113.520000 74.290000 113.590000 ;
        RECT 60.410000 136.555000 74.290000 136.625000 ;
        RECT 60.410000 159.570000 74.290000 159.640000 ;
        RECT 60.410000 183.580000 74.290000 183.650000 ;
        RECT 60.425000  81.955000 74.290000  82.025000 ;
        RECT 60.425000 104.955000 74.290000 105.025000 ;
        RECT 60.425000 127.955000 74.290000 128.025000 ;
        RECT 60.425000 151.025000 74.290000 151.095000 ;
        RECT 60.435000  30.210000 74.290000  30.280000 ;
        RECT 60.435000 173.955000 74.290000 174.025000 ;
        RECT 60.465000  59.025000 74.290000  59.095000 ;
        RECT 60.480000  44.450000 74.290000  44.520000 ;
        RECT 60.480000  67.480000 74.290000  67.550000 ;
        RECT 60.480000  90.540000 74.290000  90.610000 ;
        RECT 60.480000 113.450000 74.290000 113.520000 ;
        RECT 60.480000 136.485000 74.290000 136.555000 ;
        RECT 60.480000 159.500000 74.290000 159.570000 ;
        RECT 60.480000 183.510000 74.290000 183.580000 ;
        RECT 60.495000  82.025000 74.290000  82.095000 ;
        RECT 60.495000 105.025000 74.290000 105.095000 ;
        RECT 60.495000 128.025000 74.290000 128.095000 ;
        RECT 60.495000 151.095000 74.290000 151.165000 ;
        RECT 60.505000  30.280000 74.290000  30.350000 ;
        RECT 60.505000 174.025000 74.290000 174.095000 ;
        RECT 60.535000  59.095000 74.290000  59.165000 ;
        RECT 60.550000  44.380000 74.290000  44.450000 ;
        RECT 60.550000  67.410000 74.290000  67.480000 ;
        RECT 60.550000  90.470000 74.290000  90.540000 ;
        RECT 60.550000 113.380000 74.290000 113.450000 ;
        RECT 60.550000 136.415000 74.290000 136.485000 ;
        RECT 60.550000 159.430000 74.290000 159.500000 ;
        RECT 60.550000 183.440000 74.290000 183.510000 ;
        RECT 60.565000  82.095000 74.290000  82.165000 ;
        RECT 60.565000 105.095000 74.290000 105.165000 ;
        RECT 60.565000 128.095000 74.290000 128.165000 ;
        RECT 60.565000 151.165000 74.290000 151.235000 ;
        RECT 60.575000  30.350000 74.290000  30.420000 ;
        RECT 60.575000 174.095000 74.290000 174.165000 ;
        RECT 60.605000  59.165000 74.290000  59.235000 ;
        RECT 60.620000  44.310000 74.290000  44.380000 ;
        RECT 60.620000  67.340000 74.290000  67.410000 ;
        RECT 60.620000  90.400000 74.290000  90.470000 ;
        RECT 60.620000 113.310000 74.290000 113.380000 ;
        RECT 60.620000 136.345000 74.290000 136.415000 ;
        RECT 60.620000 159.360000 74.290000 159.430000 ;
        RECT 60.620000 183.370000 74.290000 183.440000 ;
        RECT 60.635000  82.165000 74.290000  82.235000 ;
        RECT 60.635000 105.165000 74.290000 105.235000 ;
        RECT 60.635000 128.165000 74.290000 128.235000 ;
        RECT 60.635000 151.235000 74.290000 151.305000 ;
        RECT 60.645000  30.420000 74.290000  30.490000 ;
        RECT 60.645000 174.165000 74.290000 174.235000 ;
        RECT 60.675000  59.235000 74.290000  59.305000 ;
        RECT 60.690000  44.240000 74.290000  44.310000 ;
        RECT 60.690000  67.270000 74.290000  67.340000 ;
        RECT 60.690000  90.330000 74.290000  90.400000 ;
        RECT 60.690000 113.240000 74.290000 113.310000 ;
        RECT 60.690000 136.275000 74.290000 136.345000 ;
        RECT 60.690000 159.290000 74.290000 159.360000 ;
        RECT 60.690000 183.300000 74.290000 183.370000 ;
        RECT 60.705000  82.235000 74.290000  82.305000 ;
        RECT 60.705000 105.235000 74.290000 105.305000 ;
        RECT 60.705000 128.235000 74.290000 128.305000 ;
        RECT 60.705000 151.305000 74.290000 151.375000 ;
        RECT 60.715000  30.490000 74.290000  30.560000 ;
        RECT 60.715000 174.235000 74.290000 174.305000 ;
        RECT 60.745000  59.305000 74.290000  59.375000 ;
        RECT 60.760000  44.170000 74.290000  44.240000 ;
        RECT 60.760000  67.200000 74.290000  67.270000 ;
        RECT 60.760000  90.260000 74.290000  90.330000 ;
        RECT 60.760000 113.170000 74.290000 113.240000 ;
        RECT 60.760000 136.205000 74.290000 136.275000 ;
        RECT 60.760000 159.220000 74.290000 159.290000 ;
        RECT 60.760000 183.230000 74.290000 183.300000 ;
        RECT 60.775000  82.305000 74.290000  82.375000 ;
        RECT 60.775000 105.305000 74.290000 105.375000 ;
        RECT 60.775000 128.305000 74.290000 128.375000 ;
        RECT 60.775000 151.375000 74.290000 151.445000 ;
        RECT 60.785000  30.560000 74.290000  30.630000 ;
        RECT 60.785000 174.305000 74.290000 174.375000 ;
        RECT 60.815000  59.375000 74.290000  59.445000 ;
        RECT 60.830000  44.100000 74.290000  44.170000 ;
        RECT 60.830000  67.130000 74.290000  67.200000 ;
        RECT 60.830000  90.190000 74.290000  90.260000 ;
        RECT 60.830000 113.100000 74.290000 113.170000 ;
        RECT 60.830000 136.135000 74.290000 136.205000 ;
        RECT 60.830000 159.150000 74.290000 159.220000 ;
        RECT 60.830000 183.160000 74.290000 183.230000 ;
        RECT 60.845000  82.375000 74.290000  82.445000 ;
        RECT 60.845000 105.375000 74.290000 105.445000 ;
        RECT 60.845000 128.375000 74.290000 128.445000 ;
        RECT 60.845000 151.445000 74.290000 151.515000 ;
        RECT 60.855000  30.630000 74.290000  30.700000 ;
        RECT 60.855000 174.375000 74.290000 174.445000 ;
        RECT 60.885000  59.445000 74.290000  59.515000 ;
        RECT 60.900000  44.030000 74.290000  44.100000 ;
        RECT 60.900000  67.060000 74.290000  67.130000 ;
        RECT 60.900000  90.120000 74.290000  90.190000 ;
        RECT 60.900000 113.030000 74.290000 113.100000 ;
        RECT 60.900000 136.065000 74.290000 136.135000 ;
        RECT 60.900000 159.080000 74.290000 159.150000 ;
        RECT 60.900000 183.090000 74.290000 183.160000 ;
        RECT 60.915000  82.445000 74.290000  82.515000 ;
        RECT 60.915000 105.445000 74.290000 105.515000 ;
        RECT 60.915000 128.445000 74.290000 128.515000 ;
        RECT 60.915000 151.515000 74.290000 151.585000 ;
        RECT 60.925000  30.700000 74.290000  30.770000 ;
        RECT 60.925000 174.445000 74.290000 174.515000 ;
        RECT 60.955000  59.515000 74.290000  59.585000 ;
        RECT 60.970000  43.960000 74.290000  44.030000 ;
        RECT 60.970000  66.990000 74.290000  67.060000 ;
        RECT 60.970000  90.050000 74.290000  90.120000 ;
        RECT 60.970000 112.960000 74.290000 113.030000 ;
        RECT 60.970000 135.995000 74.290000 136.065000 ;
        RECT 60.970000 159.010000 74.290000 159.080000 ;
        RECT 60.970000 183.020000 74.290000 183.090000 ;
        RECT 60.985000  82.515000 74.290000  82.585000 ;
        RECT 60.985000 105.515000 74.290000 105.585000 ;
        RECT 60.985000 128.515000 74.290000 128.585000 ;
        RECT 60.985000 151.585000 74.290000 151.655000 ;
        RECT 60.995000  30.770000 74.290000  30.840000 ;
        RECT 60.995000 174.515000 74.290000 174.585000 ;
        RECT 61.025000  59.585000 74.290000  59.655000 ;
        RECT 61.040000  43.890000 74.290000  43.960000 ;
        RECT 61.040000  66.920000 74.290000  66.990000 ;
        RECT 61.040000  89.980000 74.290000  90.050000 ;
        RECT 61.040000 112.890000 74.290000 112.960000 ;
        RECT 61.040000 135.925000 74.290000 135.995000 ;
        RECT 61.040000 158.940000 74.290000 159.010000 ;
        RECT 61.040000 182.950000 74.290000 183.020000 ;
        RECT 61.055000  82.585000 74.290000  82.655000 ;
        RECT 61.055000 105.585000 74.290000 105.655000 ;
        RECT 61.055000 128.585000 74.290000 128.655000 ;
        RECT 61.055000 151.655000 74.290000 151.725000 ;
        RECT 61.065000  30.840000 74.290000  30.910000 ;
        RECT 61.065000 174.585000 74.290000 174.655000 ;
        RECT 61.095000  59.655000 74.290000  59.725000 ;
        RECT 61.110000  30.910000 74.290000  30.955000 ;
        RECT 61.110000  30.955000 74.290000  43.820000 ;
        RECT 61.110000  43.820000 74.290000  43.890000 ;
        RECT 61.110000  59.725000 74.290000  59.740000 ;
        RECT 61.110000  59.740000 74.290000  66.850000 ;
        RECT 61.110000  66.850000 74.290000  66.920000 ;
        RECT 61.110000  82.655000 74.290000  82.710000 ;
        RECT 61.110000  82.710000 74.290000  89.910000 ;
        RECT 61.110000  89.910000 74.290000  89.980000 ;
        RECT 61.110000 105.655000 74.290000 105.710000 ;
        RECT 61.110000 105.710000 74.290000 112.820000 ;
        RECT 61.110000 112.820000 74.290000 112.890000 ;
        RECT 61.110000 128.655000 74.290000 128.710000 ;
        RECT 61.110000 128.710000 74.290000 135.855000 ;
        RECT 61.110000 135.855000 74.290000 135.925000 ;
        RECT 61.110000 151.725000 74.290000 151.780000 ;
        RECT 61.110000 151.780000 74.290000 158.870000 ;
        RECT 61.110000 158.870000 74.290000 158.940000 ;
        RECT 61.110000 174.655000 74.290000 174.700000 ;
        RECT 61.110000 174.700000 74.290000 182.880000 ;
        RECT 61.110000 182.880000 74.290000 182.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000   0.000000 48.890000  96.150000 ;
        RECT 37.890000  96.150000 48.890000  96.300000 ;
        RECT 37.890000  96.300000 49.040000  96.450000 ;
        RECT 37.890000  96.450000 49.190000  96.600000 ;
        RECT 37.890000  96.600000 49.340000  96.750000 ;
        RECT 37.890000  96.750000 49.490000  96.900000 ;
        RECT 37.890000  96.900000 49.640000  97.050000 ;
        RECT 37.890000  97.050000 49.790000  97.200000 ;
        RECT 37.890000  97.200000 49.940000  97.350000 ;
        RECT 37.890000  97.350000 50.090000  97.500000 ;
        RECT 37.890000  97.500000 50.240000  97.650000 ;
        RECT 37.890000  97.650000 50.390000  97.800000 ;
        RECT 37.890000  97.800000 50.540000  97.950000 ;
        RECT 37.890000  97.950000 50.690000  98.100000 ;
        RECT 37.890000  98.100000 50.840000  98.250000 ;
        RECT 37.890000  98.250000 50.990000  98.300000 ;
        RECT 37.890000  98.300000 51.040000  99.505000 ;
        RECT 37.890000  99.505000 43.400000  99.655000 ;
        RECT 37.890000  99.655000 43.250000  99.805000 ;
        RECT 37.890000  99.805000 43.100000  99.955000 ;
        RECT 37.890000  99.955000 42.950000 100.105000 ;
        RECT 37.890000 100.105000 42.840000 100.215000 ;
        RECT 37.890000 100.215000 42.840000 102.135000 ;
        RECT 37.890000 102.135000 42.840000 102.285000 ;
        RECT 37.890000 102.285000 42.990000 102.435000 ;
        RECT 37.890000 102.435000 43.140000 102.585000 ;
        RECT 37.890000 102.585000 43.290000 102.735000 ;
        RECT 37.890000 102.735000 43.440000 102.885000 ;
        RECT 37.890000 102.885000 43.590000 103.035000 ;
        RECT 37.890000 103.035000 43.740000 103.185000 ;
        RECT 37.890000 103.185000 43.890000 103.335000 ;
        RECT 37.890000 103.335000 44.040000 103.485000 ;
        RECT 37.890000 103.485000 44.190000 103.635000 ;
        RECT 37.890000 103.635000 44.340000 103.785000 ;
        RECT 37.890000 103.785000 44.490000 103.935000 ;
        RECT 37.890000 103.935000 44.640000 104.085000 ;
        RECT 37.890000 104.085000 44.790000 104.235000 ;
        RECT 37.890000 104.235000 44.940000 104.385000 ;
        RECT 37.890000 104.385000 45.090000 104.535000 ;
        RECT 37.890000 104.535000 45.240000 104.685000 ;
        RECT 37.890000 104.685000 45.390000 104.835000 ;
        RECT 37.890000 104.835000 45.540000 104.985000 ;
        RECT 37.890000 104.985000 45.690000 105.135000 ;
        RECT 37.890000 105.135000 45.840000 105.285000 ;
        RECT 37.890000 105.285000 45.990000 105.435000 ;
        RECT 37.890000 105.435000 46.140000 105.585000 ;
        RECT 37.890000 105.585000 46.290000 105.655000 ;
        RECT 37.965000 175.350000 48.855000 190.020000 ;
        RECT 38.040000 105.655000 46.360000 105.805000 ;
        RECT 38.055000 175.260000 48.855000 175.350000 ;
        RECT 38.190000 105.805000 46.510000 105.955000 ;
        RECT 38.205000 175.110000 48.855000 175.260000 ;
        RECT 38.340000 105.955000 46.660000 106.105000 ;
        RECT 38.355000 174.960000 48.855000 175.110000 ;
        RECT 38.490000 106.105000 46.810000 106.255000 ;
        RECT 38.505000 174.810000 48.855000 174.960000 ;
        RECT 38.640000 106.255000 46.960000 106.405000 ;
        RECT 38.655000 174.660000 48.855000 174.810000 ;
        RECT 38.790000 106.405000 47.110000 106.555000 ;
        RECT 38.805000 174.510000 48.855000 174.660000 ;
        RECT 38.940000 106.555000 47.260000 106.705000 ;
        RECT 38.955000 174.360000 48.855000 174.510000 ;
        RECT 39.090000 106.705000 47.410000 106.855000 ;
        RECT 39.105000 174.210000 48.855000 174.360000 ;
        RECT 39.240000 106.855000 47.560000 107.005000 ;
        RECT 39.255000 174.060000 48.855000 174.210000 ;
        RECT 39.390000 107.005000 47.710000 107.155000 ;
        RECT 39.405000 173.910000 48.855000 174.060000 ;
        RECT 39.540000 107.155000 47.860000 107.305000 ;
        RECT 39.555000 173.760000 48.855000 173.910000 ;
        RECT 39.690000 107.305000 48.010000 107.455000 ;
        RECT 39.705000 173.610000 48.855000 173.760000 ;
        RECT 39.840000 107.455000 48.160000 107.605000 ;
        RECT 39.855000 173.460000 48.855000 173.610000 ;
        RECT 39.990000 107.605000 48.310000 107.755000 ;
        RECT 40.005000 173.310000 48.855000 173.460000 ;
        RECT 40.140000 107.755000 48.460000 107.905000 ;
        RECT 40.155000 173.160000 48.855000 173.310000 ;
        RECT 40.290000 107.905000 48.610000 108.055000 ;
        RECT 40.305000 173.010000 48.855000 173.160000 ;
        RECT 40.385000 108.055000 48.760000 108.150000 ;
        RECT 40.455000 172.860000 48.855000 173.010000 ;
        RECT 40.535000 108.150000 48.855000 108.300000 ;
        RECT 40.605000 172.710000 48.855000 172.860000 ;
        RECT 40.685000 108.300000 48.855000 108.450000 ;
        RECT 40.755000 172.560000 48.855000 172.710000 ;
        RECT 40.835000 108.450000 48.855000 108.600000 ;
        RECT 40.905000 172.410000 48.855000 172.560000 ;
        RECT 40.985000 108.600000 48.855000 108.750000 ;
        RECT 41.055000 172.260000 48.855000 172.410000 ;
        RECT 41.135000 108.750000 48.855000 108.900000 ;
        RECT 41.205000 172.110000 48.855000 172.260000 ;
        RECT 41.285000 108.900000 48.855000 109.050000 ;
        RECT 41.355000 171.960000 48.855000 172.110000 ;
        RECT 41.435000 109.050000 48.855000 109.200000 ;
        RECT 41.505000 171.810000 48.855000 171.960000 ;
        RECT 41.585000 109.200000 48.855000 109.350000 ;
        RECT 41.655000 171.660000 48.855000 171.810000 ;
        RECT 41.735000 109.350000 48.855000 109.500000 ;
        RECT 41.805000 171.510000 48.855000 171.660000 ;
        RECT 41.885000 109.500000 48.855000 109.650000 ;
        RECT 41.955000 171.360000 48.855000 171.510000 ;
        RECT 42.035000 109.650000 48.855000 109.800000 ;
        RECT 42.105000 171.210000 48.855000 171.360000 ;
        RECT 42.185000 109.800000 48.855000 109.950000 ;
        RECT 42.255000 171.060000 48.855000 171.210000 ;
        RECT 42.335000 109.950000 48.855000 110.100000 ;
        RECT 42.405000 170.910000 48.855000 171.060000 ;
        RECT 42.485000 110.100000 48.855000 110.250000 ;
        RECT 42.555000 170.760000 48.855000 170.910000 ;
        RECT 42.635000 110.250000 48.855000 110.400000 ;
        RECT 42.705000 170.610000 48.855000 170.760000 ;
        RECT 42.785000 110.400000 48.855000 110.550000 ;
        RECT 42.855000 110.550000 48.855000 110.620000 ;
        RECT 42.855000 110.620000 48.855000 170.460000 ;
        RECT 42.855000 170.460000 48.855000 170.610000 ;
        RECT 44.655000  99.505000 51.040000  99.610000 ;
        RECT 44.760000  99.610000 51.040000  99.715000 ;
        RECT 44.910000  99.715000 51.040000  99.865000 ;
        RECT 45.060000  99.865000 51.190000 100.015000 ;
        RECT 45.210000 100.015000 51.340000 100.165000 ;
        RECT 45.260000 100.165000 51.490000 100.215000 ;
        RECT 45.260000 100.215000 51.540000 100.365000 ;
        RECT 45.260000 100.365000 51.690000 100.515000 ;
        RECT 45.260000 100.515000 51.840000 100.665000 ;
        RECT 45.260000 100.665000 51.990000 100.815000 ;
        RECT 45.260000 100.815000 52.140000 100.965000 ;
        RECT 45.260000 100.965000 52.290000 101.115000 ;
        RECT 45.260000 101.115000 52.440000 101.265000 ;
        RECT 45.260000 101.265000 52.590000 101.415000 ;
        RECT 45.260000 101.415000 52.740000 101.565000 ;
        RECT 45.260000 101.565000 52.890000 101.715000 ;
        RECT 45.260000 101.715000 53.040000 101.865000 ;
        RECT 45.260000 101.865000 53.190000 102.015000 ;
        RECT 45.260000 102.015000 53.340000 102.165000 ;
        RECT 45.260000 102.165000 53.490000 102.315000 ;
        RECT 45.260000 102.315000 53.640000 102.415000 ;
        RECT 45.410000 102.415000 53.740000 102.565000 ;
        RECT 45.560000 102.565000 53.890000 102.715000 ;
        RECT 45.710000 102.715000 54.040000 102.865000 ;
        RECT 45.860000 102.865000 54.190000 103.015000 ;
        RECT 46.010000 103.015000 54.340000 103.165000 ;
        RECT 46.160000 103.165000 54.490000 103.315000 ;
        RECT 46.310000 103.315000 54.640000 103.465000 ;
        RECT 46.460000 103.465000 54.790000 103.615000 ;
        RECT 46.610000 103.615000 54.940000 103.765000 ;
        RECT 46.760000 103.765000 55.090000 103.915000 ;
        RECT 46.910000 103.915000 55.240000 104.065000 ;
        RECT 47.060000 104.065000 55.390000 104.215000 ;
        RECT 47.210000 104.215000 55.540000 104.365000 ;
        RECT 47.360000 104.365000 55.690000 104.515000 ;
        RECT 47.510000 104.515000 55.840000 104.665000 ;
        RECT 47.660000 104.665000 55.990000 104.815000 ;
        RECT 47.810000 104.815000 56.140000 104.965000 ;
        RECT 47.960000 104.965000 56.290000 105.115000 ;
        RECT 48.110000 105.115000 56.440000 105.265000 ;
        RECT 48.260000 105.265000 56.590000 105.415000 ;
        RECT 48.410000 105.415000 56.740000 105.565000 ;
        RECT 48.560000 105.565000 56.890000 105.715000 ;
        RECT 48.710000 105.715000 57.040000 105.865000 ;
        RECT 48.860000 105.865000 57.190000 106.015000 ;
        RECT 49.010000 106.015000 57.340000 106.165000 ;
        RECT 49.160000 106.165000 57.490000 106.315000 ;
        RECT 49.310000 106.315000 57.640000 106.465000 ;
        RECT 49.460000 106.465000 57.790000 106.615000 ;
        RECT 49.610000 106.615000 57.940000 106.765000 ;
        RECT 49.760000 106.765000 58.090000 106.915000 ;
        RECT 49.775000 172.645000 59.285000 173.020000 ;
        RECT 49.775000 173.020000 59.285000 173.170000 ;
        RECT 49.775000 173.170000 59.435000 173.320000 ;
        RECT 49.775000 173.320000 59.585000 173.470000 ;
        RECT 49.775000 173.470000 59.735000 173.620000 ;
        RECT 49.775000 173.620000 59.885000 173.770000 ;
        RECT 49.775000 173.770000 60.035000 173.920000 ;
        RECT 49.775000 173.920000 60.185000 174.070000 ;
        RECT 49.775000 174.070000 60.335000 174.220000 ;
        RECT 49.775000 174.220000 60.485000 174.370000 ;
        RECT 49.775000 174.370000 60.635000 174.520000 ;
        RECT 49.775000 174.520000 60.785000 174.670000 ;
        RECT 49.775000 174.670000 60.935000 174.680000 ;
        RECT 49.775000 174.680000 60.945000 190.040000 ;
        RECT 49.835000 172.585000 59.285000 172.645000 ;
        RECT 49.910000 106.915000 58.240000 107.065000 ;
        RECT 49.985000 172.435000 59.285000 172.585000 ;
        RECT 50.060000 107.065000 58.390000 107.215000 ;
        RECT 50.135000 172.285000 59.285000 172.435000 ;
        RECT 50.210000 107.215000 58.540000 107.365000 ;
        RECT 50.285000 172.135000 59.285000 172.285000 ;
        RECT 50.360000 107.365000 58.690000 107.515000 ;
        RECT 50.435000 171.985000 59.285000 172.135000 ;
        RECT 50.510000 107.515000 58.840000 107.665000 ;
        RECT 50.585000 171.835000 59.285000 171.985000 ;
        RECT 50.660000 107.665000 58.990000 107.815000 ;
        RECT 50.735000 171.685000 59.285000 171.835000 ;
        RECT 50.805000 107.815000 59.140000 107.960000 ;
        RECT 50.885000 171.535000 59.285000 171.685000 ;
        RECT 50.955000 107.960000 59.285000 108.110000 ;
        RECT 51.035000 171.385000 59.285000 171.535000 ;
        RECT 51.105000 108.110000 59.285000 108.260000 ;
        RECT 51.185000 171.235000 59.285000 171.385000 ;
        RECT 51.255000 108.260000 59.285000 108.410000 ;
        RECT 51.335000 171.085000 59.285000 171.235000 ;
        RECT 51.405000 108.410000 59.285000 108.560000 ;
        RECT 51.485000 170.935000 59.285000 171.085000 ;
        RECT 51.555000 108.560000 59.285000 108.710000 ;
        RECT 51.635000 170.785000 59.285000 170.935000 ;
        RECT 51.705000 108.710000 59.285000 108.860000 ;
        RECT 51.785000 170.635000 59.285000 170.785000 ;
        RECT 51.855000 108.860000 59.285000 109.010000 ;
        RECT 51.935000 170.485000 59.285000 170.635000 ;
        RECT 52.005000 109.010000 59.285000 109.160000 ;
        RECT 52.085000 170.335000 59.285000 170.485000 ;
        RECT 52.155000 109.160000 59.285000 109.310000 ;
        RECT 52.235000 170.185000 59.285000 170.335000 ;
        RECT 52.305000 109.310000 59.285000 109.460000 ;
        RECT 52.385000 170.035000 59.285000 170.185000 ;
        RECT 52.455000 109.460000 59.285000 109.610000 ;
        RECT 52.535000 169.885000 59.285000 170.035000 ;
        RECT 52.605000 109.610000 59.285000 109.760000 ;
        RECT 52.685000 169.735000 59.285000 169.885000 ;
        RECT 52.755000 109.760000 59.285000 109.910000 ;
        RECT 52.835000 169.585000 59.285000 169.735000 ;
        RECT 52.905000 109.910000 59.285000 110.060000 ;
        RECT 52.985000 169.435000 59.285000 169.585000 ;
        RECT 53.055000 110.060000 59.285000 110.210000 ;
        RECT 53.135000 169.285000 59.285000 169.435000 ;
        RECT 53.205000 110.210000 59.285000 110.360000 ;
        RECT 53.285000 110.360000 59.285000 110.440000 ;
        RECT 53.285000 110.440000 59.285000 169.135000 ;
        RECT 53.285000 169.135000 59.285000 169.285000 ;
    END
  END DRN_HVC
  PIN G_CORE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.495000   0.000000 24.395000  36.510000 ;
        RECT 0.495000  46.960000 24.395000  90.500000 ;
        RECT 0.495000  90.500000 24.245000  90.650000 ;
        RECT 0.495000  90.650000 24.095000  90.800000 ;
        RECT 0.495000  90.800000 23.945000  90.950000 ;
        RECT 0.495000  90.950000 23.795000  91.100000 ;
        RECT 0.495000  91.100000 23.645000  91.250000 ;
        RECT 0.495000  91.250000 23.495000  91.400000 ;
        RECT 0.495000  91.400000 23.345000  91.550000 ;
        RECT 0.495000  91.550000 23.195000  91.700000 ;
        RECT 0.495000  91.700000 23.045000  91.850000 ;
        RECT 0.495000  91.850000 22.895000  92.000000 ;
        RECT 0.495000  92.000000 22.745000  92.150000 ;
        RECT 0.495000  92.150000 22.595000  92.300000 ;
        RECT 0.495000  92.300000 22.445000  92.450000 ;
        RECT 0.495000  92.450000 22.295000  92.600000 ;
        RECT 0.495000  92.600000 22.145000  92.750000 ;
        RECT 0.495000  92.750000 21.995000  92.900000 ;
        RECT 0.495000  92.900000 21.845000  93.050000 ;
        RECT 0.495000  93.050000 21.695000  93.200000 ;
        RECT 0.495000  93.200000 21.545000  93.350000 ;
        RECT 0.495000  93.350000 21.395000  93.500000 ;
        RECT 0.495000  93.500000 21.245000  93.650000 ;
        RECT 0.495000  93.650000 21.095000  93.800000 ;
        RECT 0.495000  93.800000 20.945000  93.950000 ;
        RECT 0.495000  93.950000 20.795000  94.100000 ;
        RECT 0.495000  94.100000 20.645000  94.250000 ;
        RECT 0.495000  94.250000 20.495000  94.400000 ;
        RECT 0.495000  94.400000 20.345000  94.550000 ;
        RECT 0.495000  94.550000 20.195000  94.700000 ;
        RECT 0.495000  94.700000 20.045000  94.850000 ;
        RECT 0.495000  94.850000 19.895000  95.000000 ;
        RECT 0.495000  95.000000 19.745000  95.150000 ;
        RECT 0.495000  95.150000 19.595000  95.300000 ;
        RECT 0.495000  95.300000 19.445000  95.450000 ;
        RECT 0.495000  95.450000 19.295000  95.600000 ;
        RECT 0.495000  95.600000 19.145000  95.750000 ;
        RECT 0.495000  95.750000 18.995000  95.900000 ;
        RECT 0.495000  95.900000 18.845000  96.050000 ;
        RECT 0.495000  96.050000 18.695000  96.200000 ;
        RECT 0.495000  96.200000 18.545000  96.350000 ;
        RECT 0.495000  96.350000 18.395000  96.500000 ;
        RECT 0.495000  96.500000 18.245000  96.650000 ;
        RECT 0.495000  96.650000 18.095000  96.800000 ;
        RECT 0.495000  96.800000 17.945000  96.950000 ;
        RECT 0.495000  96.950000 17.795000  97.100000 ;
        RECT 0.495000  97.100000 17.645000  97.250000 ;
        RECT 0.495000  97.250000 17.495000  97.400000 ;
        RECT 0.495000  97.400000 17.345000  97.550000 ;
        RECT 0.495000  97.550000 17.195000  97.700000 ;
        RECT 0.495000  97.700000 17.045000  97.850000 ;
        RECT 0.495000  97.850000 16.895000  98.000000 ;
        RECT 0.495000  98.000000 16.745000  98.150000 ;
        RECT 0.495000  98.150000 16.595000  98.300000 ;
        RECT 0.495000  98.300000 16.445000  98.450000 ;
        RECT 0.495000  98.450000 16.295000  98.600000 ;
        RECT 0.495000  98.600000 16.145000  98.750000 ;
        RECT 0.495000  98.750000 15.995000  98.900000 ;
        RECT 0.495000  98.900000 15.845000  99.050000 ;
        RECT 0.495000  99.050000 15.695000  99.200000 ;
        RECT 0.495000  99.200000 15.545000  99.350000 ;
        RECT 0.495000  99.350000 15.395000  99.500000 ;
        RECT 0.495000  99.500000 15.245000  99.650000 ;
        RECT 0.495000  99.650000 15.095000  99.800000 ;
        RECT 0.495000  99.800000 14.945000  99.950000 ;
        RECT 0.495000  99.950000 14.795000 100.100000 ;
        RECT 0.495000 100.100000 14.645000 100.250000 ;
        RECT 0.495000 100.250000 14.495000 100.400000 ;
        RECT 0.495000 100.400000 14.345000 100.550000 ;
        RECT 0.495000 100.550000 14.195000 100.700000 ;
        RECT 0.495000 100.700000 14.045000 100.850000 ;
        RECT 0.495000 100.850000 13.895000 101.000000 ;
        RECT 0.495000 101.000000 13.745000 101.150000 ;
        RECT 0.495000 101.150000 13.595000 101.300000 ;
        RECT 0.495000 101.300000 13.500000 101.395000 ;
        RECT 0.495000 101.395000 13.500000 173.155000 ;
        RECT 0.520000  46.935000 24.395000  46.960000 ;
        RECT 0.645000  36.510000 24.395000  36.660000 ;
        RECT 0.670000  46.785000 24.395000  46.935000 ;
        RECT 0.795000  36.660000 24.395000  36.810000 ;
        RECT 0.820000  46.635000 24.395000  46.785000 ;
        RECT 0.945000  36.810000 24.395000  36.960000 ;
        RECT 0.970000  36.960000 24.395000  36.985000 ;
        RECT 0.970000  36.985000 24.395000  46.485000 ;
        RECT 0.970000  46.485000 24.395000  46.635000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000   0.000000 74.290000  90.185000 ;
        RECT 50.540000  90.185000 74.290000  90.335000 ;
        RECT 50.690000  90.335000 74.290000  90.485000 ;
        RECT 50.840000  90.485000 74.290000  90.635000 ;
        RECT 50.990000  90.635000 74.290000  90.785000 ;
        RECT 51.140000  90.785000 74.290000  90.935000 ;
        RECT 51.290000  90.935000 74.290000  91.085000 ;
        RECT 51.440000  91.085000 74.290000  91.235000 ;
        RECT 51.590000  91.235000 74.290000  91.385000 ;
        RECT 51.740000  91.385000 74.290000  91.535000 ;
        RECT 51.890000  91.535000 74.290000  91.685000 ;
        RECT 52.040000  91.685000 74.290000  91.835000 ;
        RECT 52.190000  91.835000 74.290000  91.985000 ;
        RECT 52.340000  91.985000 74.290000  92.135000 ;
        RECT 52.490000  92.135000 74.290000  92.285000 ;
        RECT 52.640000  92.285000 74.290000  92.435000 ;
        RECT 52.790000  92.435000 74.290000  92.585000 ;
        RECT 52.940000  92.585000 74.290000  92.735000 ;
        RECT 53.090000  92.735000 74.290000  92.885000 ;
        RECT 53.240000  92.885000 74.290000  93.035000 ;
        RECT 53.390000  93.035000 74.290000  93.185000 ;
        RECT 53.540000  93.185000 74.290000  93.335000 ;
        RECT 53.690000  93.335000 74.290000  93.485000 ;
        RECT 53.840000  93.485000 74.290000  93.635000 ;
        RECT 53.990000  93.635000 74.290000  93.785000 ;
        RECT 54.140000  93.785000 74.290000  93.935000 ;
        RECT 54.290000  93.935000 74.290000  94.085000 ;
        RECT 54.440000  94.085000 74.290000  94.235000 ;
        RECT 54.590000  94.235000 74.290000  94.385000 ;
        RECT 54.740000  94.385000 74.290000  94.535000 ;
        RECT 54.890000  94.535000 74.290000  94.685000 ;
        RECT 55.040000  94.685000 74.290000  94.835000 ;
        RECT 55.190000  94.835000 74.290000  94.985000 ;
        RECT 55.340000  94.985000 74.290000  95.135000 ;
        RECT 55.490000  95.135000 74.290000  95.285000 ;
        RECT 55.640000  95.285000 74.290000  95.435000 ;
        RECT 55.790000  95.435000 74.290000  95.585000 ;
        RECT 55.940000  95.585000 74.290000  95.735000 ;
        RECT 56.090000  95.735000 74.290000  95.885000 ;
        RECT 56.240000  95.885000 74.290000  96.035000 ;
        RECT 56.390000  96.035000 74.290000  96.185000 ;
        RECT 56.540000  96.185000 74.290000  96.335000 ;
        RECT 56.690000  96.335000 74.290000  96.485000 ;
        RECT 56.840000  96.485000 74.290000  96.635000 ;
        RECT 56.990000  96.635000 74.290000  96.785000 ;
        RECT 57.140000  96.785000 74.290000  96.935000 ;
        RECT 57.290000  96.935000 74.290000  97.085000 ;
        RECT 57.440000  97.085000 74.290000  97.235000 ;
        RECT 57.590000  97.235000 74.290000  97.385000 ;
        RECT 57.740000  97.385000 74.290000  97.535000 ;
        RECT 57.890000  97.535000 74.290000  97.685000 ;
        RECT 58.040000  97.685000 74.290000  97.835000 ;
        RECT 58.190000  97.835000 74.290000  97.985000 ;
        RECT 58.340000  97.985000 74.290000  98.135000 ;
        RECT 58.490000  98.135000 74.290000  98.285000 ;
        RECT 58.640000  98.285000 74.290000  98.435000 ;
        RECT 58.790000  98.435000 74.290000  98.585000 ;
        RECT 58.940000  98.585000 74.290000  98.735000 ;
        RECT 59.090000  98.735000 74.290000  98.885000 ;
        RECT 59.240000  98.885000 74.290000  99.035000 ;
        RECT 59.390000  99.035000 74.290000  99.185000 ;
        RECT 59.540000  99.185000 74.290000  99.335000 ;
        RECT 59.690000  99.335000 74.290000  99.485000 ;
        RECT 59.840000  99.485000 74.290000  99.635000 ;
        RECT 59.990000  99.635000 74.290000  99.785000 ;
        RECT 60.140000  99.785000 74.290000  99.935000 ;
        RECT 60.290000  99.935000 74.290000 100.085000 ;
        RECT 60.440000 100.085000 74.290000 100.235000 ;
        RECT 60.590000 100.235000 74.290000 100.385000 ;
        RECT 60.740000 100.385000 74.290000 100.535000 ;
        RECT 60.890000 100.535000 74.290000 100.685000 ;
        RECT 61.040000 100.685000 74.290000 100.835000 ;
        RECT 61.190000 100.835000 74.290000 100.985000 ;
        RECT 61.340000 100.985000 74.290000 101.135000 ;
        RECT 61.490000 101.135000 74.290000 101.285000 ;
        RECT 61.500000 101.285000 74.290000 101.295000 ;
        RECT 61.500000 101.295000 74.290000 173.320000 ;
    END
  END G_CORE
  PIN OGC_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 25.895000 0.000000 27.895000 0.535000 ;
    END
  END OGC_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT  0.495000   0.000000 24.395000   2.055000 ;
        RECT  0.565000   2.055000 24.395000   2.125000 ;
        RECT  0.635000   2.125000 24.395000   2.195000 ;
        RECT  0.705000   2.195000 24.395000   2.265000 ;
        RECT  0.775000   2.265000 24.395000   2.335000 ;
        RECT  0.845000   2.335000 24.395000   2.405000 ;
        RECT  0.915000   2.405000 24.395000   2.475000 ;
        RECT  0.985000   2.475000 24.395000   2.545000 ;
        RECT  1.005000   2.545000 24.395000   2.565000 ;
        RECT  1.005000   2.565000 24.395000   8.595000 ;
        RECT  1.005000   8.595000 24.395000   8.665000 ;
        RECT  1.005000   8.665000 24.465000   8.735000 ;
        RECT  1.005000   8.735000 24.535000   8.805000 ;
        RECT  1.005000   8.805000 24.605000   8.875000 ;
        RECT  1.005000   8.875000 24.675000   8.945000 ;
        RECT  1.005000   8.945000 24.745000   9.015000 ;
        RECT  1.005000   9.015000 24.815000   9.085000 ;
        RECT  1.005000   9.085000 24.885000   9.155000 ;
        RECT  1.005000   9.155000 24.955000   9.225000 ;
        RECT  1.005000   9.225000 25.025000   9.295000 ;
        RECT  1.005000   9.295000 25.095000   9.365000 ;
        RECT  1.005000   9.365000 25.165000   9.435000 ;
        RECT  1.005000   9.435000 25.235000   9.505000 ;
        RECT  1.005000   9.505000 25.305000   9.575000 ;
        RECT  1.005000   9.575000 25.375000   9.645000 ;
        RECT  1.005000   9.645000 25.445000   9.715000 ;
        RECT  1.005000   9.715000 25.515000   9.785000 ;
        RECT  1.005000   9.785000 25.585000   9.855000 ;
        RECT  1.005000   9.855000 25.655000   9.925000 ;
        RECT  1.005000   9.925000 25.725000   9.995000 ;
        RECT  1.005000   9.995000 25.795000  10.065000 ;
        RECT  1.005000  10.065000 25.865000  10.135000 ;
        RECT  1.005000  10.135000 25.935000  10.205000 ;
        RECT  1.005000  10.205000 26.005000  10.275000 ;
        RECT  1.005000  10.275000 26.075000  10.345000 ;
        RECT  1.005000  10.345000 26.145000  10.415000 ;
        RECT  1.005000  10.415000 26.215000  10.485000 ;
        RECT  1.005000  10.485000 26.285000  10.555000 ;
        RECT  1.005000  10.555000 26.355000  10.625000 ;
        RECT  1.005000  10.625000 26.425000  10.695000 ;
        RECT  1.005000  10.695000 26.495000  10.765000 ;
        RECT  1.005000  10.765000 26.565000  10.835000 ;
        RECT  1.005000  10.835000 26.635000  10.905000 ;
        RECT  1.005000  10.905000 26.705000  10.975000 ;
        RECT  1.005000  10.975000 26.775000  11.045000 ;
        RECT  1.005000  11.045000 26.845000  11.115000 ;
        RECT  1.005000  11.115000 26.915000  11.185000 ;
        RECT  1.005000  11.185000 26.985000  11.255000 ;
        RECT  1.005000  11.255000 27.055000  11.325000 ;
        RECT  1.005000  11.325000 27.125000  11.395000 ;
        RECT  1.005000  11.395000 27.195000  11.465000 ;
        RECT  1.005000  11.465000 27.265000  11.535000 ;
        RECT  1.005000  11.535000 27.335000  11.605000 ;
        RECT  1.005000  11.605000 27.405000  11.675000 ;
        RECT  1.005000  11.675000 27.475000  11.745000 ;
        RECT  1.005000  11.745000 27.545000  11.815000 ;
        RECT  1.005000  11.815000 27.615000  11.885000 ;
        RECT  1.005000  11.885000 27.685000  11.955000 ;
        RECT  1.005000  11.955000 27.755000  12.025000 ;
        RECT  1.005000  12.025000 27.825000  12.095000 ;
        RECT  1.005000  12.095000 27.895000  12.165000 ;
        RECT  1.005000  12.165000 27.965000  12.235000 ;
        RECT  1.005000  12.235000 28.035000  12.305000 ;
        RECT  1.005000  12.305000 28.105000  12.375000 ;
        RECT  1.005000  12.375000 28.175000  12.400000 ;
        RECT  1.005000  12.400000 36.895000  25.700000 ;
        RECT  1.005000  25.700000 18.750000  25.770000 ;
        RECT  1.005000  25.770000 18.680000  25.840000 ;
        RECT  1.005000  25.840000 18.610000  25.910000 ;
        RECT  1.005000  25.910000 18.540000  25.980000 ;
        RECT  1.005000  25.980000 18.470000  26.050000 ;
        RECT  1.005000  26.050000 18.400000  26.120000 ;
        RECT  1.005000  26.120000 18.330000  26.190000 ;
        RECT  1.005000  26.190000 18.260000  26.260000 ;
        RECT  1.005000  26.260000 18.190000  26.330000 ;
        RECT  1.005000  26.330000 18.120000  26.400000 ;
        RECT  1.005000  26.400000 18.050000  26.470000 ;
        RECT  1.005000  26.470000 17.980000  26.540000 ;
        RECT  1.005000  26.540000 17.910000  26.610000 ;
        RECT  1.005000  26.610000 17.840000  26.680000 ;
        RECT  1.005000  26.680000 17.770000  26.750000 ;
        RECT  1.005000  26.750000 17.700000  26.820000 ;
        RECT  1.005000  26.820000 17.630000  26.890000 ;
        RECT  1.005000  26.890000 17.560000  26.960000 ;
        RECT  1.005000  26.960000 17.490000  27.030000 ;
        RECT  1.005000  27.030000 17.420000  27.100000 ;
        RECT  1.005000  27.100000 17.350000  27.170000 ;
        RECT  1.005000  27.170000 17.280000  27.240000 ;
        RECT  1.005000  27.240000 17.210000  27.310000 ;
        RECT  1.005000  27.310000 17.140000  27.380000 ;
        RECT  1.005000  27.380000 17.070000  27.450000 ;
        RECT  1.005000  27.450000 17.000000  27.520000 ;
        RECT  1.005000  27.520000 16.930000  27.590000 ;
        RECT  1.005000  27.590000 16.860000  27.660000 ;
        RECT  1.005000  27.660000 16.790000  27.730000 ;
        RECT  1.005000  27.730000 16.720000  27.800000 ;
        RECT  1.005000  27.800000 16.650000  27.870000 ;
        RECT  1.005000  27.870000 16.580000  27.940000 ;
        RECT  1.005000  27.940000 16.510000  28.010000 ;
        RECT  1.005000  28.010000 16.440000  28.080000 ;
        RECT  1.005000  28.080000 16.370000  28.150000 ;
        RECT  1.005000  28.150000 16.300000  28.220000 ;
        RECT  1.005000  28.220000 16.230000  28.290000 ;
        RECT  1.005000  28.290000 16.160000  28.360000 ;
        RECT  1.005000  28.360000 16.090000  28.430000 ;
        RECT  1.005000  28.430000 16.020000  28.500000 ;
        RECT  1.005000  28.500000 15.950000  28.570000 ;
        RECT  1.005000  28.570000 15.880000  28.640000 ;
        RECT  1.005000  28.640000 15.810000  28.710000 ;
        RECT  1.005000  28.710000 15.740000  28.780000 ;
        RECT  1.005000  28.780000 15.670000  28.850000 ;
        RECT  1.005000  28.850000 15.600000  28.920000 ;
        RECT  1.005000  28.920000 15.530000  28.990000 ;
        RECT  1.005000  28.990000 15.460000  29.060000 ;
        RECT  1.005000  29.060000 15.390000  29.130000 ;
        RECT  1.005000  29.130000 15.320000  29.200000 ;
        RECT  1.005000  29.200000 15.250000  29.270000 ;
        RECT  1.005000  29.270000 15.205000  29.315000 ;
        RECT  1.005000  29.315000 15.205000  35.665000 ;
        RECT  1.005000  35.665000 15.205000  35.735000 ;
        RECT  1.005000  35.735000 15.275000  35.805000 ;
        RECT  1.005000  35.805000 15.345000  35.875000 ;
        RECT  1.005000  35.875000 15.415000  35.945000 ;
        RECT  1.005000  35.945000 15.485000  36.015000 ;
        RECT  1.005000  36.015000 15.555000  36.085000 ;
        RECT  1.005000  36.085000 15.625000  36.155000 ;
        RECT  1.005000  36.155000 15.695000  36.225000 ;
        RECT  1.005000  36.225000 15.765000  36.295000 ;
        RECT  1.005000  36.295000 15.835000  36.365000 ;
        RECT  1.005000  36.365000 15.905000  36.435000 ;
        RECT  1.005000  36.435000 15.975000  36.505000 ;
        RECT  1.005000  36.505000 16.045000  36.575000 ;
        RECT  1.005000  36.575000 16.115000  36.640000 ;
        RECT  1.005000  47.130000 14.120000  54.215000 ;
        RECT  1.005000  54.215000 14.120000  54.285000 ;
        RECT  1.005000  54.285000 14.190000  54.355000 ;
        RECT  1.005000  54.355000 14.260000  54.425000 ;
        RECT  1.005000  54.425000 14.330000  54.495000 ;
        RECT  1.005000  54.495000 14.400000  54.565000 ;
        RECT  1.005000  54.565000 14.470000  54.635000 ;
        RECT  1.005000  54.635000 14.540000  54.705000 ;
        RECT  1.005000  54.705000 14.610000  54.775000 ;
        RECT  1.005000  54.775000 14.680000  54.845000 ;
        RECT  1.005000  54.845000 14.750000  54.915000 ;
        RECT  1.005000  54.915000 14.820000  54.985000 ;
        RECT  1.005000  54.985000 14.890000  55.055000 ;
        RECT  1.005000  55.055000 14.960000  55.125000 ;
        RECT  1.005000  55.125000 15.030000  55.195000 ;
        RECT  1.005000  55.195000 15.100000  55.265000 ;
        RECT  1.005000  55.265000 15.170000  55.335000 ;
        RECT  1.005000  55.335000 15.240000  55.405000 ;
        RECT  1.005000  55.405000 15.310000  55.475000 ;
        RECT  1.005000  55.475000 15.380000  55.545000 ;
        RECT  1.005000  55.545000 15.450000  55.615000 ;
        RECT  1.005000  55.615000 15.520000  55.685000 ;
        RECT  1.005000  55.685000 15.590000  55.755000 ;
        RECT  1.005000  55.755000 15.660000  55.825000 ;
        RECT  1.005000  55.825000 15.730000  55.895000 ;
        RECT  1.005000  55.895000 15.800000  55.965000 ;
        RECT  1.005000  55.965000 15.870000  56.035000 ;
        RECT  1.005000  56.035000 15.940000  56.105000 ;
        RECT  1.005000  56.105000 16.010000  56.175000 ;
        RECT  1.005000  56.175000 16.080000  56.245000 ;
        RECT  1.005000  56.245000 16.150000  56.315000 ;
        RECT  1.005000  56.315000 16.220000  56.385000 ;
        RECT  1.005000  56.385000 16.290000  56.455000 ;
        RECT  1.005000  56.455000 16.360000  56.525000 ;
        RECT  1.005000  56.525000 16.430000  56.595000 ;
        RECT  1.005000  56.595000 16.500000  56.665000 ;
        RECT  1.005000  56.665000 16.570000  56.735000 ;
        RECT  1.005000  56.735000 16.640000  56.805000 ;
        RECT  1.005000  56.805000 16.710000  56.875000 ;
        RECT  1.005000  56.875000 16.780000  56.945000 ;
        RECT  1.005000  56.945000 16.850000  57.015000 ;
        RECT  1.005000  57.015000 16.920000  57.085000 ;
        RECT  1.005000  57.085000 16.990000  57.155000 ;
        RECT  1.005000  57.155000 17.060000  57.225000 ;
        RECT  1.005000  57.225000 17.130000  57.295000 ;
        RECT  1.005000  57.295000 17.200000  57.365000 ;
        RECT  1.005000  57.365000 17.270000  57.435000 ;
        RECT  1.005000  57.435000 17.340000  57.505000 ;
        RECT  1.005000  57.505000 17.410000  57.575000 ;
        RECT  1.005000  57.575000 17.480000  57.645000 ;
        RECT  1.005000  57.645000 17.550000  57.715000 ;
        RECT  1.005000  57.715000 17.620000  57.780000 ;
        RECT  1.005000  57.780000 56.710000  66.480000 ;
        RECT  1.005000  66.480000 17.595000  66.550000 ;
        RECT  1.005000  66.550000 17.525000  66.620000 ;
        RECT  1.005000  66.620000 17.455000  66.690000 ;
        RECT  1.005000  66.690000 17.385000  66.760000 ;
        RECT  1.005000  66.760000 17.315000  66.830000 ;
        RECT  1.005000  66.830000 17.245000  66.900000 ;
        RECT  1.005000  66.900000 17.175000  66.970000 ;
        RECT  1.005000  66.970000 17.105000  67.040000 ;
        RECT  1.005000  67.040000 17.035000  67.110000 ;
        RECT  1.005000  67.110000 16.965000  67.180000 ;
        RECT  1.005000  67.180000 16.895000  67.250000 ;
        RECT  1.005000  67.250000 16.825000  67.320000 ;
        RECT  1.005000  67.320000 16.755000  67.390000 ;
        RECT  1.005000  67.390000 16.685000  67.460000 ;
        RECT  1.005000  67.460000 16.615000  67.530000 ;
        RECT  1.005000  67.530000 16.545000  67.600000 ;
        RECT  1.005000  67.600000 16.475000  67.670000 ;
        RECT  1.005000  67.670000 16.405000  67.740000 ;
        RECT  1.005000  67.740000 16.335000  67.810000 ;
        RECT  1.005000  67.810000 16.265000  67.880000 ;
        RECT  1.005000  67.880000 16.195000  67.950000 ;
        RECT  1.005000  67.950000 16.125000  68.020000 ;
        RECT  1.005000  68.020000 16.055000  68.090000 ;
        RECT  1.005000  68.090000 15.985000  68.160000 ;
        RECT  1.005000  68.160000 15.915000  68.230000 ;
        RECT  1.005000  68.230000 15.845000  68.300000 ;
        RECT  1.005000  68.300000 15.775000  68.370000 ;
        RECT  1.005000  68.370000 15.705000  68.440000 ;
        RECT  1.005000  68.440000 15.635000  68.510000 ;
        RECT  1.005000  68.510000 15.565000  68.580000 ;
        RECT  1.005000  68.580000 15.495000  68.650000 ;
        RECT  1.005000  68.650000 15.425000  68.720000 ;
        RECT  1.005000  68.720000 15.355000  68.790000 ;
        RECT  1.005000  68.790000 15.285000  68.860000 ;
        RECT  1.005000  68.860000 15.215000  68.930000 ;
        RECT  1.005000  68.930000 15.145000  69.000000 ;
        RECT  1.005000  69.000000 15.075000  69.070000 ;
        RECT  1.005000  69.070000 15.005000  69.140000 ;
        RECT  1.005000  69.140000 14.935000  69.210000 ;
        RECT  1.005000  69.210000 14.865000  69.280000 ;
        RECT  1.005000  69.280000 14.795000  69.350000 ;
        RECT  1.005000  69.350000 14.725000  69.420000 ;
        RECT  1.005000  69.420000 14.655000  69.490000 ;
        RECT  1.005000  69.490000 14.585000  69.560000 ;
        RECT  1.005000  69.560000 14.515000  69.630000 ;
        RECT  1.005000  69.630000 14.445000  69.700000 ;
        RECT  1.005000  69.700000 14.375000  69.770000 ;
        RECT  1.005000  69.770000 14.305000  69.840000 ;
        RECT  1.005000  69.840000 14.235000  69.910000 ;
        RECT  1.005000  69.910000 14.165000  69.980000 ;
        RECT  1.005000  69.980000 14.120000  70.025000 ;
        RECT  1.005000  70.025000 14.120000  77.240000 ;
        RECT  1.005000  77.240000 14.120000  77.310000 ;
        RECT  1.005000  77.310000 14.190000  77.380000 ;
        RECT  1.005000  77.380000 14.260000  77.450000 ;
        RECT  1.005000  77.450000 14.330000  77.520000 ;
        RECT  1.005000  77.520000 14.400000  77.590000 ;
        RECT  1.005000  77.590000 14.470000  77.660000 ;
        RECT  1.005000  77.660000 14.540000  77.730000 ;
        RECT  1.005000  77.730000 14.610000  77.800000 ;
        RECT  1.005000  77.800000 14.680000  77.870000 ;
        RECT  1.005000  77.870000 14.750000  77.940000 ;
        RECT  1.005000  77.940000 14.820000  78.010000 ;
        RECT  1.005000  78.010000 14.890000  78.080000 ;
        RECT  1.005000  78.080000 14.960000  78.150000 ;
        RECT  1.005000  78.150000 15.030000  78.220000 ;
        RECT  1.005000  78.220000 15.100000  78.290000 ;
        RECT  1.005000  78.290000 15.170000  78.360000 ;
        RECT  1.005000  78.360000 15.240000  78.430000 ;
        RECT  1.005000  78.430000 15.310000  78.500000 ;
        RECT  1.005000  78.500000 15.380000  78.570000 ;
        RECT  1.005000  78.570000 15.450000  78.640000 ;
        RECT  1.005000  78.640000 15.520000  78.710000 ;
        RECT  1.005000  78.710000 15.590000  78.780000 ;
        RECT  1.005000  78.780000 15.660000  78.850000 ;
        RECT  1.005000  78.850000 15.730000  78.920000 ;
        RECT  1.005000  78.920000 15.800000  78.990000 ;
        RECT  1.005000  78.990000 15.870000  79.060000 ;
        RECT  1.005000  79.060000 15.940000  79.130000 ;
        RECT  1.005000  79.130000 16.010000  79.200000 ;
        RECT  1.005000  79.200000 16.080000  79.270000 ;
        RECT  1.005000  79.270000 16.150000  79.340000 ;
        RECT  1.005000  79.340000 16.220000  79.410000 ;
        RECT  1.005000  79.410000 16.290000  79.480000 ;
        RECT  1.005000  79.480000 16.360000  79.550000 ;
        RECT  1.005000  79.550000 16.430000  79.620000 ;
        RECT  1.005000  79.620000 16.500000  79.690000 ;
        RECT  1.005000  79.690000 16.570000  79.760000 ;
        RECT  1.005000  79.760000 16.640000  79.830000 ;
        RECT  1.005000  79.830000 16.710000  79.900000 ;
        RECT  1.005000  79.900000 16.780000  79.970000 ;
        RECT  1.005000  79.970000 16.850000  80.040000 ;
        RECT  1.005000  80.040000 16.920000  80.110000 ;
        RECT  1.005000  80.110000 16.990000  80.180000 ;
        RECT  1.005000  80.180000 17.060000  80.250000 ;
        RECT  1.005000  80.250000 17.130000  80.320000 ;
        RECT  1.005000  80.320000 17.200000  80.390000 ;
        RECT  1.005000  80.390000 17.270000  80.460000 ;
        RECT  1.005000  80.460000 17.340000  80.530000 ;
        RECT  1.005000  80.530000 17.410000  80.600000 ;
        RECT  1.005000  80.600000 17.480000  80.670000 ;
        RECT  1.005000  80.670000 17.550000  80.740000 ;
        RECT  1.005000  80.740000 17.620000  80.780000 ;
        RECT  1.005000  80.780000 56.705000  89.480000 ;
        RECT  1.005000  89.480000 17.595000  89.550000 ;
        RECT  1.005000  89.550000 17.525000  89.620000 ;
        RECT  1.005000  89.620000 17.455000  89.690000 ;
        RECT  1.005000  89.690000 17.385000  89.760000 ;
        RECT  1.005000  89.760000 17.315000  89.830000 ;
        RECT  1.005000  89.830000 17.245000  89.900000 ;
        RECT  1.005000  89.900000 17.175000  89.970000 ;
        RECT  1.005000  89.970000 17.105000  90.040000 ;
        RECT  1.005000  90.040000 17.035000  90.110000 ;
        RECT  1.005000  90.110000 16.965000  90.180000 ;
        RECT  1.005000  90.180000 16.895000  90.250000 ;
        RECT  1.005000  90.250000 16.825000  90.320000 ;
        RECT  1.005000  90.320000 16.755000  90.390000 ;
        RECT  1.005000  90.390000 16.685000  90.460000 ;
        RECT  1.005000  90.460000 16.615000  90.530000 ;
        RECT  1.005000  90.530000 16.545000  90.600000 ;
        RECT  1.005000  90.600000 16.475000  90.670000 ;
        RECT  1.005000  90.670000 16.405000  90.740000 ;
        RECT  1.005000  90.740000 16.335000  90.810000 ;
        RECT  1.005000  90.810000 16.265000  90.880000 ;
        RECT  1.005000  90.880000 16.195000  90.950000 ;
        RECT  1.005000  90.950000 16.125000  91.020000 ;
        RECT  1.005000  91.020000 16.055000  91.090000 ;
        RECT  1.005000  91.090000 15.985000  91.160000 ;
        RECT  1.005000  91.160000 15.915000  91.230000 ;
        RECT  1.005000  91.230000 15.845000  91.300000 ;
        RECT  1.005000  91.300000 15.775000  91.370000 ;
        RECT  1.005000  91.370000 15.705000  91.440000 ;
        RECT  1.005000  91.440000 15.635000  91.510000 ;
        RECT  1.005000  91.510000 15.565000  91.580000 ;
        RECT  1.005000  91.580000 15.495000  91.650000 ;
        RECT  1.005000  91.650000 15.425000  91.720000 ;
        RECT  1.005000  91.720000 15.355000  91.790000 ;
        RECT  1.005000  91.790000 15.285000  91.860000 ;
        RECT  1.005000  91.860000 15.215000  91.930000 ;
        RECT  1.005000  91.930000 15.145000  92.000000 ;
        RECT  1.005000  92.000000 15.075000  92.070000 ;
        RECT  1.005000  92.070000 15.005000  92.140000 ;
        RECT  1.005000  92.140000 14.935000  92.210000 ;
        RECT  1.005000  92.210000 14.865000  92.280000 ;
        RECT  1.005000  92.280000 14.795000  92.350000 ;
        RECT  1.005000  92.350000 14.725000  92.420000 ;
        RECT  1.005000  92.420000 14.655000  92.490000 ;
        RECT  1.005000  92.490000 14.585000  92.560000 ;
        RECT  1.005000  92.560000 14.515000  92.630000 ;
        RECT  1.005000  92.630000 14.445000  92.700000 ;
        RECT  1.005000  92.700000 14.375000  92.770000 ;
        RECT  1.005000  92.770000 14.305000  92.840000 ;
        RECT  1.005000  92.840000 14.235000  92.910000 ;
        RECT  1.005000  92.910000 14.165000  92.980000 ;
        RECT  1.005000  92.980000 14.120000  93.025000 ;
        RECT  1.005000  93.025000 14.120000 100.240000 ;
        RECT  1.005000 100.240000 14.120000 100.310000 ;
        RECT  1.005000 100.310000 14.190000 100.380000 ;
        RECT  1.005000 100.380000 14.260000 100.450000 ;
        RECT  1.005000 100.450000 14.330000 100.520000 ;
        RECT  1.005000 100.520000 14.400000 100.590000 ;
        RECT  1.005000 100.590000 14.470000 100.660000 ;
        RECT  1.005000 100.660000 14.540000 100.730000 ;
        RECT  1.005000 100.730000 14.610000 100.800000 ;
        RECT  1.005000 100.800000 14.680000 100.870000 ;
        RECT  1.005000 100.870000 14.750000 100.940000 ;
        RECT  1.005000 100.940000 14.820000 101.010000 ;
        RECT  1.005000 101.010000 14.890000 101.080000 ;
        RECT  1.005000 101.080000 14.960000 101.150000 ;
        RECT  1.005000 101.150000 15.030000 101.220000 ;
        RECT  1.005000 101.220000 15.100000 101.290000 ;
        RECT  1.005000 101.290000 15.170000 101.360000 ;
        RECT  1.005000 101.360000 15.240000 101.430000 ;
        RECT  1.005000 101.430000 15.310000 101.500000 ;
        RECT  1.005000 101.500000 15.380000 101.570000 ;
        RECT  1.005000 101.570000 15.450000 101.640000 ;
        RECT  1.005000 101.640000 15.520000 101.710000 ;
        RECT  1.005000 101.710000 15.590000 101.780000 ;
        RECT  1.005000 101.780000 15.660000 101.850000 ;
        RECT  1.005000 101.850000 15.730000 101.920000 ;
        RECT  1.005000 101.920000 15.800000 101.990000 ;
        RECT  1.005000 101.990000 15.870000 102.060000 ;
        RECT  1.005000 102.060000 15.940000 102.130000 ;
        RECT  1.005000 102.130000 16.010000 102.200000 ;
        RECT  1.005000 102.200000 16.080000 102.270000 ;
        RECT  1.005000 102.270000 16.150000 102.340000 ;
        RECT  1.005000 102.340000 16.220000 102.410000 ;
        RECT  1.005000 102.410000 16.290000 102.480000 ;
        RECT  1.005000 102.480000 16.360000 102.550000 ;
        RECT  1.005000 102.550000 16.430000 102.620000 ;
        RECT  1.005000 102.620000 16.500000 102.690000 ;
        RECT  1.005000 102.690000 16.570000 102.760000 ;
        RECT  1.005000 102.760000 16.640000 102.830000 ;
        RECT  1.005000 102.830000 16.710000 102.900000 ;
        RECT  1.005000 102.900000 16.780000 102.970000 ;
        RECT  1.005000 102.970000 16.850000 103.040000 ;
        RECT  1.005000 103.040000 16.920000 103.110000 ;
        RECT  1.005000 103.110000 16.990000 103.180000 ;
        RECT  1.005000 103.180000 17.060000 103.250000 ;
        RECT  1.005000 103.250000 17.130000 103.320000 ;
        RECT  1.005000 103.320000 17.200000 103.390000 ;
        RECT  1.005000 103.390000 17.270000 103.460000 ;
        RECT  1.005000 103.460000 17.340000 103.530000 ;
        RECT  1.005000 103.530000 17.410000 103.600000 ;
        RECT  1.005000 103.600000 17.480000 103.670000 ;
        RECT  1.005000 103.670000 17.550000 103.740000 ;
        RECT  1.005000 103.740000 17.620000 103.780000 ;
        RECT  1.005000 103.780000 56.705000 112.480000 ;
        RECT  1.005000 112.480000 17.635000 112.550000 ;
        RECT  1.005000 112.550000 17.565000 112.620000 ;
        RECT  1.005000 112.620000 17.495000 112.690000 ;
        RECT  1.005000 112.690000 17.425000 112.760000 ;
        RECT  1.005000 112.760000 17.355000 112.830000 ;
        RECT  1.005000 112.830000 17.285000 112.900000 ;
        RECT  1.005000 112.900000 17.215000 112.970000 ;
        RECT  1.005000 112.970000 17.145000 113.040000 ;
        RECT  1.005000 113.040000 17.075000 113.110000 ;
        RECT  1.005000 113.110000 17.005000 113.180000 ;
        RECT  1.005000 113.180000 16.935000 113.250000 ;
        RECT  1.005000 113.250000 16.865000 113.320000 ;
        RECT  1.005000 113.320000 16.795000 113.390000 ;
        RECT  1.005000 113.390000 16.725000 113.460000 ;
        RECT  1.005000 113.460000 16.655000 113.530000 ;
        RECT  1.005000 113.530000 16.585000 113.600000 ;
        RECT  1.005000 113.600000 16.515000 113.670000 ;
        RECT  1.005000 113.670000 16.445000 113.740000 ;
        RECT  1.005000 113.740000 16.375000 113.810000 ;
        RECT  1.005000 113.810000 16.305000 113.880000 ;
        RECT  1.005000 113.880000 16.235000 113.950000 ;
        RECT  1.005000 113.950000 16.165000 114.020000 ;
        RECT  1.005000 114.020000 16.095000 114.090000 ;
        RECT  1.005000 114.090000 16.025000 114.160000 ;
        RECT  1.005000 114.160000 15.955000 114.230000 ;
        RECT  1.005000 114.230000 15.885000 114.300000 ;
        RECT  1.005000 114.300000 15.815000 114.370000 ;
        RECT  1.005000 114.370000 15.745000 114.440000 ;
        RECT  1.005000 114.440000 15.675000 114.510000 ;
        RECT  1.005000 114.510000 15.605000 114.580000 ;
        RECT  1.005000 114.580000 15.535000 114.650000 ;
        RECT  1.005000 114.650000 15.465000 114.720000 ;
        RECT  1.005000 114.720000 15.395000 114.790000 ;
        RECT  1.005000 114.790000 15.325000 114.860000 ;
        RECT  1.005000 114.860000 15.255000 114.930000 ;
        RECT  1.005000 114.930000 15.185000 115.000000 ;
        RECT  1.005000 115.000000 15.115000 115.070000 ;
        RECT  1.005000 115.070000 15.045000 115.140000 ;
        RECT  1.005000 115.140000 14.975000 115.210000 ;
        RECT  1.005000 115.210000 14.905000 115.280000 ;
        RECT  1.005000 115.280000 14.835000 115.350000 ;
        RECT  1.005000 115.350000 14.765000 115.420000 ;
        RECT  1.005000 115.420000 14.695000 115.490000 ;
        RECT  1.005000 115.490000 14.625000 115.560000 ;
        RECT  1.005000 115.560000 14.555000 115.630000 ;
        RECT  1.005000 115.630000 14.485000 115.700000 ;
        RECT  1.005000 115.700000 14.415000 115.770000 ;
        RECT  1.005000 115.770000 14.345000 115.840000 ;
        RECT  1.005000 115.840000 14.275000 115.910000 ;
        RECT  1.005000 115.910000 14.205000 115.980000 ;
        RECT  1.005000 115.980000 14.135000 116.050000 ;
        RECT  1.005000 116.050000 14.120000 116.065000 ;
        RECT  1.005000 116.065000 14.120000 123.145000 ;
        RECT  1.005000 123.145000 14.120000 123.215000 ;
        RECT  1.005000 123.215000 14.190000 123.285000 ;
        RECT  1.005000 123.285000 14.260000 123.355000 ;
        RECT  1.005000 123.355000 14.330000 123.425000 ;
        RECT  1.005000 123.425000 14.400000 123.495000 ;
        RECT  1.005000 123.495000 14.470000 123.565000 ;
        RECT  1.005000 123.565000 14.540000 123.635000 ;
        RECT  1.005000 123.635000 14.610000 123.705000 ;
        RECT  1.005000 123.705000 14.680000 123.775000 ;
        RECT  1.005000 123.775000 14.750000 123.845000 ;
        RECT  1.005000 123.845000 14.820000 123.915000 ;
        RECT  1.005000 123.915000 14.890000 123.985000 ;
        RECT  1.005000 123.985000 14.960000 124.055000 ;
        RECT  1.005000 124.055000 15.030000 124.125000 ;
        RECT  1.005000 124.125000 15.100000 124.195000 ;
        RECT  1.005000 124.195000 15.170000 124.265000 ;
        RECT  1.005000 124.265000 15.240000 124.335000 ;
        RECT  1.005000 124.335000 15.310000 124.405000 ;
        RECT  1.005000 124.405000 15.380000 124.475000 ;
        RECT  1.005000 124.475000 15.450000 124.545000 ;
        RECT  1.005000 124.545000 15.520000 124.615000 ;
        RECT  1.005000 124.615000 15.590000 124.685000 ;
        RECT  1.005000 124.685000 15.660000 124.755000 ;
        RECT  1.005000 124.755000 15.730000 124.825000 ;
        RECT  1.005000 124.825000 15.800000 124.895000 ;
        RECT  1.005000 124.895000 15.870000 124.965000 ;
        RECT  1.005000 124.965000 15.940000 125.035000 ;
        RECT  1.005000 125.035000 16.010000 125.105000 ;
        RECT  1.005000 125.105000 16.080000 125.175000 ;
        RECT  1.005000 125.175000 16.150000 125.245000 ;
        RECT  1.005000 125.245000 16.220000 125.315000 ;
        RECT  1.005000 125.315000 16.290000 125.385000 ;
        RECT  1.005000 125.385000 16.360000 125.455000 ;
        RECT  1.005000 125.455000 16.430000 125.525000 ;
        RECT  1.005000 125.525000 16.500000 125.595000 ;
        RECT  1.005000 125.595000 16.570000 125.665000 ;
        RECT  1.005000 125.665000 16.640000 125.735000 ;
        RECT  1.005000 125.735000 16.710000 125.805000 ;
        RECT  1.005000 125.805000 16.780000 125.875000 ;
        RECT  1.005000 125.875000 16.850000 125.945000 ;
        RECT  1.005000 125.945000 16.920000 126.015000 ;
        RECT  1.005000 126.015000 16.990000 126.085000 ;
        RECT  1.005000 126.085000 17.060000 126.155000 ;
        RECT  1.005000 126.155000 17.130000 126.225000 ;
        RECT  1.005000 126.225000 17.200000 126.295000 ;
        RECT  1.005000 126.295000 17.270000 126.365000 ;
        RECT  1.005000 126.365000 17.340000 126.435000 ;
        RECT  1.005000 126.435000 17.410000 126.505000 ;
        RECT  1.005000 126.505000 17.480000 126.575000 ;
        RECT  1.005000 126.575000 17.550000 126.645000 ;
        RECT  1.005000 126.645000 17.620000 126.715000 ;
        RECT  1.005000 126.715000 17.690000 126.780000 ;
        RECT  1.005000 126.780000 56.705000 135.480000 ;
        RECT  1.005000 135.480000 17.740000 135.550000 ;
        RECT  1.005000 135.550000 17.670000 135.620000 ;
        RECT  1.005000 135.620000 17.600000 135.690000 ;
        RECT  1.005000 135.690000 17.530000 135.760000 ;
        RECT  1.005000 135.760000 17.460000 135.830000 ;
        RECT  1.005000 135.830000 17.390000 135.900000 ;
        RECT  1.005000 135.900000 17.320000 135.970000 ;
        RECT  1.005000 135.970000 17.250000 136.040000 ;
        RECT  1.005000 136.040000 17.180000 136.110000 ;
        RECT  1.005000 136.110000 17.110000 136.180000 ;
        RECT  1.005000 136.180000 17.040000 136.250000 ;
        RECT  1.005000 136.250000 16.970000 136.320000 ;
        RECT  1.005000 136.320000 16.900000 136.390000 ;
        RECT  1.005000 136.390000 16.830000 136.460000 ;
        RECT  1.005000 136.460000 16.760000 136.530000 ;
        RECT  1.005000 136.530000 16.690000 136.600000 ;
        RECT  1.005000 136.600000 16.620000 136.670000 ;
        RECT  1.005000 136.670000 16.550000 136.740000 ;
        RECT  1.005000 136.740000 16.480000 136.810000 ;
        RECT  1.005000 136.810000 16.410000 136.880000 ;
        RECT  1.005000 136.880000 16.340000 136.950000 ;
        RECT  1.005000 136.950000 16.270000 137.020000 ;
        RECT  1.005000 137.020000 16.200000 137.090000 ;
        RECT  1.005000 137.090000 16.130000 137.160000 ;
        RECT  1.005000 137.160000 16.060000 137.230000 ;
        RECT  1.005000 137.230000 15.990000 137.300000 ;
        RECT  1.005000 137.300000 15.920000 137.370000 ;
        RECT  1.005000 137.370000 15.850000 137.440000 ;
        RECT  1.005000 137.440000 15.780000 137.510000 ;
        RECT  1.005000 137.510000 15.710000 137.580000 ;
        RECT  1.005000 137.580000 15.640000 137.650000 ;
        RECT  1.005000 137.650000 15.570000 137.720000 ;
        RECT  1.005000 137.720000 15.500000 137.790000 ;
        RECT  1.005000 137.790000 15.430000 137.860000 ;
        RECT  1.005000 137.860000 15.360000 137.930000 ;
        RECT  1.005000 137.930000 15.290000 138.000000 ;
        RECT  1.005000 138.000000 15.220000 138.070000 ;
        RECT  1.005000 138.070000 15.150000 138.140000 ;
        RECT  1.005000 138.140000 15.080000 138.210000 ;
        RECT  1.005000 138.210000 15.010000 138.280000 ;
        RECT  1.005000 138.280000 14.940000 138.350000 ;
        RECT  1.005000 138.350000 14.870000 138.420000 ;
        RECT  1.005000 138.420000 14.800000 138.490000 ;
        RECT  1.005000 138.490000 14.730000 138.560000 ;
        RECT  1.005000 138.560000 14.660000 138.630000 ;
        RECT  1.005000 138.630000 14.590000 138.700000 ;
        RECT  1.005000 138.700000 14.520000 138.770000 ;
        RECT  1.005000 138.770000 14.450000 138.840000 ;
        RECT  1.005000 138.840000 14.380000 138.910000 ;
        RECT  1.005000 138.910000 14.310000 138.980000 ;
        RECT  1.005000 138.980000 14.240000 139.050000 ;
        RECT  1.005000 139.050000 14.170000 139.120000 ;
        RECT  1.005000 139.120000 14.120000 139.170000 ;
        RECT  1.005000 139.170000 14.120000 146.215000 ;
        RECT  1.005000 146.215000 14.120000 146.285000 ;
        RECT  1.005000 146.285000 14.190000 146.355000 ;
        RECT  1.005000 146.355000 14.260000 146.425000 ;
        RECT  1.005000 146.425000 14.330000 146.495000 ;
        RECT  1.005000 146.495000 14.400000 146.565000 ;
        RECT  1.005000 146.565000 14.470000 146.635000 ;
        RECT  1.005000 146.635000 14.540000 146.705000 ;
        RECT  1.005000 146.705000 14.610000 146.775000 ;
        RECT  1.005000 146.775000 14.680000 146.845000 ;
        RECT  1.005000 146.845000 14.750000 146.915000 ;
        RECT  1.005000 146.915000 14.820000 146.985000 ;
        RECT  1.005000 146.985000 14.890000 147.055000 ;
        RECT  1.005000 147.055000 14.960000 147.125000 ;
        RECT  1.005000 147.125000 15.030000 147.195000 ;
        RECT  1.005000 147.195000 15.100000 147.265000 ;
        RECT  1.005000 147.265000 15.170000 147.335000 ;
        RECT  1.005000 147.335000 15.240000 147.405000 ;
        RECT  1.005000 147.405000 15.310000 147.475000 ;
        RECT  1.005000 147.475000 15.380000 147.545000 ;
        RECT  1.005000 147.545000 15.450000 147.615000 ;
        RECT  1.005000 147.615000 15.520000 147.685000 ;
        RECT  1.005000 147.685000 15.590000 147.755000 ;
        RECT  1.005000 147.755000 15.660000 147.825000 ;
        RECT  1.005000 147.825000 15.730000 147.895000 ;
        RECT  1.005000 147.895000 15.800000 147.965000 ;
        RECT  1.005000 147.965000 15.870000 148.035000 ;
        RECT  1.005000 148.035000 15.940000 148.105000 ;
        RECT  1.005000 148.105000 16.010000 148.175000 ;
        RECT  1.005000 148.175000 16.080000 148.245000 ;
        RECT  1.005000 148.245000 16.150000 148.315000 ;
        RECT  1.005000 148.315000 16.220000 148.385000 ;
        RECT  1.005000 148.385000 16.290000 148.455000 ;
        RECT  1.005000 148.455000 16.360000 148.525000 ;
        RECT  1.005000 148.525000 16.430000 148.595000 ;
        RECT  1.005000 148.595000 16.500000 148.665000 ;
        RECT  1.005000 148.665000 16.570000 148.735000 ;
        RECT  1.005000 148.735000 16.640000 148.805000 ;
        RECT  1.005000 148.805000 16.710000 148.875000 ;
        RECT  1.005000 148.875000 16.780000 148.945000 ;
        RECT  1.005000 148.945000 16.850000 149.015000 ;
        RECT  1.005000 149.015000 16.920000 149.085000 ;
        RECT  1.005000 149.085000 16.990000 149.155000 ;
        RECT  1.005000 149.155000 17.060000 149.225000 ;
        RECT  1.005000 149.225000 17.130000 149.295000 ;
        RECT  1.005000 149.295000 17.200000 149.365000 ;
        RECT  1.005000 149.365000 17.270000 149.435000 ;
        RECT  1.005000 149.435000 17.340000 149.505000 ;
        RECT  1.005000 149.505000 17.410000 149.575000 ;
        RECT  1.005000 149.575000 17.480000 149.645000 ;
        RECT  1.005000 149.645000 17.550000 149.715000 ;
        RECT  1.005000 149.715000 17.620000 149.780000 ;
        RECT  1.005000 149.780000 56.705000 158.480000 ;
        RECT  1.005000 158.480000 17.650000 158.550000 ;
        RECT  1.005000 158.550000 17.580000 158.620000 ;
        RECT  1.005000 158.620000 17.510000 158.690000 ;
        RECT  1.005000 158.690000 17.440000 158.760000 ;
        RECT  1.005000 158.760000 17.370000 158.830000 ;
        RECT  1.005000 158.830000 17.300000 158.900000 ;
        RECT  1.005000 158.900000 17.230000 158.970000 ;
        RECT  1.005000 158.970000 17.160000 159.040000 ;
        RECT  1.005000 159.040000 17.090000 159.110000 ;
        RECT  1.005000 159.110000 17.020000 159.180000 ;
        RECT  1.005000 159.180000 16.950000 159.250000 ;
        RECT  1.005000 159.250000 16.880000 159.320000 ;
        RECT  1.005000 159.320000 16.810000 159.390000 ;
        RECT  1.005000 159.390000 16.740000 159.460000 ;
        RECT  1.005000 159.460000 16.670000 159.530000 ;
        RECT  1.005000 159.530000 16.600000 159.600000 ;
        RECT  1.005000 159.600000 16.530000 159.670000 ;
        RECT  1.005000 159.670000 16.460000 159.740000 ;
        RECT  1.005000 159.740000 16.390000 159.810000 ;
        RECT  1.005000 159.810000 16.320000 159.880000 ;
        RECT  1.005000 159.880000 16.250000 159.950000 ;
        RECT  1.005000 159.950000 16.180000 160.020000 ;
        RECT  1.005000 160.020000 16.110000 160.090000 ;
        RECT  1.005000 160.090000 16.040000 160.160000 ;
        RECT  1.005000 160.160000 15.970000 160.230000 ;
        RECT  1.005000 160.230000 15.900000 160.300000 ;
        RECT  1.005000 160.300000 15.830000 160.370000 ;
        RECT  1.005000 160.370000 15.760000 160.440000 ;
        RECT  1.005000 160.440000 15.690000 160.510000 ;
        RECT  1.005000 160.510000 15.620000 160.580000 ;
        RECT  1.005000 160.580000 15.550000 160.650000 ;
        RECT  1.005000 160.650000 15.480000 160.720000 ;
        RECT  1.005000 160.720000 15.410000 160.790000 ;
        RECT  1.005000 160.790000 15.340000 160.860000 ;
        RECT  1.005000 160.860000 15.270000 160.930000 ;
        RECT  1.005000 160.930000 15.200000 161.000000 ;
        RECT  1.005000 161.000000 15.130000 161.070000 ;
        RECT  1.005000 161.070000 15.060000 161.140000 ;
        RECT  1.005000 161.140000 14.990000 161.210000 ;
        RECT  1.005000 161.210000 14.920000 161.280000 ;
        RECT  1.005000 161.280000 14.850000 161.350000 ;
        RECT  1.005000 161.350000 14.780000 161.420000 ;
        RECT  1.005000 161.420000 14.710000 161.490000 ;
        RECT  1.005000 161.490000 14.640000 161.560000 ;
        RECT  1.005000 161.560000 14.570000 161.630000 ;
        RECT  1.005000 161.630000 14.500000 161.700000 ;
        RECT  1.005000 161.700000 14.430000 161.770000 ;
        RECT  1.005000 161.770000 14.360000 161.840000 ;
        RECT  1.005000 161.840000 14.290000 161.910000 ;
        RECT  1.005000 161.910000 14.220000 161.980000 ;
        RECT  1.005000 161.980000 14.150000 162.050000 ;
        RECT  1.005000 162.050000 14.120000 162.080000 ;
        RECT  1.005000 162.080000 14.120000 169.220000 ;
        RECT  1.005000 169.220000 14.120000 169.290000 ;
        RECT  1.005000 169.290000 14.190000 169.360000 ;
        RECT  1.005000 169.360000 14.260000 169.430000 ;
        RECT  1.005000 169.430000 14.330000 169.500000 ;
        RECT  1.005000 169.500000 14.400000 169.570000 ;
        RECT  1.005000 169.570000 14.470000 169.640000 ;
        RECT  1.005000 169.640000 14.540000 169.710000 ;
        RECT  1.005000 169.710000 14.610000 169.780000 ;
        RECT  1.005000 169.780000 14.680000 169.850000 ;
        RECT  1.005000 169.850000 14.750000 169.920000 ;
        RECT  1.005000 169.920000 14.820000 169.990000 ;
        RECT  1.005000 169.990000 14.890000 170.060000 ;
        RECT  1.005000 170.060000 14.960000 170.130000 ;
        RECT  1.005000 170.130000 15.030000 170.200000 ;
        RECT  1.005000 170.200000 15.100000 170.270000 ;
        RECT  1.005000 170.270000 15.170000 170.340000 ;
        RECT  1.005000 170.340000 15.240000 170.410000 ;
        RECT  1.005000 170.410000 15.310000 170.480000 ;
        RECT  1.005000 170.480000 15.380000 170.550000 ;
        RECT  1.005000 170.550000 15.450000 170.620000 ;
        RECT  1.005000 170.620000 15.520000 170.690000 ;
        RECT  1.005000 170.690000 15.590000 170.760000 ;
        RECT  1.005000 170.760000 15.660000 170.830000 ;
        RECT  1.005000 170.830000 15.730000 170.900000 ;
        RECT  1.005000 170.900000 15.800000 170.970000 ;
        RECT  1.005000 170.970000 15.870000 171.040000 ;
        RECT  1.005000 171.040000 15.940000 171.110000 ;
        RECT  1.005000 171.110000 16.010000 171.180000 ;
        RECT  1.005000 171.180000 16.080000 171.250000 ;
        RECT  1.005000 171.250000 16.150000 171.320000 ;
        RECT  1.005000 171.320000 16.220000 171.390000 ;
        RECT  1.005000 171.390000 16.290000 171.460000 ;
        RECT  1.005000 171.460000 16.360000 171.530000 ;
        RECT  1.005000 171.530000 16.430000 171.600000 ;
        RECT  1.005000 171.600000 16.500000 171.670000 ;
        RECT  1.005000 171.670000 16.570000 171.740000 ;
        RECT  1.005000 171.740000 16.640000 171.810000 ;
        RECT  1.005000 171.810000 16.710000 171.880000 ;
        RECT  1.005000 171.880000 16.780000 171.950000 ;
        RECT  1.005000 171.950000 16.850000 172.020000 ;
        RECT  1.005000 172.020000 16.920000 172.090000 ;
        RECT  1.005000 172.090000 16.990000 172.160000 ;
        RECT  1.005000 172.160000 17.060000 172.230000 ;
        RECT  1.005000 172.230000 17.130000 172.300000 ;
        RECT  1.005000 172.300000 17.200000 172.370000 ;
        RECT  1.005000 172.370000 17.270000 172.440000 ;
        RECT  1.005000 172.440000 17.340000 172.510000 ;
        RECT  1.005000 172.510000 17.410000 172.580000 ;
        RECT  1.005000 172.580000 17.480000 172.650000 ;
        RECT  1.005000 172.650000 17.550000 172.720000 ;
        RECT  1.005000 172.720000 17.620000 172.780000 ;
        RECT  1.005000 172.780000 57.960000 181.480000 ;
        RECT  1.005000 181.480000 17.625000 181.550000 ;
        RECT  1.005000 181.550000 17.555000 181.620000 ;
        RECT  1.005000 181.620000 17.485000 181.690000 ;
        RECT  1.005000 181.690000 17.415000 181.760000 ;
        RECT  1.005000 181.760000 17.345000 181.830000 ;
        RECT  1.005000 181.830000 17.275000 181.900000 ;
        RECT  1.005000 181.900000 17.205000 181.970000 ;
        RECT  1.005000 181.970000 17.135000 182.040000 ;
        RECT  1.005000 182.040000 17.065000 182.110000 ;
        RECT  1.005000 182.110000 16.995000 182.180000 ;
        RECT  1.005000 182.180000 16.925000 182.250000 ;
        RECT  1.005000 182.250000 16.855000 182.320000 ;
        RECT  1.005000 182.320000 16.785000 182.390000 ;
        RECT  1.005000 182.390000 16.715000 182.460000 ;
        RECT  1.005000 182.460000 16.645000 182.530000 ;
        RECT  1.005000 182.530000 16.575000 182.600000 ;
        RECT  1.005000 182.600000 16.505000 182.670000 ;
        RECT  1.005000 182.670000 16.435000 182.740000 ;
        RECT  1.005000 182.740000 16.365000 182.810000 ;
        RECT  1.005000 182.810000 16.295000 182.880000 ;
        RECT  1.005000 182.880000 16.225000 182.950000 ;
        RECT  1.005000 182.950000 16.155000 183.020000 ;
        RECT  1.005000 183.020000 16.085000 183.090000 ;
        RECT  1.005000 183.090000 16.015000 183.160000 ;
        RECT  1.005000 183.160000 15.945000 183.230000 ;
        RECT  1.005000 183.230000 15.875000 183.300000 ;
        RECT  1.005000 183.300000 15.805000 183.370000 ;
        RECT  1.005000 183.370000 15.735000 183.440000 ;
        RECT  1.005000 183.440000 15.665000 183.510000 ;
        RECT  1.005000 183.510000 15.595000 183.580000 ;
        RECT  1.005000 183.580000 15.525000 183.650000 ;
        RECT  1.005000 183.650000 15.455000 183.720000 ;
        RECT  1.005000 183.720000 15.385000 183.790000 ;
        RECT  1.005000 183.790000 15.315000 183.860000 ;
        RECT  1.005000 183.860000 15.245000 183.930000 ;
        RECT  1.005000 183.930000 15.175000 184.000000 ;
        RECT  1.005000 184.000000 15.105000 184.070000 ;
        RECT  1.005000 184.070000 15.035000 184.140000 ;
        RECT  1.005000 184.140000 14.965000 184.210000 ;
        RECT  1.005000 184.210000 14.895000 184.280000 ;
        RECT  1.005000 184.280000 14.825000 184.350000 ;
        RECT  1.005000 184.350000 14.755000 184.420000 ;
        RECT  1.005000 184.420000 14.685000 184.490000 ;
        RECT  1.005000 184.490000 14.615000 184.560000 ;
        RECT  1.005000 184.560000 14.545000 184.630000 ;
        RECT  1.005000 184.630000 14.475000 184.700000 ;
        RECT  1.005000 184.700000 14.405000 184.770000 ;
        RECT  1.005000 184.770000 14.335000 184.840000 ;
        RECT  1.005000 184.840000 14.265000 184.910000 ;
        RECT  1.005000 184.910000 14.195000 184.980000 ;
        RECT  1.005000 184.980000 14.125000 185.050000 ;
        RECT  1.005000 185.050000 14.120000 185.055000 ;
        RECT  1.005000 185.055000 14.120000 189.585000 ;
        RECT  1.005000 189.585000 14.120000 189.655000 ;
        RECT  1.005000 189.655000 14.190000 189.725000 ;
        RECT  1.005000 189.725000 14.260000 189.795000 ;
        RECT  1.005000 189.795000 14.330000 189.865000 ;
        RECT  1.005000 189.865000 14.400000 189.935000 ;
        RECT  1.005000 189.935000 14.470000 190.005000 ;
        RECT  1.005000 190.005000 14.540000 190.075000 ;
        RECT  1.005000 190.075000 14.610000 190.145000 ;
        RECT  1.005000 190.145000 14.680000 190.215000 ;
        RECT  1.005000 190.215000 14.750000 190.285000 ;
        RECT  1.005000 190.285000 14.820000 190.355000 ;
        RECT  1.005000 190.355000 14.890000 190.425000 ;
        RECT  1.005000 190.425000 14.960000 190.495000 ;
        RECT  1.005000 190.495000 15.030000 190.560000 ;
        RECT  1.005000 190.560000 67.200000 195.075000 ;
        RECT  1.010000  47.125000 14.120000  47.130000 ;
        RECT  1.045000  36.640000 16.180000  36.680000 ;
        RECT  1.050000  47.085000 14.120000  47.125000 ;
        RECT  1.085000  36.680000 16.220000  36.720000 ;
        RECT  1.090000  36.720000 16.260000  36.725000 ;
        RECT  1.090000  36.725000 16.265000  36.795000 ;
        RECT  1.090000  36.795000 16.335000  36.865000 ;
        RECT  1.090000  36.865000 16.405000  36.935000 ;
        RECT  1.090000  36.935000 16.475000  37.005000 ;
        RECT  1.090000  37.005000 16.545000  37.075000 ;
        RECT  1.090000  37.075000 16.615000  37.145000 ;
        RECT  1.090000  37.145000 16.685000  37.215000 ;
        RECT  1.090000  37.215000 16.755000  37.285000 ;
        RECT  1.090000  37.285000 16.825000  37.355000 ;
        RECT  1.090000  37.355000 16.895000  37.425000 ;
        RECT  1.090000  37.425000 16.965000  37.495000 ;
        RECT  1.090000  37.495000 17.035000  37.565000 ;
        RECT  1.090000  37.565000 17.105000  37.635000 ;
        RECT  1.090000  37.635000 17.175000  37.705000 ;
        RECT  1.090000  37.705000 17.245000  37.775000 ;
        RECT  1.090000  37.775000 17.315000  37.845000 ;
        RECT  1.090000  37.845000 17.385000  37.915000 ;
        RECT  1.090000  37.915000 17.455000  37.985000 ;
        RECT  1.090000  37.985000 17.525000  38.055000 ;
        RECT  1.090000  38.055000 17.595000  38.125000 ;
        RECT  1.090000  38.125000 17.665000  38.195000 ;
        RECT  1.090000  38.195000 17.735000  38.265000 ;
        RECT  1.090000  38.265000 17.805000  38.335000 ;
        RECT  1.090000  38.335000 17.875000  38.405000 ;
        RECT  1.090000  38.405000 17.945000  38.475000 ;
        RECT  1.090000  38.475000 18.015000  38.545000 ;
        RECT  1.090000  38.545000 18.085000  38.615000 ;
        RECT  1.090000  38.615000 18.155000  38.685000 ;
        RECT  1.090000  38.685000 18.225000  38.755000 ;
        RECT  1.090000  38.755000 18.295000  38.825000 ;
        RECT  1.090000  38.825000 18.365000  38.895000 ;
        RECT  1.090000  38.895000 18.435000  38.965000 ;
        RECT  1.090000  38.965000 18.505000  39.035000 ;
        RECT  1.090000  39.035000 18.575000  39.105000 ;
        RECT  1.090000  39.105000 18.645000  39.175000 ;
        RECT  1.090000  39.175000 18.715000  39.245000 ;
        RECT  1.090000  39.245000 18.785000  39.315000 ;
        RECT  1.090000  39.315000 18.855000  39.385000 ;
        RECT  1.090000  39.385000 18.925000  39.455000 ;
        RECT  1.090000  39.455000 18.995000  39.525000 ;
        RECT  1.090000  39.525000 19.065000  39.595000 ;
        RECT  1.090000  39.595000 19.135000  39.665000 ;
        RECT  1.090000  39.665000 19.205000  39.735000 ;
        RECT  1.090000  39.735000 19.275000  39.805000 ;
        RECT  1.090000  39.805000 19.345000  39.875000 ;
        RECT  1.090000  39.875000 19.415000  39.945000 ;
        RECT  1.090000  39.945000 19.485000  40.015000 ;
        RECT  1.090000  40.015000 19.555000  40.085000 ;
        RECT  1.090000  40.085000 19.625000  40.155000 ;
        RECT  1.090000  40.155000 19.695000  40.225000 ;
        RECT  1.090000  40.225000 19.765000  40.295000 ;
        RECT  1.090000  40.295000 19.835000  40.350000 ;
        RECT  1.090000  40.350000 56.160000  40.420000 ;
        RECT  1.090000  40.420000 56.090000  40.490000 ;
        RECT  1.090000  40.490000 56.020000  40.560000 ;
        RECT  1.090000  40.560000 55.950000  40.630000 ;
        RECT  1.090000  40.630000 55.880000  40.700000 ;
        RECT  1.090000  40.700000 55.810000  40.770000 ;
        RECT  1.090000  40.770000 55.740000  40.840000 ;
        RECT  1.090000  40.840000 55.670000  40.910000 ;
        RECT  1.090000  40.910000 55.600000  40.980000 ;
        RECT  1.090000  40.980000 55.530000  41.050000 ;
        RECT  1.090000  41.050000 55.460000  41.120000 ;
        RECT  1.090000  41.120000 55.390000  41.190000 ;
        RECT  1.090000  41.190000 55.320000  41.260000 ;
        RECT  1.090000  41.260000 55.250000  41.330000 ;
        RECT  1.090000  41.330000 55.180000  41.400000 ;
        RECT  1.090000  41.400000 55.110000  41.470000 ;
        RECT  1.090000  41.470000 55.040000  41.540000 ;
        RECT  1.090000  41.540000 54.970000  41.610000 ;
        RECT  1.090000  41.610000 54.900000  41.680000 ;
        RECT  1.090000  41.680000 54.830000  41.750000 ;
        RECT  1.090000  41.750000 54.760000  41.820000 ;
        RECT  1.090000  41.820000 54.690000  41.890000 ;
        RECT  1.090000  41.890000 54.620000  41.960000 ;
        RECT  1.090000  41.960000 54.550000  42.030000 ;
        RECT  1.090000  42.030000 54.480000  42.100000 ;
        RECT  1.090000  42.100000 54.410000  42.170000 ;
        RECT  1.090000  42.170000 54.340000  42.240000 ;
        RECT  1.090000  42.240000 54.270000  42.310000 ;
        RECT  1.090000  42.310000 54.200000  42.380000 ;
        RECT  1.090000  42.380000 16.985000  42.450000 ;
        RECT  1.090000  42.450000 16.915000  42.520000 ;
        RECT  1.090000  42.520000 16.845000  42.590000 ;
        RECT  1.090000  42.590000 16.775000  42.660000 ;
        RECT  1.090000  42.660000 16.705000  42.730000 ;
        RECT  1.090000  42.730000 16.635000  42.800000 ;
        RECT  1.090000  42.800000 16.565000  42.870000 ;
        RECT  1.090000  42.870000 16.495000  42.940000 ;
        RECT  1.090000  42.940000 16.425000  43.010000 ;
        RECT  1.090000  43.010000 16.355000  43.080000 ;
        RECT  1.090000  43.080000 16.285000  43.150000 ;
        RECT  1.090000  43.150000 16.215000  43.220000 ;
        RECT  1.090000  43.220000 16.145000  43.290000 ;
        RECT  1.090000  43.290000 16.075000  43.360000 ;
        RECT  1.090000  43.360000 16.005000  43.430000 ;
        RECT  1.090000  43.430000 15.935000  43.500000 ;
        RECT  1.090000  43.500000 15.865000  43.570000 ;
        RECT  1.090000  43.570000 15.795000  43.640000 ;
        RECT  1.090000  43.640000 15.725000  43.710000 ;
        RECT  1.090000  43.710000 15.655000  43.780000 ;
        RECT  1.090000  43.780000 15.585000  43.850000 ;
        RECT  1.090000  43.850000 15.515000  43.920000 ;
        RECT  1.090000  43.920000 15.445000  43.990000 ;
        RECT  1.090000  43.990000 15.375000  44.060000 ;
        RECT  1.090000  44.060000 15.305000  44.130000 ;
        RECT  1.090000  44.130000 15.235000  44.200000 ;
        RECT  1.090000  44.200000 15.165000  44.270000 ;
        RECT  1.090000  44.270000 15.095000  44.340000 ;
        RECT  1.090000  44.340000 15.025000  44.410000 ;
        RECT  1.090000  44.410000 14.955000  44.480000 ;
        RECT  1.090000  44.480000 14.885000  44.550000 ;
        RECT  1.090000  44.550000 14.815000  44.620000 ;
        RECT  1.090000  44.620000 14.745000  44.690000 ;
        RECT  1.090000  44.690000 14.675000  44.760000 ;
        RECT  1.090000  44.760000 14.605000  44.830000 ;
        RECT  1.090000  44.830000 14.535000  44.900000 ;
        RECT  1.090000  44.900000 14.465000  44.970000 ;
        RECT  1.090000  44.970000 14.395000  45.040000 ;
        RECT  1.090000  45.040000 14.325000  45.110000 ;
        RECT  1.090000  45.110000 14.255000  45.180000 ;
        RECT  1.090000  45.180000 14.185000  45.250000 ;
        RECT  1.090000  45.250000 14.120000  45.315000 ;
        RECT  1.090000  45.315000 14.120000  47.045000 ;
        RECT  1.090000  47.045000 14.120000  47.085000 ;
        RECT 52.630000  40.295000 56.230000  40.350000 ;
        RECT 52.700000  40.225000 56.285000  40.295000 ;
        RECT 52.770000  40.155000 56.355000  40.225000 ;
        RECT 52.840000  40.085000 56.425000  40.155000 ;
        RECT 52.910000  40.015000 56.495000  40.085000 ;
        RECT 52.980000  39.945000 56.565000  40.015000 ;
        RECT 53.050000  39.875000 56.635000  39.945000 ;
        RECT 53.120000  39.805000 56.705000  39.875000 ;
        RECT 53.190000  39.735000 56.775000  39.805000 ;
        RECT 53.260000  39.665000 56.845000  39.735000 ;
        RECT 53.270000  39.655000 56.915000  39.665000 ;
        RECT 53.340000  39.585000 56.915000  39.655000 ;
        RECT 53.410000  39.515000 56.915000  39.585000 ;
        RECT 53.480000  39.445000 56.915000  39.515000 ;
        RECT 53.550000  39.375000 56.915000  39.445000 ;
        RECT 53.620000  39.305000 56.915000  39.375000 ;
        RECT 53.690000  39.235000 56.915000  39.305000 ;
        RECT 53.760000  39.165000 56.915000  39.235000 ;
        RECT 53.830000  39.095000 56.915000  39.165000 ;
        RECT 53.900000  39.025000 56.915000  39.095000 ;
        RECT 53.970000  38.955000 56.915000  39.025000 ;
        RECT 54.040000  38.885000 56.915000  38.955000 ;
        RECT 54.110000  38.815000 56.915000  38.885000 ;
        RECT 54.180000  38.745000 56.915000  38.815000 ;
        RECT 54.250000  38.675000 56.915000  38.745000 ;
        RECT 54.320000  38.605000 56.915000  38.675000 ;
        RECT 54.390000  38.535000 56.915000  38.605000 ;
        RECT 54.460000  38.465000 56.915000  38.535000 ;
        RECT 54.530000  38.395000 56.915000  38.465000 ;
        RECT 54.600000  38.325000 56.915000  38.395000 ;
        RECT 54.670000  36.115000 56.915000  38.255000 ;
        RECT 54.670000  38.255000 56.915000  38.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.050000 172.755000 25.010000 195.100000 ;
        RECT 14.055000 172.750000 25.010000 172.755000 ;
        RECT 14.110000 172.695000 25.010000 172.750000 ;
        RECT 14.165000 172.640000 25.010000 172.695000 ;
        RECT 14.300000 172.505000 24.875000 172.640000 ;
        RECT 14.450000 172.355000 24.725000 172.505000 ;
        RECT 14.600000 172.205000 24.575000 172.355000 ;
        RECT 14.750000 172.055000 24.425000 172.205000 ;
        RECT 14.900000 171.905000 24.275000 172.055000 ;
        RECT 15.050000 171.755000 24.125000 171.905000 ;
        RECT 15.200000 171.605000 23.975000 171.755000 ;
        RECT 15.350000 171.455000 23.825000 171.605000 ;
        RECT 15.500000 102.200000 23.830000 102.350000 ;
        RECT 15.500000 102.350000 23.680000 102.500000 ;
        RECT 15.500000 102.500000 23.530000 102.650000 ;
        RECT 15.500000 102.650000 23.380000 102.800000 ;
        RECT 15.500000 102.800000 23.230000 102.950000 ;
        RECT 15.500000 102.950000 23.080000 103.100000 ;
        RECT 15.500000 103.100000 22.930000 103.250000 ;
        RECT 15.500000 103.250000 22.780000 103.400000 ;
        RECT 15.500000 103.400000 22.630000 103.550000 ;
        RECT 15.500000 103.550000 22.480000 103.700000 ;
        RECT 15.500000 103.700000 22.330000 103.850000 ;
        RECT 15.500000 103.850000 22.180000 104.000000 ;
        RECT 15.500000 104.000000 22.030000 104.150000 ;
        RECT 15.500000 104.150000 21.880000 104.300000 ;
        RECT 15.500000 104.300000 21.730000 104.450000 ;
        RECT 15.500000 104.450000 21.580000 104.600000 ;
        RECT 15.500000 104.600000 21.500000 104.680000 ;
        RECT 15.500000 104.680000 21.500000 169.130000 ;
        RECT 15.500000 169.130000 21.500000 169.280000 ;
        RECT 15.500000 169.280000 21.650000 169.430000 ;
        RECT 15.500000 169.430000 21.800000 169.580000 ;
        RECT 15.500000 169.580000 21.950000 169.730000 ;
        RECT 15.500000 169.730000 22.100000 169.880000 ;
        RECT 15.500000 169.880000 22.250000 170.030000 ;
        RECT 15.500000 170.030000 22.400000 170.180000 ;
        RECT 15.500000 170.180000 22.550000 170.330000 ;
        RECT 15.500000 170.330000 22.700000 170.480000 ;
        RECT 15.500000 170.480000 22.850000 170.630000 ;
        RECT 15.500000 170.630000 23.000000 170.780000 ;
        RECT 15.500000 170.780000 23.150000 170.930000 ;
        RECT 15.500000 170.930000 23.300000 171.080000 ;
        RECT 15.500000 171.080000 23.450000 171.230000 ;
        RECT 15.500000 171.230000 23.600000 171.305000 ;
        RECT 15.500000 171.305000 23.675000 171.455000 ;
        RECT 15.645000 102.055000 23.980000 102.200000 ;
        RECT 15.795000 101.905000 24.125000 102.055000 ;
        RECT 15.945000 101.755000 24.275000 101.905000 ;
        RECT 16.095000 101.605000 24.425000 101.755000 ;
        RECT 16.245000 101.455000 24.575000 101.605000 ;
        RECT 16.395000 101.305000 24.725000 101.455000 ;
        RECT 16.545000 101.155000 24.875000 101.305000 ;
        RECT 16.695000 101.005000 25.025000 101.155000 ;
        RECT 16.845000 100.855000 25.175000 101.005000 ;
        RECT 16.995000 100.705000 25.325000 100.855000 ;
        RECT 17.145000 100.555000 25.475000 100.705000 ;
        RECT 17.295000 100.405000 25.625000 100.555000 ;
        RECT 17.445000 100.255000 25.775000 100.405000 ;
        RECT 17.595000 100.105000 25.925000 100.255000 ;
        RECT 17.745000  99.955000 26.075000 100.105000 ;
        RECT 17.895000  99.805000 26.225000  99.955000 ;
        RECT 18.045000  99.655000 26.375000  99.805000 ;
        RECT 18.195000  99.505000 26.525000  99.655000 ;
        RECT 18.345000  99.355000 26.675000  99.505000 ;
        RECT 18.495000  99.205000 26.825000  99.355000 ;
        RECT 18.645000  99.055000 26.975000  99.205000 ;
        RECT 18.795000  98.905000 27.125000  99.055000 ;
        RECT 18.945000  98.755000 27.275000  98.905000 ;
        RECT 19.095000  98.605000 27.425000  98.755000 ;
        RECT 19.245000  98.455000 27.575000  98.605000 ;
        RECT 19.395000  98.305000 27.725000  98.455000 ;
        RECT 19.545000  98.155000 27.875000  98.305000 ;
        RECT 19.695000  98.005000 28.025000  98.155000 ;
        RECT 19.845000  97.855000 28.175000  98.005000 ;
        RECT 19.995000  97.705000 28.325000  97.855000 ;
        RECT 20.145000  97.555000 28.475000  97.705000 ;
        RECT 20.295000  97.405000 28.625000  97.555000 ;
        RECT 20.445000  97.255000 28.775000  97.405000 ;
        RECT 20.595000  97.105000 28.925000  97.255000 ;
        RECT 20.745000  96.955000 29.075000  97.105000 ;
        RECT 20.895000  96.805000 29.225000  96.955000 ;
        RECT 21.045000  96.655000 29.375000  96.805000 ;
        RECT 21.195000  96.505000 29.525000  96.655000 ;
        RECT 21.345000  96.355000 29.525000  96.505000 ;
        RECT 21.495000  96.205000 29.525000  96.355000 ;
        RECT 21.645000  96.055000 29.525000  96.205000 ;
        RECT 21.795000  95.905000 29.525000  96.055000 ;
        RECT 21.945000  95.755000 29.525000  95.905000 ;
        RECT 22.095000  95.605000 29.525000  95.755000 ;
        RECT 22.245000  95.455000 29.525000  95.605000 ;
        RECT 22.395000  95.305000 29.525000  95.455000 ;
        RECT 22.545000  95.155000 29.525000  95.305000 ;
        RECT 22.695000  95.005000 29.525000  95.155000 ;
        RECT 22.845000  94.855000 29.525000  95.005000 ;
        RECT 22.995000  94.705000 29.525000  94.855000 ;
        RECT 23.145000  94.555000 29.525000  94.705000 ;
        RECT 23.295000  94.405000 29.525000  94.555000 ;
        RECT 23.445000  94.255000 29.525000  94.405000 ;
        RECT 23.595000  94.105000 29.525000  94.255000 ;
        RECT 23.745000  92.540000 29.935000  92.690000 ;
        RECT 23.745000  92.690000 29.785000  92.840000 ;
        RECT 23.745000  92.840000 29.635000  92.990000 ;
        RECT 23.745000  92.990000 29.525000  93.100000 ;
        RECT 23.745000  93.100000 29.525000  93.955000 ;
        RECT 23.745000  93.955000 29.525000  94.105000 ;
        RECT 23.820000  92.465000 30.085000  92.540000 ;
        RECT 23.895000  92.390000 30.160000  92.465000 ;
        RECT 23.945000  92.340000 36.895000  92.390000 ;
        RECT 24.095000  92.190000 36.895000  92.340000 ;
        RECT 24.245000  92.040000 36.895000  92.190000 ;
        RECT 24.395000  91.890000 36.895000  92.040000 ;
        RECT 24.545000  91.740000 36.895000  91.890000 ;
        RECT 24.695000  91.590000 36.895000  91.740000 ;
        RECT 24.845000  91.440000 36.895000  91.590000 ;
        RECT 24.995000  91.290000 36.895000  91.440000 ;
        RECT 25.145000  91.140000 36.895000  91.290000 ;
        RECT 25.295000  90.990000 36.895000  91.140000 ;
        RECT 25.445000  90.840000 36.895000  90.990000 ;
        RECT 25.595000  90.690000 36.895000  90.840000 ;
        RECT 25.745000  90.540000 36.895000  90.690000 ;
        RECT 25.895000   0.000000 36.895000  90.390000 ;
        RECT 25.895000  90.390000 36.895000  90.540000 ;
        RECT 25.930000 102.390000 34.250000 102.540000 ;
        RECT 25.930000 102.540000 34.100000 102.690000 ;
        RECT 25.930000 102.690000 33.950000 102.840000 ;
        RECT 25.930000 102.840000 33.800000 102.990000 ;
        RECT 25.930000 102.990000 33.650000 103.140000 ;
        RECT 25.930000 103.140000 33.500000 103.290000 ;
        RECT 25.930000 103.290000 33.350000 103.440000 ;
        RECT 25.930000 103.440000 33.200000 103.590000 ;
        RECT 25.930000 103.590000 33.050000 103.740000 ;
        RECT 25.930000 103.740000 32.900000 103.890000 ;
        RECT 25.930000 103.890000 32.750000 104.040000 ;
        RECT 25.930000 104.040000 32.600000 104.190000 ;
        RECT 25.930000 104.190000 32.450000 104.340000 ;
        RECT 25.930000 104.340000 32.300000 104.490000 ;
        RECT 25.930000 104.490000 32.150000 104.640000 ;
        RECT 25.930000 104.640000 32.000000 104.790000 ;
        RECT 25.930000 104.790000 31.930000 104.860000 ;
        RECT 25.930000 104.860000 31.930000 170.460000 ;
        RECT 25.930000 170.460000 31.930000 170.610000 ;
        RECT 25.930000 170.610000 32.080000 170.760000 ;
        RECT 25.930000 170.760000 32.230000 170.910000 ;
        RECT 25.930000 170.910000 32.380000 171.060000 ;
        RECT 25.930000 171.060000 32.530000 171.210000 ;
        RECT 25.930000 171.210000 32.680000 171.360000 ;
        RECT 25.930000 171.360000 32.830000 171.510000 ;
        RECT 25.930000 171.510000 32.980000 171.660000 ;
        RECT 25.930000 171.660000 33.130000 171.810000 ;
        RECT 25.930000 171.810000 33.280000 171.960000 ;
        RECT 25.930000 171.960000 33.430000 172.110000 ;
        RECT 25.930000 172.110000 33.580000 172.260000 ;
        RECT 25.930000 172.260000 33.730000 172.410000 ;
        RECT 25.930000 172.410000 33.880000 172.560000 ;
        RECT 25.930000 172.560000 34.030000 172.710000 ;
        RECT 25.930000 172.710000 34.180000 172.860000 ;
        RECT 25.930000 172.860000 34.330000 173.010000 ;
        RECT 25.930000 173.010000 34.480000 173.160000 ;
        RECT 25.930000 173.160000 34.630000 173.310000 ;
        RECT 25.930000 173.310000 34.780000 173.460000 ;
        RECT 25.930000 173.460000 34.930000 173.610000 ;
        RECT 25.930000 173.610000 35.080000 173.760000 ;
        RECT 25.930000 173.760000 35.230000 173.910000 ;
        RECT 25.930000 173.910000 35.380000 174.060000 ;
        RECT 25.930000 174.060000 35.530000 174.210000 ;
        RECT 25.930000 174.210000 35.680000 174.360000 ;
        RECT 25.930000 174.360000 35.830000 174.510000 ;
        RECT 25.930000 174.510000 35.980000 174.660000 ;
        RECT 25.930000 174.660000 36.130000 174.810000 ;
        RECT 25.930000 174.810000 36.280000 174.960000 ;
        RECT 25.930000 174.960000 36.430000 175.110000 ;
        RECT 25.930000 175.110000 36.580000 175.260000 ;
        RECT 25.930000 175.260000 36.730000 175.350000 ;
        RECT 25.930000 175.350000 36.820000 195.100000 ;
        RECT 26.025000 102.295000 34.400000 102.390000 ;
        RECT 26.175000 102.145000 34.495000 102.295000 ;
        RECT 26.325000 101.995000 34.645000 102.145000 ;
        RECT 26.475000 101.845000 34.795000 101.995000 ;
        RECT 26.625000 101.695000 34.945000 101.845000 ;
        RECT 26.775000 101.545000 35.095000 101.695000 ;
        RECT 26.925000 101.395000 35.245000 101.545000 ;
        RECT 27.075000 101.245000 35.395000 101.395000 ;
        RECT 27.225000 101.095000 35.545000 101.245000 ;
        RECT 27.375000 100.945000 35.695000 101.095000 ;
        RECT 27.525000 100.795000 35.845000 100.945000 ;
        RECT 27.675000 100.645000 35.995000 100.795000 ;
        RECT 27.825000 100.495000 36.145000 100.645000 ;
        RECT 27.975000 100.345000 36.295000 100.495000 ;
        RECT 28.125000 100.195000 36.445000 100.345000 ;
        RECT 28.275000 100.045000 36.595000 100.195000 ;
        RECT 28.425000  99.895000 36.745000 100.045000 ;
        RECT 28.495000  99.825000 36.895000  99.895000 ;
        RECT 28.645000  99.675000 36.895000  99.825000 ;
        RECT 28.795000  99.525000 36.895000  99.675000 ;
        RECT 28.945000  99.375000 36.895000  99.525000 ;
        RECT 29.095000  99.225000 36.895000  99.375000 ;
        RECT 29.245000  99.075000 36.895000  99.225000 ;
        RECT 29.395000  98.925000 36.895000  99.075000 ;
        RECT 29.545000  98.775000 36.895000  98.925000 ;
        RECT 29.695000  98.625000 36.895000  98.775000 ;
        RECT 29.845000  98.475000 36.895000  98.625000 ;
        RECT 29.995000  98.325000 36.895000  98.475000 ;
        RECT 30.145000  98.175000 36.895000  98.325000 ;
        RECT 30.295000  98.025000 36.895000  98.175000 ;
        RECT 30.445000  97.875000 36.895000  98.025000 ;
        RECT 30.595000  97.725000 36.895000  97.875000 ;
        RECT 30.745000  97.575000 36.895000  97.725000 ;
        RECT 30.895000  97.425000 36.895000  97.575000 ;
        RECT 31.045000  97.275000 36.895000  97.425000 ;
        RECT 31.195000  97.125000 36.895000  97.275000 ;
        RECT 31.345000  96.975000 36.895000  97.125000 ;
        RECT 31.385000  92.390000 36.895000  92.540000 ;
        RECT 31.495000  96.825000 36.895000  96.975000 ;
        RECT 31.535000  92.540000 36.895000  92.690000 ;
        RECT 31.645000  96.675000 36.895000  96.825000 ;
        RECT 31.685000  92.690000 36.895000  92.840000 ;
        RECT 31.795000  96.525000 36.895000  96.675000 ;
        RECT 31.835000  92.840000 36.895000  92.990000 ;
        RECT 31.945000  92.990000 36.895000  93.100000 ;
        RECT 31.945000  93.100000 36.895000  96.375000 ;
        RECT 31.945000  96.375000 36.895000  96.525000 ;
    END
  END SRC_BDY_HVC
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  1.145000  43.280000  1.315000  43.810000 ;
      RECT  3.100000  27.160000 48.200000  28.030000 ;
      RECT  3.100000  28.030000  4.020000  38.695000 ;
      RECT  3.100000  38.695000 48.200000  39.565000 ;
      RECT  3.130000  27.140000 48.200000  27.160000 ;
      RECT  3.130000  39.565000 48.200000  39.585000 ;
      RECT  4.735000  29.230000 45.955000  29.430000 ;
      RECT  4.735000  29.430000  4.905000  37.425000 ;
      RECT  4.735000  37.425000 45.955000  37.595000 ;
      RECT  6.115000  33.340000  6.285000  36.490000 ;
      RECT  6.340000  36.970000 45.060000  37.230000 ;
      RECT  6.895000  29.775000  7.065000  32.860000 ;
      RECT  7.675000  33.335000  7.845000  36.490000 ;
      RECT  8.050000  43.270000  8.580000  43.440000 ;
      RECT  8.455000  29.770000  8.625000  32.860000 ;
      RECT  8.510000 162.655000 10.360000 169.150000 ;
      RECT  9.135000  43.505000 70.125000  44.755000 ;
      RECT  9.135000  44.755000 10.385000  71.570000 ;
      RECT  9.135000  71.570000 21.085000  72.820000 ;
      RECT  9.150000 169.400000 10.400000 198.445000 ;
      RECT  9.150000 198.445000 70.125000 199.695000 ;
      RECT  9.170000 133.350000 20.990000 134.540000 ;
      RECT  9.170000 134.540000 10.360000 162.655000 ;
      RECT  9.170000 169.150000 10.360000 169.400000 ;
      RECT  9.200000 133.205000 14.190000 133.350000 ;
      RECT  9.235000  33.340000  9.405000  36.490000 ;
      RECT  9.405000  74.180000  9.935000  74.350000 ;
      RECT 10.015000  29.775000 10.185000  32.860000 ;
      RECT 10.770000 162.655000 11.975000 169.905000 ;
      RECT 10.795000  33.335000 10.965000  36.490000 ;
      RECT 11.100000 170.415000 11.990000 196.835000 ;
      RECT 11.100000 196.835000 68.155000 197.725000 ;
      RECT 11.105000  45.460000 68.155000  46.350000 ;
      RECT 11.105000  46.350000 11.995000  69.975000 ;
      RECT 11.105000  69.975000 22.680000  70.865000 ;
      RECT 11.125000 135.315000 22.660000 136.165000 ;
      RECT 11.125000 136.165000 12.100000 158.915000 ;
      RECT 11.125000 158.915000 11.975000 162.655000 ;
      RECT 11.125000 169.905000 11.975000 170.415000 ;
      RECT 11.575000  29.770000 11.745000  32.860000 ;
      RECT 12.065000   1.000000 70.650000   1.890000 ;
      RECT 12.065000   1.890000 13.045000  22.230000 ;
      RECT 12.065000  22.230000 56.085000  22.350000 ;
      RECT 12.065000  22.350000 56.105000  23.240000 ;
      RECT 12.355000  33.340000 12.525000  36.490000 ;
      RECT 12.400000 159.555000 64.500000 161.990000 ;
      RECT 12.830000 182.570000 66.685000 184.990000 ;
      RECT 13.085000  46.815000 64.500000  46.990000 ;
      RECT 13.085000  46.990000 13.255000  67.965000 ;
      RECT 13.090000  46.740000 64.500000  46.815000 ;
      RECT 13.135000  29.775000 13.305000  32.860000 ;
      RECT 13.915000  33.335000 14.085000  36.490000 ;
      RECT 14.385000  47.160000 15.415000  66.930000 ;
      RECT 14.385000 139.160000 15.415000 158.930000 ;
      RECT 14.385000 162.160000 15.415000 181.930000 ;
      RECT 14.385000 185.160000 15.435000 195.185000 ;
      RECT 14.695000  29.770000 14.865000  32.860000 ;
      RECT 15.475000  33.340000 15.645000  36.490000 ;
      RECT 15.705000  67.340000 64.500000  68.995000 ;
      RECT 15.780000 136.540000 64.500000 138.990000 ;
      RECT 15.780000 159.340000 64.500000 159.555000 ;
      RECT 15.780000 182.340000 66.685000 182.570000 ;
      RECT 15.780000 195.370000 16.490000 195.540000 ;
      RECT 16.255000  29.770000 16.425000  32.860000 ;
      RECT 17.035000  33.335000 17.205000  36.490000 ;
      RECT 17.790000 195.370000 18.500000 195.540000 ;
      RECT 17.815000  29.770000 17.985000  32.860000 ;
      RECT 17.835000 133.145000 20.990000 133.350000 ;
      RECT 18.470000  74.200000 19.000000  74.370000 ;
      RECT 18.595000  33.340000 18.765000  36.490000 ;
      RECT 18.985000  47.515000 19.875000  66.855000 ;
      RECT 18.985000 139.515000 19.875000 158.810000 ;
      RECT 18.985000 162.515000 19.875000 181.810000 ;
      RECT 18.985000 185.515000 19.875000 195.075000 ;
      RECT 19.375000  29.775000 19.545000  32.860000 ;
      RECT 19.565000  97.500000 20.990000 133.145000 ;
      RECT 19.800000  72.820000 21.085000  96.895000 ;
      RECT 19.800000  96.895000 20.990000  97.500000 ;
      RECT 20.155000  33.335000 20.325000  36.490000 ;
      RECT 20.380000 195.370000 21.090000 195.540000 ;
      RECT 20.935000  29.770000 21.105000  32.860000 ;
      RECT 21.715000  33.340000 21.885000  36.490000 ;
      RECT 21.790000  70.865000 22.680000  97.450000 ;
      RECT 21.810000  97.450000 22.660000 135.315000 ;
      RECT 22.390000 195.370000 23.100000 195.540000 ;
      RECT 22.495000  29.775000 22.665000  32.860000 ;
      RECT 23.025000  90.495000 64.500000  92.990000 ;
      RECT 23.055000 113.340000 64.500000 115.990000 ;
      RECT 23.275000  33.335000 23.445000  36.490000 ;
      RECT 23.510000  68.995000 64.500000  69.990000 ;
      RECT 23.585000  47.515000 24.475000  66.810000 ;
      RECT 23.585000  70.160000 24.615000  89.930000 ;
      RECT 23.585000  93.160000 24.615000 112.930000 ;
      RECT 23.585000 116.160000 24.615000 135.930000 ;
      RECT 23.585000 139.515000 24.475000 158.765000 ;
      RECT 23.585000 162.515000 24.475000 181.765000 ;
      RECT 23.585000 185.515000 24.475000 195.030000 ;
      RECT 24.055000  29.770000 24.225000  32.860000 ;
      RECT 24.835000  33.340000 25.005000  36.490000 ;
      RECT 24.980000  90.370000 64.500000  90.495000 ;
      RECT 24.980000 136.370000 64.500000 136.540000 ;
      RECT 24.980000 195.370000 25.690000 195.540000 ;
      RECT 25.615000  29.775000 25.785000  32.860000 ;
      RECT 25.670000  90.340000 64.500000  90.370000 ;
      RECT 25.670000 136.340000 64.500000 136.370000 ;
      RECT 26.395000  33.335000 26.565000  36.490000 ;
      RECT 26.990000 195.370000 27.700000 195.540000 ;
      RECT 27.175000  29.770000 27.345000  32.860000 ;
      RECT 27.955000  33.340000 28.125000  36.490000 ;
      RECT 28.185000  47.515000 29.075000  66.810000 ;
      RECT 28.185000  70.515000 29.075000  89.810000 ;
      RECT 28.185000  93.515000 29.075000 112.855000 ;
      RECT 28.185000 116.515000 29.075000 135.810000 ;
      RECT 28.185000 139.515000 29.075000 158.765000 ;
      RECT 28.185000 162.515000 29.075000 181.765000 ;
      RECT 28.185000 185.515000 29.075000 195.030000 ;
      RECT 28.735000  29.775000 28.905000  32.860000 ;
      RECT 29.515000  33.335000 29.685000  36.490000 ;
      RECT 29.580000 195.370000 30.290000 195.540000 ;
      RECT 30.295000  29.770000 30.465000  32.860000 ;
      RECT 31.075000  33.340000 31.245000  36.490000 ;
      RECT 31.590000 195.370000 32.300000 195.540000 ;
      RECT 31.855000  29.775000 32.025000  32.860000 ;
      RECT 32.635000  33.335000 32.805000  36.490000 ;
      RECT 32.785000  47.515000 33.675000  66.810000 ;
      RECT 32.785000  70.515000 33.675000  89.765000 ;
      RECT 32.785000  93.515000 33.675000 112.810000 ;
      RECT 32.785000 116.515000 33.675000 135.765000 ;
      RECT 32.785000 139.515000 33.675000 158.765000 ;
      RECT 32.785000 162.515000 33.675000 181.765000 ;
      RECT 32.785000 185.515000 33.675000 195.030000 ;
      RECT 33.415000  29.770000 33.585000  32.860000 ;
      RECT 34.180000 195.370000 34.890000 195.540000 ;
      RECT 34.195000  33.340000 34.365000  36.490000 ;
      RECT 34.975000  29.775000 35.145000  32.860000 ;
      RECT 35.755000  33.335000 35.925000  36.490000 ;
      RECT 36.190000 195.370000 36.900000 195.540000 ;
      RECT 36.535000  29.770000 36.705000  32.860000 ;
      RECT 37.315000  33.340000 37.485000  36.490000 ;
      RECT 37.385000  47.515000 38.275000  66.810000 ;
      RECT 37.385000  70.515000 38.275000  89.765000 ;
      RECT 37.385000  93.515000 38.275000 112.810000 ;
      RECT 37.385000 116.515000 38.275000 135.765000 ;
      RECT 37.385000 139.515000 38.275000 158.765000 ;
      RECT 37.385000 162.515000 38.275000 181.765000 ;
      RECT 37.385000 185.515000 38.275000 195.030000 ;
      RECT 38.095000  29.775000 38.265000  32.860000 ;
      RECT 38.780000 195.370000 39.490000 195.540000 ;
      RECT 38.875000  33.335000 39.045000  36.490000 ;
      RECT 39.655000  29.770000 39.825000  32.860000 ;
      RECT 40.435000  33.335000 40.605000  36.490000 ;
      RECT 40.790000 195.370000 41.500000 195.540000 ;
      RECT 41.215000  29.770000 41.385000  32.860000 ;
      RECT 41.985000  47.515000 42.875000  66.810000 ;
      RECT 41.985000  70.515000 42.875000  89.765000 ;
      RECT 41.985000  93.515000 42.875000 112.810000 ;
      RECT 41.985000 116.515000 42.875000 135.765000 ;
      RECT 41.985000 139.515000 42.875000 158.765000 ;
      RECT 41.985000 162.515000 42.875000 181.765000 ;
      RECT 41.985000 185.515000 42.875000 195.030000 ;
      RECT 41.995000  33.340000 42.165000  36.490000 ;
      RECT 42.775000  29.775000 42.945000  32.860000 ;
      RECT 43.380000 195.370000 44.090000 195.540000 ;
      RECT 43.555000  33.335000 43.725000  36.490000 ;
      RECT 44.335000  29.770000 44.505000  32.860000 ;
      RECT 45.115000  33.340000 45.285000  36.490000 ;
      RECT 45.390000 195.370000 46.100000 195.540000 ;
      RECT 45.755000  29.430000 45.955000  37.425000 ;
      RECT 46.585000  47.515000 47.475000  66.810000 ;
      RECT 46.585000  70.515000 47.475000  89.765000 ;
      RECT 46.585000  93.515000 47.475000 112.810000 ;
      RECT 46.585000 116.515000 47.475000 135.765000 ;
      RECT 46.585000 139.515000 47.475000 158.765000 ;
      RECT 46.585000 162.515000 47.475000 181.765000 ;
      RECT 46.585000 185.515000 47.475000 195.030000 ;
      RECT 47.310000  28.030000 48.200000  29.215000 ;
      RECT 47.310000  29.525000 48.200000  38.695000 ;
      RECT 47.330000  29.215000 48.180000  29.525000 ;
      RECT 47.980000 195.370000 48.690000 195.540000 ;
      RECT 49.990000 195.370000 50.700000 195.540000 ;
      RECT 51.185000  47.515000 52.075000  66.810000 ;
      RECT 51.185000  70.515000 52.075000  89.765000 ;
      RECT 51.185000  93.515000 52.075000 112.810000 ;
      RECT 51.185000 116.515000 52.075000 135.765000 ;
      RECT 51.185000 139.515000 52.075000 158.765000 ;
      RECT 51.185000 162.515000 52.075000 181.765000 ;
      RECT 51.185000 185.515000 52.075000 195.030000 ;
      RECT 52.320000  29.300000 68.865000  31.060000 ;
      RECT 52.320000  31.060000 53.210000  41.455000 ;
      RECT 52.320000  41.455000 68.865000  42.495000 ;
      RECT 52.580000 195.370000 53.290000 195.540000 ;
      RECT 53.960000  31.835000 67.140000  32.005000 ;
      RECT 53.960000  32.005000 54.130000  40.410000 ;
      RECT 53.960000  40.410000 67.140000  40.580000 ;
      RECT 54.590000 195.370000 55.300000 195.540000 ;
      RECT 54.695000  36.190000 54.865000  39.290000 ;
      RECT 54.940000  39.770000 66.335000  39.940000 ;
      RECT 55.215000  23.240000 56.105000  28.345000 ;
      RECT 55.215000  28.345000 70.630000  29.300000 ;
      RECT 55.465000  32.620000 55.635000  35.770000 ;
      RECT 55.785000  47.515000 56.675000  66.810000 ;
      RECT 55.785000  70.515000 56.675000  89.765000 ;
      RECT 55.785000  93.515000 56.675000 112.810000 ;
      RECT 55.785000 116.515000 56.675000 135.765000 ;
      RECT 55.785000 139.515000 56.675000 158.765000 ;
      RECT 55.785000 162.515000 56.675000 181.765000 ;
      RECT 55.785000 185.515000 56.675000 195.140000 ;
      RECT 56.255000  36.190000 56.425000  39.290000 ;
      RECT 56.820000  23.480000 57.050000  27.485000 ;
      RECT 56.820000  27.485000 62.810000  27.715000 ;
      RECT 56.850000  21.465000 57.020000  23.480000 ;
      RECT 57.025000  32.620000 57.195000  35.770000 ;
      RECT 57.180000 195.370000 57.890000 195.540000 ;
      RECT 57.555000  23.480000 57.785000  26.430000 ;
      RECT 57.815000  21.735000 61.815000  21.965000 ;
      RECT 57.815000  36.190000 57.985000  39.290000 ;
      RECT 58.585000  32.620000 58.755000  35.770000 ;
      RECT 59.190000 195.370000 59.900000 195.540000 ;
      RECT 59.375000  36.190000 59.545000  39.290000 ;
      RECT 60.145000  32.620000 60.315000  35.770000 ;
      RECT 60.385000  47.515000 61.275000  66.810000 ;
      RECT 60.385000  70.515000 61.275000  89.765000 ;
      RECT 60.385000  93.515000 61.275000 112.810000 ;
      RECT 60.385000 116.515000 61.275000 135.765000 ;
      RECT 60.385000 139.515000 61.275000 158.765000 ;
      RECT 60.385000 162.515000 61.275000 181.765000 ;
      RECT 60.385000 185.515000 61.275000 195.140000 ;
      RECT 60.935000  36.190000 61.105000  39.290000 ;
      RECT 61.705000  32.620000 61.875000  35.770000 ;
      RECT 61.780000 195.370000 62.490000 195.540000 ;
      RECT 61.850000  23.480000 62.080000  26.430000 ;
      RECT 62.495000  36.190000 62.665000  39.290000 ;
      RECT 62.580000  23.480000 62.810000  27.485000 ;
      RECT 62.610000  21.465000 62.780000  23.480000 ;
      RECT 63.265000  32.620000 63.435000  35.770000 ;
      RECT 63.790000 195.370000 64.500000 195.540000 ;
      RECT 64.055000  36.190000 64.225000  39.290000 ;
      RECT 64.825000  32.620000 64.995000  35.770000 ;
      RECT 64.845000  47.160000 65.875000  66.930000 ;
      RECT 64.845000  70.160000 65.875000  72.950000 ;
      RECT 64.845000  87.140000 65.875000  89.930000 ;
      RECT 64.845000  93.160000 65.875000  95.950000 ;
      RECT 64.845000 110.145000 65.875000 112.935000 ;
      RECT 64.845000 116.160000 65.875000 118.950000 ;
      RECT 64.845000 133.140000 65.875000 135.930000 ;
      RECT 64.845000 139.160000 65.875000 158.930000 ;
      RECT 64.845000 162.160000 65.875000 181.930000 ;
      RECT 64.845000 185.160000 65.875000 195.180000 ;
      RECT 64.985000  72.950000 65.875000  87.140000 ;
      RECT 64.985000  95.950000 65.875000 110.145000 ;
      RECT 64.985000 118.950000 65.875000 133.140000 ;
      RECT 65.615000  36.190000 65.785000  39.290000 ;
      RECT 66.385000  32.620000 66.555000  35.770000 ;
      RECT 66.935000  32.005000 67.140000  36.065000 ;
      RECT 66.935000  36.275000 67.140000  40.410000 ;
      RECT 66.970000  36.065000 67.140000  36.275000 ;
      RECT 67.265000  46.350000 68.155000 101.315000 ;
      RECT 67.265000 166.045000 68.155000 196.835000 ;
      RECT 67.290000 101.315000 68.140000 101.710000 ;
      RECT 67.290000 101.710000 68.155000 165.645000 ;
      RECT 67.290000 165.645000 68.140000 166.045000 ;
      RECT 67.975000  31.060000 68.865000  40.480000 ;
      RECT 67.975000  41.315000 68.865000  41.455000 ;
      RECT 68.000000  40.480000 68.830000  41.315000 ;
      RECT 68.875000  44.755000 70.125000  45.995000 ;
      RECT 68.875000  46.185000 70.125000 198.445000 ;
      RECT 68.905000  45.995000 70.095000  46.185000 ;
      RECT 69.740000  22.520000 70.630000  28.345000 ;
      RECT 69.760000   1.890000 70.650000   2.770000 ;
      RECT 69.765000   3.845000 70.630000   8.915000 ;
      RECT 69.765000   9.845000 70.630000  14.915000 ;
      RECT 69.765000  16.165000 70.630000  21.235000 ;
      RECT 69.780000   2.770000 70.630000   3.845000 ;
      RECT 69.780000   8.915000 70.630000   9.845000 ;
      RECT 69.780000  14.915000 70.630000  16.165000 ;
      RECT 69.780000  21.235000 70.630000  22.520000 ;
      RECT 70.470000  42.820000 71.055000  42.990000 ;
      RECT 70.725000  42.735000 71.055000  42.820000 ;
      RECT 72.245000 199.210000 72.775000 199.380000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  0.215000   2.170000 ;
      RECT  0.000000   0.000000  0.215000   2.170000 ;
      RECT  0.000000   2.170000  0.215000   2.240000 ;
      RECT  0.000000   2.170000  0.725000   2.680000 ;
      RECT  0.000000   2.240000  0.285000   2.310000 ;
      RECT  0.000000   2.310000  0.355000   2.380000 ;
      RECT  0.000000   2.380000  0.425000   2.450000 ;
      RECT  0.000000   2.450000  0.495000   2.520000 ;
      RECT  0.000000   2.520000  0.565000   2.590000 ;
      RECT  0.000000   2.590000  0.635000   2.660000 ;
      RECT  0.000000   2.660000  0.705000   2.680000 ;
      RECT  0.000000   2.680000  0.725000  36.755000 ;
      RECT  0.000000   2.680000  0.725000  36.755000 ;
      RECT  0.000000  36.755000  0.725000  36.800000 ;
      RECT  0.000000  36.755000  0.810000  36.840000 ;
      RECT  0.000000  36.800000  0.770000  36.840000 ;
      RECT  0.000000  36.840000  0.810000  46.930000 ;
      RECT  0.000000  36.840000  0.810000  46.930000 ;
      RECT  0.000000  46.930000  0.725000  47.015000 ;
      RECT  0.000000  46.930000  0.770000  46.970000 ;
      RECT  0.000000  46.970000  0.730000  47.010000 ;
      RECT  0.000000  47.010000  0.725000  47.015000 ;
      RECT  0.000000  47.015000  0.725000 195.355000 ;
      RECT  0.000000  47.015000  0.725000 195.355000 ;
      RECT  0.000000 195.355000 67.480000 200.000000 ;
      RECT  0.000000 195.355000 75.000000 200.000000 ;
      RECT 14.400000  45.430000 57.415000  47.315000 ;
      RECT 14.400000  45.430000 59.035000  45.500000 ;
      RECT 14.400000  45.430000 59.035000  45.500000 ;
      RECT 14.400000  45.500000 58.965000  45.570000 ;
      RECT 14.400000  45.500000 58.965000  45.570000 ;
      RECT 14.400000  45.570000 58.895000  45.640000 ;
      RECT 14.400000  45.570000 58.895000  45.640000 ;
      RECT 14.400000  45.640000 58.825000  45.710000 ;
      RECT 14.400000  45.640000 58.825000  45.710000 ;
      RECT 14.400000  45.710000 58.755000  45.780000 ;
      RECT 14.400000  45.710000 58.755000  45.780000 ;
      RECT 14.400000  45.780000 58.685000  45.850000 ;
      RECT 14.400000  45.780000 58.685000  45.850000 ;
      RECT 14.400000  45.850000 58.615000  45.920000 ;
      RECT 14.400000  45.850000 58.615000  45.920000 ;
      RECT 14.400000  45.920000 58.545000  45.990000 ;
      RECT 14.400000  45.920000 58.545000  45.990000 ;
      RECT 14.400000  45.990000 58.475000  46.060000 ;
      RECT 14.400000  45.990000 58.475000  46.060000 ;
      RECT 14.400000  46.060000 58.405000  46.130000 ;
      RECT 14.400000  46.060000 58.405000  46.130000 ;
      RECT 14.400000  46.130000 58.335000  46.200000 ;
      RECT 14.400000  46.130000 58.335000  46.200000 ;
      RECT 14.400000  46.200000 58.265000  46.270000 ;
      RECT 14.400000  46.200000 58.265000  46.270000 ;
      RECT 14.400000  46.270000 58.195000  46.340000 ;
      RECT 14.400000  46.270000 58.195000  46.340000 ;
      RECT 14.400000  46.340000 58.125000  46.410000 ;
      RECT 14.400000  46.340000 58.125000  46.410000 ;
      RECT 14.400000  46.410000 58.055000  46.480000 ;
      RECT 14.400000  46.410000 58.055000  46.480000 ;
      RECT 14.400000  46.480000 57.985000  46.550000 ;
      RECT 14.400000  46.480000 57.985000  46.550000 ;
      RECT 14.400000  46.550000 57.915000  46.620000 ;
      RECT 14.400000  46.550000 57.915000  46.620000 ;
      RECT 14.400000  46.620000 57.845000  46.690000 ;
      RECT 14.400000  46.620000 57.845000  46.690000 ;
      RECT 14.400000  46.690000 57.775000  46.760000 ;
      RECT 14.400000  46.690000 57.775000  46.760000 ;
      RECT 14.400000  46.760000 57.705000  46.830000 ;
      RECT 14.400000  46.760000 57.705000  46.830000 ;
      RECT 14.400000  46.830000 57.635000  46.900000 ;
      RECT 14.400000  46.830000 57.635000  46.900000 ;
      RECT 14.400000  46.900000 57.565000  46.970000 ;
      RECT 14.400000  46.900000 57.565000  46.970000 ;
      RECT 14.400000  46.970000 57.495000  47.040000 ;
      RECT 14.400000  46.970000 57.495000  47.040000 ;
      RECT 14.400000  47.040000 57.425000  47.110000 ;
      RECT 14.400000  47.040000 57.425000  47.110000 ;
      RECT 14.400000  47.110000 57.360000  47.175000 ;
      RECT 14.400000  47.110000 57.360000  47.175000 ;
      RECT 14.400000  47.175000 16.525000  54.100000 ;
      RECT 14.400000  47.315000 16.665000  54.100000 ;
      RECT 14.400000  54.100000 16.665000  54.905000 ;
      RECT 14.400000  70.140000 57.405000  70.160000 ;
      RECT 14.400000  70.140000 57.405000  70.160000 ;
      RECT 14.400000  70.140000 57.445000  70.315000 ;
      RECT 14.400000  70.160000 57.390000  70.175000 ;
      RECT 14.400000  70.160000 57.390000  70.175000 ;
      RECT 14.400000  70.175000 24.540000  72.870000 ;
      RECT 14.400000  70.315000 24.680000  72.925000 ;
      RECT 14.400000  72.870000 24.470000  72.940000 ;
      RECT 14.400000  72.870000 24.470000  72.940000 ;
      RECT 14.400000  72.925000 23.590000  74.015000 ;
      RECT 14.400000  72.940000 24.400000  73.010000 ;
      RECT 14.400000  72.940000 24.400000  73.010000 ;
      RECT 14.400000  73.010000 24.330000  73.080000 ;
      RECT 14.400000  73.010000 24.330000  73.080000 ;
      RECT 14.400000  73.080000 24.260000  73.150000 ;
      RECT 14.400000  73.080000 24.260000  73.150000 ;
      RECT 14.400000  73.150000 24.190000  73.220000 ;
      RECT 14.400000  73.150000 24.190000  73.220000 ;
      RECT 14.400000  73.220000 24.120000  73.290000 ;
      RECT 14.400000  73.220000 24.120000  73.290000 ;
      RECT 14.400000  73.290000 24.050000  73.360000 ;
      RECT 14.400000  73.290000 24.050000  73.360000 ;
      RECT 14.400000  73.360000 23.980000  73.430000 ;
      RECT 14.400000  73.360000 23.980000  73.430000 ;
      RECT 14.400000  73.430000 23.910000  73.500000 ;
      RECT 14.400000  73.430000 23.910000  73.500000 ;
      RECT 14.400000  73.500000 23.840000  73.570000 ;
      RECT 14.400000  73.500000 23.840000  73.570000 ;
      RECT 14.400000  73.570000 23.770000  73.640000 ;
      RECT 14.400000  73.570000 23.770000  73.640000 ;
      RECT 14.400000  73.640000 23.700000  73.710000 ;
      RECT 14.400000  73.640000 23.700000  73.710000 ;
      RECT 14.400000  73.710000 23.630000  73.780000 ;
      RECT 14.400000  73.710000 23.630000  73.780000 ;
      RECT 14.400000  73.780000 23.560000  73.850000 ;
      RECT 14.400000  73.780000 23.560000  73.850000 ;
      RECT 14.400000  73.850000 23.535000  73.875000 ;
      RECT 14.400000  73.850000 23.535000  73.875000 ;
      RECT 14.400000  73.875000 18.130000  74.695000 ;
      RECT 14.400000  74.015000 18.270000  74.555000 ;
      RECT 14.400000  74.555000 24.680000  75.675000 ;
      RECT 14.400000  74.695000 23.505000  74.765000 ;
      RECT 14.400000  74.695000 23.505000  74.765000 ;
      RECT 14.400000  74.765000 23.575000  74.835000 ;
      RECT 14.400000  74.765000 23.575000  74.835000 ;
      RECT 14.400000  74.835000 23.645000  74.905000 ;
      RECT 14.400000  74.835000 23.645000  74.905000 ;
      RECT 14.400000  74.905000 23.715000  74.975000 ;
      RECT 14.400000  74.905000 23.715000  74.975000 ;
      RECT 14.400000  74.975000 23.785000  75.045000 ;
      RECT 14.400000  74.975000 23.785000  75.045000 ;
      RECT 14.400000  75.045000 23.855000  75.115000 ;
      RECT 14.400000  75.045000 23.855000  75.115000 ;
      RECT 14.400000  75.115000 23.925000  75.185000 ;
      RECT 14.400000  75.115000 23.925000  75.185000 ;
      RECT 14.400000  75.185000 23.995000  75.255000 ;
      RECT 14.400000  75.185000 23.995000  75.255000 ;
      RECT 14.400000  75.255000 24.065000  75.325000 ;
      RECT 14.400000  75.255000 24.065000  75.325000 ;
      RECT 14.400000  75.325000 24.135000  75.395000 ;
      RECT 14.400000  75.325000 24.135000  75.395000 ;
      RECT 14.400000  75.395000 24.205000  75.465000 ;
      RECT 14.400000  75.395000 24.205000  75.465000 ;
      RECT 14.400000  75.465000 24.275000  75.535000 ;
      RECT 14.400000  75.465000 24.275000  75.535000 ;
      RECT 14.400000  75.535000 24.345000  75.605000 ;
      RECT 14.400000  75.535000 24.345000  75.605000 ;
      RECT 14.400000  75.605000 24.415000  75.675000 ;
      RECT 14.400000  75.605000 24.415000  75.675000 ;
      RECT 14.400000  75.675000 24.485000  75.730000 ;
      RECT 14.400000  75.675000 24.485000  75.730000 ;
      RECT 14.400000  75.675000 24.680000  77.125000 ;
      RECT 14.400000  75.730000 24.540000  77.125000 ;
      RECT 14.400000  77.125000 24.680000  79.295000 ;
      RECT 14.400000  93.140000 57.465000  93.160000 ;
      RECT 14.400000  93.140000 57.465000  93.160000 ;
      RECT 14.400000  93.140000 57.505000  93.315000 ;
      RECT 14.400000  93.160000 57.450000  93.175000 ;
      RECT 14.400000  93.160000 57.450000  93.175000 ;
      RECT 14.400000  93.175000 24.540000 100.125000 ;
      RECT 14.400000  93.315000 24.680000 100.125000 ;
      RECT 14.400000 100.125000 24.680000 102.295000 ;
      RECT 14.400000 116.180000 24.540000 123.030000 ;
      RECT 14.400000 116.180000 57.415000 116.315000 ;
      RECT 14.400000 116.315000 24.680000 123.030000 ;
      RECT 14.400000 123.030000 24.680000 125.295000 ;
      RECT 14.400000 139.285000 16.525000 146.100000 ;
      RECT 14.400000 139.285000 57.450000 139.315000 ;
      RECT 14.400000 139.315000 16.665000 146.100000 ;
      RECT 14.400000 146.100000 16.665000 146.770000 ;
      RECT 14.400000 162.195000 16.525000 169.105000 ;
      RECT 14.400000 162.195000 57.465000 162.315000 ;
      RECT 14.400000 162.315000 16.665000 169.105000 ;
      RECT 14.400000 169.105000 16.665000 171.295000 ;
      RECT 14.400000 185.170000 15.340000 189.470000 ;
      RECT 14.400000 185.170000 15.480000 189.470000 ;
      RECT 14.400000 189.470000 15.480000 190.155000 ;
      RECT 14.405000 116.175000 24.540000 116.180000 ;
      RECT 14.405000 116.175000 24.540000 116.180000 ;
      RECT 14.410000 162.185000 16.525000 162.195000 ;
      RECT 14.415000 185.155000 15.340000 185.170000 ;
      RECT 14.415000 185.155000 15.480000 185.170000 ;
      RECT 14.420000  70.120000 57.425000  70.140000 ;
      RECT 14.420000  70.120000 57.425000  70.140000 ;
      RECT 14.420000 162.175000 16.525000 162.185000 ;
      RECT 14.445000  45.385000 59.105000  45.430000 ;
      RECT 14.445000  45.385000 59.105000  45.430000 ;
      RECT 14.455000  93.085000 57.485000  93.140000 ;
      RECT 14.455000  93.085000 57.485000  93.140000 ;
      RECT 14.455000 139.230000 16.525000 139.285000 ;
      RECT 14.460000 116.120000 57.360000 116.175000 ;
      RECT 14.460000 116.120000 57.360000 116.175000 ;
      RECT 14.470000  54.100000 16.525000  54.170000 ;
      RECT 14.470000  77.125000 24.540000  77.195000 ;
      RECT 14.470000  77.125000 24.540000  77.195000 ;
      RECT 14.470000 100.125000 24.540000 100.195000 ;
      RECT 14.470000 100.125000 24.540000 100.195000 ;
      RECT 14.470000 123.030000 24.540000 123.100000 ;
      RECT 14.470000 123.030000 24.540000 123.100000 ;
      RECT 14.470000 146.100000 16.525000 146.170000 ;
      RECT 14.470000 169.105000 16.525000 169.175000 ;
      RECT 14.470000 189.470000 15.340000 189.540000 ;
      RECT 14.475000 162.120000 57.410000 162.175000 ;
      RECT 14.475000 162.120000 57.410000 162.175000 ;
      RECT 14.485000 185.085000 15.340000 185.155000 ;
      RECT 14.490000  70.050000 57.445000  70.120000 ;
      RECT 14.490000  70.050000 57.445000  70.120000 ;
      RECT 14.510000 139.175000 16.525000 139.230000 ;
      RECT 14.515000  45.315000 59.150000  45.385000 ;
      RECT 14.515000  45.315000 59.150000  45.385000 ;
      RECT 14.525000  93.015000 57.540000  93.085000 ;
      RECT 14.525000  93.015000 57.540000  93.085000 ;
      RECT 14.530000 116.050000 57.415000 116.120000 ;
      RECT 14.530000 116.050000 57.415000 116.120000 ;
      RECT 14.540000  54.170000 16.525000  54.240000 ;
      RECT 14.540000  77.195000 24.540000  77.265000 ;
      RECT 14.540000  77.195000 24.540000  77.265000 ;
      RECT 14.540000 100.195000 24.540000 100.265000 ;
      RECT 14.540000 100.195000 24.540000 100.265000 ;
      RECT 14.540000 123.100000 24.540000 123.170000 ;
      RECT 14.540000 123.100000 24.540000 123.170000 ;
      RECT 14.540000 146.170000 16.525000 146.240000 ;
      RECT 14.540000 169.175000 16.525000 169.245000 ;
      RECT 14.540000 189.540000 15.340000 189.610000 ;
      RECT 14.545000 162.050000 57.465000 162.120000 ;
      RECT 14.545000 162.050000 57.465000 162.120000 ;
      RECT 14.555000 185.015000 15.340000 185.085000 ;
      RECT 14.560000  69.980000 57.515000  70.050000 ;
      RECT 14.560000  69.980000 57.515000  70.050000 ;
      RECT 14.565000 139.120000 57.395000 139.175000 ;
      RECT 14.565000 139.120000 57.395000 139.175000 ;
      RECT 14.565000 185.005000 58.580000 185.015000 ;
      RECT 14.585000  45.245000 59.220000  45.315000 ;
      RECT 14.585000  45.245000 59.220000  45.315000 ;
      RECT 14.595000  92.945000 57.610000  93.015000 ;
      RECT 14.595000  92.945000 57.610000  93.015000 ;
      RECT 14.600000 115.980000 57.485000 116.050000 ;
      RECT 14.600000 115.980000 57.485000 116.050000 ;
      RECT 14.610000  54.240000 16.525000  54.310000 ;
      RECT 14.610000  77.265000 24.540000  77.335000 ;
      RECT 14.610000  77.265000 24.540000  77.335000 ;
      RECT 14.610000 100.265000 24.540000 100.335000 ;
      RECT 14.610000 100.265000 24.540000 100.335000 ;
      RECT 14.610000 123.170000 24.540000 123.240000 ;
      RECT 14.610000 123.170000 24.540000 123.240000 ;
      RECT 14.610000 146.240000 16.525000 146.310000 ;
      RECT 14.610000 169.245000 16.525000 169.315000 ;
      RECT 14.610000 189.610000 15.340000 189.680000 ;
      RECT 14.615000 161.980000 57.535000 162.050000 ;
      RECT 14.615000 161.980000 57.535000 162.050000 ;
      RECT 14.630000  69.910000 57.585000  69.980000 ;
      RECT 14.630000  69.910000 57.585000  69.980000 ;
      RECT 14.635000 139.050000 57.450000 139.120000 ;
      RECT 14.635000 139.050000 57.450000 139.120000 ;
      RECT 14.635000 184.935000 58.590000 185.005000 ;
      RECT 14.655000  45.175000 59.290000  45.245000 ;
      RECT 14.655000  45.175000 59.290000  45.245000 ;
      RECT 14.665000  92.875000 57.680000  92.945000 ;
      RECT 14.665000  92.875000 57.680000  92.945000 ;
      RECT 14.670000 115.910000 57.555000 115.980000 ;
      RECT 14.670000 115.910000 57.555000 115.980000 ;
      RECT 14.680000  54.310000 16.525000  54.380000 ;
      RECT 14.680000  77.335000 24.540000  77.405000 ;
      RECT 14.680000  77.335000 24.540000  77.405000 ;
      RECT 14.680000 100.335000 24.540000 100.405000 ;
      RECT 14.680000 100.335000 24.540000 100.405000 ;
      RECT 14.680000 123.240000 24.540000 123.310000 ;
      RECT 14.680000 123.240000 24.540000 123.310000 ;
      RECT 14.680000 146.310000 16.525000 146.380000 ;
      RECT 14.680000 169.315000 16.525000 169.385000 ;
      RECT 14.680000 189.680000 15.340000 189.750000 ;
      RECT 14.685000 161.910000 57.605000 161.980000 ;
      RECT 14.685000 161.910000 57.605000 161.980000 ;
      RECT 14.700000  69.840000 57.655000  69.910000 ;
      RECT 14.700000  69.840000 57.655000  69.910000 ;
      RECT 14.705000 138.980000 57.520000 139.050000 ;
      RECT 14.705000 138.980000 57.520000 139.050000 ;
      RECT 14.705000 184.865000 58.660000 184.935000 ;
      RECT 14.725000  45.105000 59.360000  45.175000 ;
      RECT 14.725000  45.105000 59.360000  45.175000 ;
      RECT 14.735000  92.805000 57.750000  92.875000 ;
      RECT 14.735000  92.805000 57.750000  92.875000 ;
      RECT 14.740000 115.840000 57.625000 115.910000 ;
      RECT 14.740000 115.840000 57.625000 115.910000 ;
      RECT 14.750000  54.380000 16.525000  54.450000 ;
      RECT 14.750000  77.405000 24.540000  77.475000 ;
      RECT 14.750000  77.405000 24.540000  77.475000 ;
      RECT 14.750000 100.405000 24.540000 100.475000 ;
      RECT 14.750000 100.405000 24.540000 100.475000 ;
      RECT 14.750000 123.310000 24.540000 123.380000 ;
      RECT 14.750000 123.310000 24.540000 123.380000 ;
      RECT 14.750000 146.380000 16.525000 146.450000 ;
      RECT 14.750000 169.385000 16.525000 169.455000 ;
      RECT 14.750000 189.750000 15.340000 189.820000 ;
      RECT 14.755000 161.840000 57.675000 161.910000 ;
      RECT 14.755000 161.840000 57.675000 161.910000 ;
      RECT 14.770000  69.770000 57.725000  69.840000 ;
      RECT 14.770000  69.770000 57.725000  69.840000 ;
      RECT 14.775000 138.910000 57.590000 138.980000 ;
      RECT 14.775000 138.910000 57.590000 138.980000 ;
      RECT 14.775000 184.795000 58.730000 184.865000 ;
      RECT 14.795000  45.035000 59.430000  45.105000 ;
      RECT 14.795000  45.035000 59.430000  45.105000 ;
      RECT 14.805000  92.735000 57.820000  92.805000 ;
      RECT 14.805000  92.735000 57.820000  92.805000 ;
      RECT 14.810000 115.770000 57.695000 115.840000 ;
      RECT 14.810000 115.770000 57.695000 115.840000 ;
      RECT 14.820000  54.450000 16.525000  54.520000 ;
      RECT 14.820000  77.475000 24.540000  77.545000 ;
      RECT 14.820000  77.475000 24.540000  77.545000 ;
      RECT 14.820000 100.475000 24.540000 100.545000 ;
      RECT 14.820000 100.475000 24.540000 100.545000 ;
      RECT 14.820000 123.380000 24.540000 123.450000 ;
      RECT 14.820000 123.380000 24.540000 123.450000 ;
      RECT 14.820000 146.450000 16.525000 146.520000 ;
      RECT 14.820000 169.455000 16.525000 169.525000 ;
      RECT 14.820000 189.820000 15.340000 189.890000 ;
      RECT 14.825000 161.770000 57.745000 161.840000 ;
      RECT 14.825000 161.770000 57.745000 161.840000 ;
      RECT 14.840000  69.700000 57.795000  69.770000 ;
      RECT 14.840000  69.700000 57.795000  69.770000 ;
      RECT 14.845000 138.840000 57.660000 138.910000 ;
      RECT 14.845000 138.840000 57.660000 138.910000 ;
      RECT 14.845000 184.725000 58.800000 184.795000 ;
      RECT 14.865000  44.965000 59.500000  45.035000 ;
      RECT 14.865000  44.965000 59.500000  45.035000 ;
      RECT 14.875000  92.665000 57.890000  92.735000 ;
      RECT 14.875000  92.665000 57.890000  92.735000 ;
      RECT 14.880000 115.700000 57.765000 115.770000 ;
      RECT 14.880000 115.700000 57.765000 115.770000 ;
      RECT 14.890000  54.520000 16.525000  54.590000 ;
      RECT 14.890000  77.545000 24.540000  77.615000 ;
      RECT 14.890000  77.545000 24.540000  77.615000 ;
      RECT 14.890000 100.545000 24.540000 100.615000 ;
      RECT 14.890000 100.545000 24.540000 100.615000 ;
      RECT 14.890000 123.450000 24.540000 123.520000 ;
      RECT 14.890000 123.450000 24.540000 123.520000 ;
      RECT 14.890000 146.520000 16.525000 146.590000 ;
      RECT 14.890000 169.525000 16.525000 169.595000 ;
      RECT 14.890000 189.890000 15.340000 189.960000 ;
      RECT 14.895000 161.700000 57.815000 161.770000 ;
      RECT 14.895000 161.700000 57.815000 161.770000 ;
      RECT 14.910000  69.630000 57.865000  69.700000 ;
      RECT 14.910000  69.630000 57.865000  69.700000 ;
      RECT 14.915000 138.770000 57.730000 138.840000 ;
      RECT 14.915000 138.770000 57.730000 138.840000 ;
      RECT 14.915000 184.655000 58.870000 184.725000 ;
      RECT 14.935000  44.895000 59.570000  44.965000 ;
      RECT 14.935000  44.895000 59.570000  44.965000 ;
      RECT 14.945000  92.595000 57.960000  92.665000 ;
      RECT 14.945000  92.595000 57.960000  92.665000 ;
      RECT 14.950000 115.630000 57.835000 115.700000 ;
      RECT 14.950000 115.630000 57.835000 115.700000 ;
      RECT 14.960000  54.590000 16.525000  54.660000 ;
      RECT 14.960000  77.615000 24.540000  77.685000 ;
      RECT 14.960000  77.615000 24.540000  77.685000 ;
      RECT 14.960000 100.615000 24.540000 100.685000 ;
      RECT 14.960000 100.615000 24.540000 100.685000 ;
      RECT 14.960000 123.520000 24.540000 123.590000 ;
      RECT 14.960000 123.520000 24.540000 123.590000 ;
      RECT 14.960000 146.590000 16.525000 146.660000 ;
      RECT 14.960000 169.595000 16.525000 169.665000 ;
      RECT 14.960000 189.960000 15.340000 190.030000 ;
      RECT 14.965000 161.630000 57.885000 161.700000 ;
      RECT 14.965000 161.630000 57.885000 161.700000 ;
      RECT 14.980000  69.560000 57.935000  69.630000 ;
      RECT 14.980000  69.560000 57.935000  69.630000 ;
      RECT 14.985000 138.700000 57.800000 138.770000 ;
      RECT 14.985000 138.700000 57.800000 138.770000 ;
      RECT 14.985000 184.585000 58.940000 184.655000 ;
      RECT 15.005000  44.825000 59.640000  44.895000 ;
      RECT 15.005000  44.825000 59.640000  44.895000 ;
      RECT 15.015000  92.525000 58.030000  92.595000 ;
      RECT 15.015000  92.525000 58.030000  92.595000 ;
      RECT 15.020000 115.560000 57.905000 115.630000 ;
      RECT 15.020000 115.560000 57.905000 115.630000 ;
      RECT 15.030000  54.660000 16.525000  54.730000 ;
      RECT 15.030000  77.685000 24.540000  77.755000 ;
      RECT 15.030000  77.685000 24.540000  77.755000 ;
      RECT 15.030000 100.685000 24.540000 100.755000 ;
      RECT 15.030000 100.685000 24.540000 100.755000 ;
      RECT 15.030000 123.590000 24.540000 123.660000 ;
      RECT 15.030000 123.590000 24.540000 123.660000 ;
      RECT 15.030000 146.660000 16.525000 146.730000 ;
      RECT 15.030000 169.665000 16.525000 169.735000 ;
      RECT 15.030000 190.030000 15.340000 190.100000 ;
      RECT 15.035000 161.560000 57.955000 161.630000 ;
      RECT 15.035000 161.560000 57.955000 161.630000 ;
      RECT 15.050000  69.490000 58.005000  69.560000 ;
      RECT 15.050000  69.490000 58.005000  69.560000 ;
      RECT 15.055000 138.630000 57.870000 138.700000 ;
      RECT 15.055000 138.630000 57.870000 138.700000 ;
      RECT 15.055000 184.515000 59.010000 184.585000 ;
      RECT 15.070000 146.770000 18.190000 148.295000 ;
      RECT 15.075000  44.755000 59.710000  44.825000 ;
      RECT 15.075000  44.755000 59.710000  44.825000 ;
      RECT 15.085000  92.455000 58.100000  92.525000 ;
      RECT 15.085000  92.455000 58.100000  92.525000 ;
      RECT 15.085000 190.155000 75.000000 190.280000 ;
      RECT 15.090000 115.490000 57.975000 115.560000 ;
      RECT 15.090000 115.490000 57.975000 115.560000 ;
      RECT 15.100000  54.730000 16.525000  54.800000 ;
      RECT 15.100000  77.755000 24.540000  77.825000 ;
      RECT 15.100000  77.755000 24.540000  77.825000 ;
      RECT 15.100000 100.755000 24.540000 100.825000 ;
      RECT 15.100000 100.755000 24.540000 100.825000 ;
      RECT 15.100000 123.660000 24.540000 123.730000 ;
      RECT 15.100000 123.660000 24.540000 123.730000 ;
      RECT 15.100000 146.730000 16.525000 146.800000 ;
      RECT 15.100000 169.735000 16.525000 169.805000 ;
      RECT 15.100000 190.100000 15.340000 190.170000 ;
      RECT 15.105000 161.490000 58.025000 161.560000 ;
      RECT 15.105000 161.490000 58.025000 161.560000 ;
      RECT 15.120000  69.420000 58.075000  69.490000 ;
      RECT 15.120000  69.420000 58.075000  69.490000 ;
      RECT 15.125000 138.560000 57.940000 138.630000 ;
      RECT 15.125000 138.560000 57.940000 138.630000 ;
      RECT 15.125000 146.800000 16.525000 146.825000 ;
      RECT 15.125000 184.445000 59.080000 184.515000 ;
      RECT 15.145000  44.685000 59.780000  44.755000 ;
      RECT 15.145000  44.685000 59.780000  44.755000 ;
      RECT 15.155000  92.385000 58.170000  92.455000 ;
      RECT 15.155000  92.385000 58.170000  92.455000 ;
      RECT 15.160000 115.420000 58.045000 115.490000 ;
      RECT 15.160000 115.420000 58.045000 115.490000 ;
      RECT 15.170000  54.800000 16.525000  54.870000 ;
      RECT 15.170000  77.825000 24.540000  77.895000 ;
      RECT 15.170000  77.825000 24.540000  77.895000 ;
      RECT 15.170000 100.825000 24.540000 100.895000 ;
      RECT 15.170000 100.825000 24.540000 100.895000 ;
      RECT 15.170000 123.730000 24.540000 123.800000 ;
      RECT 15.170000 123.730000 24.540000 123.800000 ;
      RECT 15.170000 169.805000 16.525000 169.875000 ;
      RECT 15.170000 190.170000 15.340000 190.240000 ;
      RECT 15.175000 161.420000 58.095000 161.490000 ;
      RECT 15.175000 161.420000 58.095000 161.490000 ;
      RECT 15.190000  69.350000 58.145000  69.420000 ;
      RECT 15.190000  69.350000 58.145000  69.420000 ;
      RECT 15.195000 138.490000 58.010000 138.560000 ;
      RECT 15.195000 138.490000 58.010000 138.560000 ;
      RECT 15.195000 146.825000 16.525000 146.895000 ;
      RECT 15.195000 184.375000 59.150000 184.445000 ;
      RECT 15.205000  54.905000 18.790000  56.295000 ;
      RECT 15.210000 190.240000 15.340000 190.280000 ;
      RECT 15.215000  44.615000 59.850000  44.685000 ;
      RECT 15.215000  44.615000 59.850000  44.685000 ;
      RECT 15.225000  92.315000 58.240000  92.385000 ;
      RECT 15.225000  92.315000 58.240000  92.385000 ;
      RECT 15.230000 115.350000 58.115000 115.420000 ;
      RECT 15.230000 115.350000 58.115000 115.420000 ;
      RECT 15.240000  54.870000 16.525000  54.940000 ;
      RECT 15.240000  77.895000 24.540000  77.965000 ;
      RECT 15.240000  77.895000 24.540000  77.965000 ;
      RECT 15.240000 100.895000 24.540000 100.965000 ;
      RECT 15.240000 100.895000 24.540000 100.965000 ;
      RECT 15.240000 123.800000 24.540000 123.870000 ;
      RECT 15.240000 123.800000 24.540000 123.870000 ;
      RECT 15.240000 169.875000 16.525000 169.945000 ;
      RECT 15.245000 161.350000 58.165000 161.420000 ;
      RECT 15.245000 161.350000 58.165000 161.420000 ;
      RECT 15.260000  69.280000 58.215000  69.350000 ;
      RECT 15.260000  69.280000 58.215000  69.350000 ;
      RECT 15.265000 138.420000 58.080000 138.490000 ;
      RECT 15.265000 138.420000 58.080000 138.490000 ;
      RECT 15.265000 146.895000 16.595000 146.965000 ;
      RECT 15.265000 184.305000 59.220000 184.375000 ;
      RECT 15.285000  44.545000 59.920000  44.615000 ;
      RECT 15.285000  44.545000 59.920000  44.615000 ;
      RECT 15.295000  92.245000 58.310000  92.315000 ;
      RECT 15.295000  92.245000 58.310000  92.315000 ;
      RECT 15.300000 115.280000 58.185000 115.350000 ;
      RECT 15.300000 115.280000 58.185000 115.350000 ;
      RECT 15.310000  54.940000 16.525000  55.010000 ;
      RECT 15.310000  77.965000 24.540000  78.035000 ;
      RECT 15.310000  77.965000 24.540000  78.035000 ;
      RECT 15.310000 100.965000 24.540000 101.035000 ;
      RECT 15.310000 100.965000 24.540000 101.035000 ;
      RECT 15.310000 123.870000 24.540000 123.940000 ;
      RECT 15.310000 123.870000 24.540000 123.940000 ;
      RECT 15.310000 169.945000 16.525000 170.015000 ;
      RECT 15.315000 161.280000 58.235000 161.350000 ;
      RECT 15.315000 161.280000 58.235000 161.350000 ;
      RECT 15.330000  69.210000 58.285000  69.280000 ;
      RECT 15.330000  69.210000 58.285000  69.280000 ;
      RECT 15.335000 138.350000 58.150000 138.420000 ;
      RECT 15.335000 138.350000 58.150000 138.420000 ;
      RECT 15.335000 146.965000 16.665000 147.035000 ;
      RECT 15.335000 184.235000 59.290000 184.305000 ;
      RECT 15.345000  55.010000 16.525000  55.045000 ;
      RECT 15.355000  44.475000 59.990000  44.545000 ;
      RECT 15.355000  44.475000 59.990000  44.545000 ;
      RECT 15.365000  92.175000 58.380000  92.245000 ;
      RECT 15.365000  92.175000 58.380000  92.245000 ;
      RECT 15.370000 115.210000 58.255000 115.280000 ;
      RECT 15.370000 115.210000 58.255000 115.280000 ;
      RECT 15.380000  78.035000 24.540000  78.105000 ;
      RECT 15.380000  78.035000 24.540000  78.105000 ;
      RECT 15.380000 101.035000 24.540000 101.105000 ;
      RECT 15.380000 101.035000 24.540000 101.105000 ;
      RECT 15.380000 123.940000 24.540000 124.010000 ;
      RECT 15.380000 123.940000 24.540000 124.010000 ;
      RECT 15.380000 170.015000 16.525000 170.085000 ;
      RECT 15.385000 161.210000 58.305000 161.280000 ;
      RECT 15.385000 161.210000 58.305000 161.280000 ;
      RECT 15.400000  69.140000 58.355000  69.210000 ;
      RECT 15.400000  69.140000 58.355000  69.210000 ;
      RECT 15.405000 138.280000 58.220000 138.350000 ;
      RECT 15.405000 138.280000 58.220000 138.350000 ;
      RECT 15.405000 147.035000 16.735000 147.105000 ;
      RECT 15.405000 184.165000 59.360000 184.235000 ;
      RECT 15.415000  55.045000 17.345000  55.115000 ;
      RECT 15.425000  44.405000 60.060000  44.475000 ;
      RECT 15.425000  44.405000 60.060000  44.475000 ;
      RECT 15.435000  92.105000 58.450000  92.175000 ;
      RECT 15.435000  92.105000 58.450000  92.175000 ;
      RECT 15.440000 115.140000 58.325000 115.210000 ;
      RECT 15.440000 115.140000 58.325000 115.210000 ;
      RECT 15.450000  78.105000 24.540000  78.175000 ;
      RECT 15.450000  78.105000 24.540000  78.175000 ;
      RECT 15.450000 101.105000 24.540000 101.175000 ;
      RECT 15.450000 101.105000 24.540000 101.175000 ;
      RECT 15.450000 124.010000 24.540000 124.080000 ;
      RECT 15.450000 124.010000 24.540000 124.080000 ;
      RECT 15.450000 170.085000 16.525000 170.155000 ;
      RECT 15.455000 161.140000 58.375000 161.210000 ;
      RECT 15.455000 161.140000 58.375000 161.210000 ;
      RECT 15.470000  69.070000 58.425000  69.140000 ;
      RECT 15.470000  69.070000 58.425000  69.140000 ;
      RECT 15.475000 138.210000 58.290000 138.280000 ;
      RECT 15.475000 138.210000 58.290000 138.280000 ;
      RECT 15.475000 147.105000 16.805000 147.175000 ;
      RECT 15.475000 184.095000 59.430000 184.165000 ;
      RECT 15.485000  29.430000 59.190000  29.500000 ;
      RECT 15.485000  29.430000 59.190000  29.500000 ;
      RECT 15.485000  29.430000 60.970000  31.015000 ;
      RECT 15.485000  29.500000 59.260000  29.570000 ;
      RECT 15.485000  29.500000 59.260000  29.570000 ;
      RECT 15.485000  29.570000 59.330000  29.640000 ;
      RECT 15.485000  29.570000 59.330000  29.640000 ;
      RECT 15.485000  29.640000 59.400000  29.710000 ;
      RECT 15.485000  29.640000 59.400000  29.710000 ;
      RECT 15.485000  29.710000 59.470000  29.780000 ;
      RECT 15.485000  29.710000 59.470000  29.780000 ;
      RECT 15.485000  29.780000 59.540000  29.850000 ;
      RECT 15.485000  29.780000 59.540000  29.850000 ;
      RECT 15.485000  29.850000 59.610000  29.920000 ;
      RECT 15.485000  29.850000 59.610000  29.920000 ;
      RECT 15.485000  29.920000 59.680000  29.990000 ;
      RECT 15.485000  29.920000 59.680000  29.990000 ;
      RECT 15.485000  29.990000 59.750000  30.060000 ;
      RECT 15.485000  29.990000 59.750000  30.060000 ;
      RECT 15.485000  30.060000 59.820000  30.130000 ;
      RECT 15.485000  30.060000 59.820000  30.130000 ;
      RECT 15.485000  30.130000 59.890000  30.200000 ;
      RECT 15.485000  30.130000 59.890000  30.200000 ;
      RECT 15.485000  30.200000 59.960000  30.270000 ;
      RECT 15.485000  30.200000 59.960000  30.270000 ;
      RECT 15.485000  30.270000 60.030000  30.340000 ;
      RECT 15.485000  30.270000 60.030000  30.340000 ;
      RECT 15.485000  30.340000 60.100000  30.410000 ;
      RECT 15.485000  30.340000 60.100000  30.410000 ;
      RECT 15.485000  30.410000 60.170000  30.480000 ;
      RECT 15.485000  30.410000 60.170000  30.480000 ;
      RECT 15.485000  30.480000 60.240000  30.550000 ;
      RECT 15.485000  30.480000 60.240000  30.550000 ;
      RECT 15.485000  30.550000 60.310000  30.620000 ;
      RECT 15.485000  30.550000 60.310000  30.620000 ;
      RECT 15.485000  30.620000 60.380000  30.690000 ;
      RECT 15.485000  30.620000 60.380000  30.690000 ;
      RECT 15.485000  30.690000 60.450000  30.760000 ;
      RECT 15.485000  30.690000 60.450000  30.760000 ;
      RECT 15.485000  30.760000 60.520000  30.830000 ;
      RECT 15.485000  30.760000 60.520000  30.830000 ;
      RECT 15.485000  30.830000 60.590000  30.900000 ;
      RECT 15.485000  30.830000 60.590000  30.900000 ;
      RECT 15.485000  30.900000 60.660000  30.970000 ;
      RECT 15.485000  30.900000 60.660000  30.970000 ;
      RECT 15.485000  30.970000 60.730000  31.040000 ;
      RECT 15.485000  30.970000 60.730000  31.040000 ;
      RECT 15.485000  31.015000 60.970000  35.550000 ;
      RECT 15.485000  31.040000 60.800000  31.070000 ;
      RECT 15.485000  31.040000 60.800000  31.070000 ;
      RECT 15.485000  31.070000 60.830000  35.550000 ;
      RECT 15.485000  35.550000 60.970000  35.975000 ;
      RECT 15.485000  55.115000 17.415000  55.185000 ;
      RECT 15.495000  44.335000 60.130000  44.405000 ;
      RECT 15.495000  44.335000 60.130000  44.405000 ;
      RECT 15.505000  29.410000 59.170000  29.430000 ;
      RECT 15.505000  29.410000 59.170000  29.430000 ;
      RECT 15.505000  92.035000 58.520000  92.105000 ;
      RECT 15.505000  92.035000 58.520000  92.105000 ;
      RECT 15.510000 115.070000 58.395000 115.140000 ;
      RECT 15.510000 115.070000 58.395000 115.140000 ;
      RECT 15.520000  78.175000 24.540000  78.245000 ;
      RECT 15.520000  78.175000 24.540000  78.245000 ;
      RECT 15.520000 101.175000 24.540000 101.245000 ;
      RECT 15.520000 101.175000 24.540000 101.245000 ;
      RECT 15.520000 124.080000 24.540000 124.150000 ;
      RECT 15.520000 124.080000 24.540000 124.150000 ;
      RECT 15.520000 170.155000 16.525000 170.225000 ;
      RECT 15.525000 161.070000 58.445000 161.140000 ;
      RECT 15.525000 161.070000 58.445000 161.140000 ;
      RECT 15.540000  69.000000 58.495000  69.070000 ;
      RECT 15.540000  69.000000 58.495000  69.070000 ;
      RECT 15.545000 138.140000 58.360000 138.210000 ;
      RECT 15.545000 138.140000 58.360000 138.210000 ;
      RECT 15.545000 147.175000 16.875000 147.245000 ;
      RECT 15.545000 184.025000 59.500000 184.095000 ;
      RECT 15.555000  35.550000 60.830000  35.620000 ;
      RECT 15.555000  35.550000 60.830000  35.620000 ;
      RECT 15.555000  55.185000 17.485000  55.255000 ;
      RECT 15.565000  44.265000 60.200000  44.335000 ;
      RECT 15.565000  44.265000 60.200000  44.335000 ;
      RECT 15.575000  29.340000 59.100000  29.410000 ;
      RECT 15.575000  29.340000 59.100000  29.410000 ;
      RECT 15.575000  91.965000 58.590000  92.035000 ;
      RECT 15.575000  91.965000 58.590000  92.035000 ;
      RECT 15.580000 115.000000 58.465000 115.070000 ;
      RECT 15.580000 115.000000 58.465000 115.070000 ;
      RECT 15.590000  78.245000 24.540000  78.315000 ;
      RECT 15.590000  78.245000 24.540000  78.315000 ;
      RECT 15.590000 101.245000 24.540000 101.315000 ;
      RECT 15.590000 101.245000 24.540000 101.315000 ;
      RECT 15.590000 124.150000 24.540000 124.220000 ;
      RECT 15.590000 124.150000 24.540000 124.220000 ;
      RECT 15.590000 170.225000 16.525000 170.295000 ;
      RECT 15.595000 161.000000 58.515000 161.070000 ;
      RECT 15.595000 161.000000 58.515000 161.070000 ;
      RECT 15.610000  68.930000 58.565000  69.000000 ;
      RECT 15.610000  68.930000 58.565000  69.000000 ;
      RECT 15.615000 138.070000 58.430000 138.140000 ;
      RECT 15.615000 138.070000 58.430000 138.140000 ;
      RECT 15.615000 147.245000 16.945000 147.315000 ;
      RECT 15.615000 183.955000 59.570000 184.025000 ;
      RECT 15.625000  35.620000 60.830000  35.690000 ;
      RECT 15.625000  35.620000 60.830000  35.690000 ;
      RECT 15.625000  55.255000 17.555000  55.325000 ;
      RECT 15.635000  44.195000 60.270000  44.265000 ;
      RECT 15.635000  44.195000 60.270000  44.265000 ;
      RECT 15.645000  29.270000 59.030000  29.340000 ;
      RECT 15.645000  29.270000 59.030000  29.340000 ;
      RECT 15.645000  91.895000 58.660000  91.965000 ;
      RECT 15.645000  91.895000 58.660000  91.965000 ;
      RECT 15.650000 114.930000 58.535000 115.000000 ;
      RECT 15.650000 114.930000 58.535000 115.000000 ;
      RECT 15.660000  78.315000 24.540000  78.385000 ;
      RECT 15.660000  78.315000 24.540000  78.385000 ;
      RECT 15.660000 101.315000 24.540000 101.385000 ;
      RECT 15.660000 101.315000 24.540000 101.385000 ;
      RECT 15.660000 124.220000 24.540000 124.290000 ;
      RECT 15.660000 124.220000 24.540000 124.290000 ;
      RECT 15.660000 170.295000 16.525000 170.365000 ;
      RECT 15.665000 160.930000 58.585000 161.000000 ;
      RECT 15.665000 160.930000 58.585000 161.000000 ;
      RECT 15.680000  68.860000 58.635000  68.930000 ;
      RECT 15.680000  68.860000 58.635000  68.930000 ;
      RECT 15.685000 138.000000 58.500000 138.070000 ;
      RECT 15.685000 138.000000 58.500000 138.070000 ;
      RECT 15.685000 147.315000 17.015000 147.385000 ;
      RECT 15.685000 183.885000 59.640000 183.955000 ;
      RECT 15.695000  35.690000 60.830000  35.760000 ;
      RECT 15.695000  35.690000 60.830000  35.760000 ;
      RECT 15.695000  55.325000 17.625000  55.395000 ;
      RECT 15.705000  44.125000 60.340000  44.195000 ;
      RECT 15.705000  44.125000 60.340000  44.195000 ;
      RECT 15.715000  29.200000 58.960000  29.270000 ;
      RECT 15.715000  29.200000 58.960000  29.270000 ;
      RECT 15.715000  91.825000 58.730000  91.895000 ;
      RECT 15.715000  91.825000 58.730000  91.895000 ;
      RECT 15.720000 114.860000 58.605000 114.930000 ;
      RECT 15.720000 114.860000 58.605000 114.930000 ;
      RECT 15.730000  78.385000 24.540000  78.455000 ;
      RECT 15.730000  78.385000 24.540000  78.455000 ;
      RECT 15.730000 101.385000 24.540000 101.455000 ;
      RECT 15.730000 101.385000 24.540000 101.455000 ;
      RECT 15.730000 124.290000 24.540000 124.360000 ;
      RECT 15.730000 124.290000 24.540000 124.360000 ;
      RECT 15.730000 170.365000 16.525000 170.435000 ;
      RECT 15.735000 160.860000 58.655000 160.930000 ;
      RECT 15.735000 160.860000 58.655000 160.930000 ;
      RECT 15.750000  68.790000 58.705000  68.860000 ;
      RECT 15.750000  68.790000 58.705000  68.860000 ;
      RECT 15.755000 137.930000 58.570000 138.000000 ;
      RECT 15.755000 137.930000 58.570000 138.000000 ;
      RECT 15.755000 147.385000 17.085000 147.455000 ;
      RECT 15.755000 183.815000 59.710000 183.885000 ;
      RECT 15.765000  35.760000 60.830000  35.830000 ;
      RECT 15.765000  35.760000 60.830000  35.830000 ;
      RECT 15.765000  55.395000 17.695000  55.465000 ;
      RECT 15.770000  35.830000 60.830000  35.835000 ;
      RECT 15.770000  35.830000 60.830000  35.835000 ;
      RECT 15.775000  44.055000 60.410000  44.125000 ;
      RECT 15.775000  44.055000 60.410000  44.125000 ;
      RECT 15.785000  29.130000 58.890000  29.200000 ;
      RECT 15.785000  29.130000 58.890000  29.200000 ;
      RECT 15.785000  91.755000 58.800000  91.825000 ;
      RECT 15.785000  91.755000 58.800000  91.825000 ;
      RECT 15.790000 114.790000 58.675000 114.860000 ;
      RECT 15.790000 114.790000 58.675000 114.860000 ;
      RECT 15.800000  78.455000 24.540000  78.525000 ;
      RECT 15.800000  78.455000 24.540000  78.525000 ;
      RECT 15.800000 101.455000 24.540000 101.525000 ;
      RECT 15.800000 101.455000 24.540000 101.525000 ;
      RECT 15.800000 124.360000 24.540000 124.430000 ;
      RECT 15.800000 124.360000 24.540000 124.430000 ;
      RECT 15.800000 170.435000 16.525000 170.505000 ;
      RECT 15.805000 160.790000 58.725000 160.860000 ;
      RECT 15.805000 160.790000 58.725000 160.860000 ;
      RECT 15.820000  68.720000 58.775000  68.790000 ;
      RECT 15.820000  68.720000 58.775000  68.790000 ;
      RECT 15.825000 137.860000 58.640000 137.930000 ;
      RECT 15.825000 137.860000 58.640000 137.930000 ;
      RECT 15.825000 147.455000 17.155000 147.525000 ;
      RECT 15.825000 183.745000 59.780000 183.815000 ;
      RECT 15.835000  55.465000 17.765000  55.535000 ;
      RECT 15.840000  35.835000 54.390000  35.905000 ;
      RECT 15.840000  35.835000 54.390000  35.905000 ;
      RECT 15.845000  43.985000 60.480000  44.055000 ;
      RECT 15.845000  43.985000 60.480000  44.055000 ;
      RECT 15.855000  29.060000 58.820000  29.130000 ;
      RECT 15.855000  29.060000 58.820000  29.130000 ;
      RECT 15.855000  91.685000 58.870000  91.755000 ;
      RECT 15.855000  91.685000 58.870000  91.755000 ;
      RECT 15.860000 114.720000 58.745000 114.790000 ;
      RECT 15.860000 114.720000 58.745000 114.790000 ;
      RECT 15.870000  78.525000 24.540000  78.595000 ;
      RECT 15.870000  78.525000 24.540000  78.595000 ;
      RECT 15.870000 101.525000 24.540000 101.595000 ;
      RECT 15.870000 101.525000 24.540000 101.595000 ;
      RECT 15.870000 124.430000 24.540000 124.500000 ;
      RECT 15.870000 124.430000 24.540000 124.500000 ;
      RECT 15.870000 170.505000 16.525000 170.575000 ;
      RECT 15.875000 160.720000 58.795000 160.790000 ;
      RECT 15.875000 160.720000 58.795000 160.790000 ;
      RECT 15.890000  68.650000 58.845000  68.720000 ;
      RECT 15.890000  68.650000 58.845000  68.720000 ;
      RECT 15.895000 137.790000 58.710000 137.860000 ;
      RECT 15.895000 137.790000 58.710000 137.860000 ;
      RECT 15.895000 147.525000 17.225000 147.595000 ;
      RECT 15.895000 183.675000 59.850000 183.745000 ;
      RECT 15.905000  55.535000 17.835000  55.605000 ;
      RECT 15.910000  35.905000 54.390000  35.975000 ;
      RECT 15.910000  35.905000 54.390000  35.975000 ;
      RECT 15.910000  35.975000 54.530000  38.195000 ;
      RECT 15.915000  43.915000 60.550000  43.985000 ;
      RECT 15.915000  43.915000 60.550000  43.985000 ;
      RECT 15.925000  28.990000 58.750000  29.060000 ;
      RECT 15.925000  28.990000 58.750000  29.060000 ;
      RECT 15.925000  91.615000 58.940000  91.685000 ;
      RECT 15.925000  91.615000 58.940000  91.685000 ;
      RECT 15.930000 114.650000 58.815000 114.720000 ;
      RECT 15.930000 114.650000 58.815000 114.720000 ;
      RECT 15.940000  78.595000 24.540000  78.665000 ;
      RECT 15.940000  78.595000 24.540000  78.665000 ;
      RECT 15.940000 101.595000 24.540000 101.665000 ;
      RECT 15.940000 101.595000 24.540000 101.665000 ;
      RECT 15.940000 124.500000 24.540000 124.570000 ;
      RECT 15.940000 124.500000 24.540000 124.570000 ;
      RECT 15.940000 170.575000 16.525000 170.645000 ;
      RECT 15.945000 160.650000 58.865000 160.720000 ;
      RECT 15.945000 160.650000 58.865000 160.720000 ;
      RECT 15.960000  68.580000 58.915000  68.650000 ;
      RECT 15.960000  68.580000 58.915000  68.650000 ;
      RECT 15.965000 137.720000 58.780000 137.790000 ;
      RECT 15.965000 137.720000 58.780000 137.790000 ;
      RECT 15.965000 147.595000 17.295000 147.665000 ;
      RECT 15.965000 183.605000 59.920000 183.675000 ;
      RECT 15.975000  55.605000 17.905000  55.675000 ;
      RECT 15.980000  35.975000 54.390000  36.045000 ;
      RECT 15.980000  35.975000 54.390000  36.045000 ;
      RECT 15.985000  43.845000 60.620000  43.915000 ;
      RECT 15.985000  43.845000 60.620000  43.915000 ;
      RECT 15.995000  28.920000 58.680000  28.990000 ;
      RECT 15.995000  28.920000 58.680000  28.990000 ;
      RECT 15.995000  91.545000 59.010000  91.615000 ;
      RECT 15.995000  91.545000 59.010000  91.615000 ;
      RECT 16.000000 114.580000 58.885000 114.650000 ;
      RECT 16.000000 114.580000 58.885000 114.650000 ;
      RECT 16.010000  78.665000 24.540000  78.735000 ;
      RECT 16.010000  78.665000 24.540000  78.735000 ;
      RECT 16.010000 101.665000 24.540000 101.735000 ;
      RECT 16.010000 101.665000 24.540000 101.735000 ;
      RECT 16.010000 124.570000 24.540000 124.640000 ;
      RECT 16.010000 124.570000 24.540000 124.640000 ;
      RECT 16.010000 170.645000 16.525000 170.715000 ;
      RECT 16.015000 160.580000 58.935000 160.650000 ;
      RECT 16.015000 160.580000 58.935000 160.650000 ;
      RECT 16.030000  68.510000 58.985000  68.580000 ;
      RECT 16.030000  68.510000 58.985000  68.580000 ;
      RECT 16.035000 137.650000 58.850000 137.720000 ;
      RECT 16.035000 137.650000 58.850000 137.720000 ;
      RECT 16.035000 147.665000 17.365000 147.735000 ;
      RECT 16.035000 183.535000 59.990000 183.605000 ;
      RECT 16.045000  55.675000 17.975000  55.745000 ;
      RECT 16.050000  36.045000 54.390000  36.115000 ;
      RECT 16.050000  36.045000 54.390000  36.115000 ;
      RECT 16.055000  43.775000 60.690000  43.845000 ;
      RECT 16.055000  43.775000 60.690000  43.845000 ;
      RECT 16.065000  28.850000 58.610000  28.920000 ;
      RECT 16.065000  28.850000 58.610000  28.920000 ;
      RECT 16.065000  91.475000 59.080000  91.545000 ;
      RECT 16.065000  91.475000 59.080000  91.545000 ;
      RECT 16.070000  43.760000 59.300000  45.430000 ;
      RECT 16.070000 114.510000 58.955000 114.580000 ;
      RECT 16.070000 114.510000 58.955000 114.580000 ;
      RECT 16.080000  78.735000 24.540000  78.805000 ;
      RECT 16.080000  78.735000 24.540000  78.805000 ;
      RECT 16.080000 101.735000 24.540000 101.805000 ;
      RECT 16.080000 101.735000 24.540000 101.805000 ;
      RECT 16.080000 124.640000 24.540000 124.710000 ;
      RECT 16.080000 124.640000 24.540000 124.710000 ;
      RECT 16.080000 170.715000 16.525000 170.785000 ;
      RECT 16.085000 160.510000 59.005000 160.580000 ;
      RECT 16.085000 160.510000 59.005000 160.580000 ;
      RECT 16.100000  68.440000 59.055000  68.510000 ;
      RECT 16.100000  68.440000 59.055000  68.510000 ;
      RECT 16.105000 137.580000 58.920000 137.650000 ;
      RECT 16.105000 137.580000 58.920000 137.650000 ;
      RECT 16.105000 147.735000 17.435000 147.805000 ;
      RECT 16.105000 183.465000 60.060000 183.535000 ;
      RECT 16.115000  55.745000 18.045000  55.815000 ;
      RECT 16.120000  36.115000 54.390000  36.185000 ;
      RECT 16.120000  36.115000 54.390000  36.185000 ;
      RECT 16.125000  43.705000 60.760000  43.775000 ;
      RECT 16.125000  43.705000 60.760000  43.775000 ;
      RECT 16.135000  28.780000 58.540000  28.850000 ;
      RECT 16.135000  28.780000 58.540000  28.850000 ;
      RECT 16.135000  91.405000 59.150000  91.475000 ;
      RECT 16.135000  91.405000 59.150000  91.475000 ;
      RECT 16.140000 114.440000 59.025000 114.510000 ;
      RECT 16.140000 114.440000 59.025000 114.510000 ;
      RECT 16.150000  78.805000 24.540000  78.875000 ;
      RECT 16.150000  78.805000 24.540000  78.875000 ;
      RECT 16.150000 101.805000 24.540000 101.875000 ;
      RECT 16.150000 101.805000 24.540000 101.875000 ;
      RECT 16.150000 124.710000 24.540000 124.780000 ;
      RECT 16.150000 124.710000 24.540000 124.780000 ;
      RECT 16.150000 170.785000 16.525000 170.855000 ;
      RECT 16.155000 160.440000 59.075000 160.510000 ;
      RECT 16.155000 160.440000 59.075000 160.510000 ;
      RECT 16.170000  68.370000 59.125000  68.440000 ;
      RECT 16.170000  68.370000 59.125000  68.440000 ;
      RECT 16.175000 137.510000 58.990000 137.580000 ;
      RECT 16.175000 137.510000 58.990000 137.580000 ;
      RECT 16.175000 147.805000 17.505000 147.875000 ;
      RECT 16.175000 183.395000 60.130000 183.465000 ;
      RECT 16.185000  55.815000 18.115000  55.885000 ;
      RECT 16.190000  36.185000 54.390000  36.255000 ;
      RECT 16.190000  36.185000 54.390000  36.255000 ;
      RECT 16.190000  43.640000 60.830000  43.705000 ;
      RECT 16.190000  43.640000 60.830000  43.705000 ;
      RECT 16.205000  28.710000 58.470000  28.780000 ;
      RECT 16.205000  28.710000 58.470000  28.780000 ;
      RECT 16.205000  91.335000 59.220000  91.405000 ;
      RECT 16.205000  91.335000 59.220000  91.405000 ;
      RECT 16.210000 114.370000 59.095000 114.440000 ;
      RECT 16.210000 114.370000 59.095000 114.440000 ;
      RECT 16.220000  78.875000 24.540000  78.945000 ;
      RECT 16.220000  78.875000 24.540000  78.945000 ;
      RECT 16.220000 101.875000 24.540000 101.945000 ;
      RECT 16.220000 101.875000 24.540000 101.945000 ;
      RECT 16.220000 124.780000 24.540000 124.850000 ;
      RECT 16.220000 124.780000 24.540000 124.850000 ;
      RECT 16.220000 170.855000 16.525000 170.925000 ;
      RECT 16.225000 160.370000 59.145000 160.440000 ;
      RECT 16.225000 160.370000 59.145000 160.440000 ;
      RECT 16.240000  68.300000 59.195000  68.370000 ;
      RECT 16.240000  68.300000 59.195000  68.370000 ;
      RECT 16.245000 137.440000 59.060000 137.510000 ;
      RECT 16.245000 137.440000 59.060000 137.510000 ;
      RECT 16.245000 147.875000 17.575000 147.945000 ;
      RECT 16.245000 183.325000 60.200000 183.395000 ;
      RECT 16.255000  55.885000 18.185000  55.955000 ;
      RECT 16.260000  36.255000 54.390000  36.325000 ;
      RECT 16.260000  36.255000 54.390000  36.325000 ;
      RECT 16.260000  43.570000 60.830000  43.640000 ;
      RECT 16.260000  43.570000 60.830000  43.640000 ;
      RECT 16.275000  28.640000 58.400000  28.710000 ;
      RECT 16.275000  28.640000 58.400000  28.710000 ;
      RECT 16.275000  91.265000 59.290000  91.335000 ;
      RECT 16.275000  91.265000 59.290000  91.335000 ;
      RECT 16.280000 114.300000 59.165000 114.370000 ;
      RECT 16.280000 114.300000 59.165000 114.370000 ;
      RECT 16.290000  78.945000 24.540000  79.015000 ;
      RECT 16.290000  78.945000 24.540000  79.015000 ;
      RECT 16.290000 101.945000 24.540000 102.015000 ;
      RECT 16.290000 101.945000 24.540000 102.015000 ;
      RECT 16.290000 124.850000 24.540000 124.920000 ;
      RECT 16.290000 124.850000 24.540000 124.920000 ;
      RECT 16.290000 170.925000 16.525000 170.995000 ;
      RECT 16.295000 160.300000 59.215000 160.370000 ;
      RECT 16.295000 160.300000 59.215000 160.370000 ;
      RECT 16.310000  68.230000 59.265000  68.300000 ;
      RECT 16.310000  68.230000 59.265000  68.300000 ;
      RECT 16.315000 137.370000 59.130000 137.440000 ;
      RECT 16.315000 137.370000 59.130000 137.440000 ;
      RECT 16.315000 147.945000 17.645000 148.015000 ;
      RECT 16.315000 183.255000 60.270000 183.325000 ;
      RECT 16.325000  55.955000 18.255000  56.025000 ;
      RECT 16.330000  36.325000 54.390000  36.395000 ;
      RECT 16.330000  36.325000 54.390000  36.395000 ;
      RECT 16.330000  43.500000 60.830000  43.570000 ;
      RECT 16.330000  43.500000 60.830000  43.570000 ;
      RECT 16.345000  28.570000 58.330000  28.640000 ;
      RECT 16.345000  28.570000 58.330000  28.640000 ;
      RECT 16.345000  91.195000 59.360000  91.265000 ;
      RECT 16.345000  91.195000 59.360000  91.265000 ;
      RECT 16.350000 114.230000 59.235000 114.300000 ;
      RECT 16.350000 114.230000 59.235000 114.300000 ;
      RECT 16.360000  79.015000 24.540000  79.085000 ;
      RECT 16.360000  79.015000 24.540000  79.085000 ;
      RECT 16.360000 102.015000 24.540000 102.085000 ;
      RECT 16.360000 102.015000 24.540000 102.085000 ;
      RECT 16.360000 124.920000 24.540000 124.990000 ;
      RECT 16.360000 124.920000 24.540000 124.990000 ;
      RECT 16.360000 170.995000 16.525000 171.065000 ;
      RECT 16.365000 160.230000 59.285000 160.300000 ;
      RECT 16.365000 160.230000 59.285000 160.300000 ;
      RECT 16.380000  68.160000 59.335000  68.230000 ;
      RECT 16.380000  68.160000 59.335000  68.230000 ;
      RECT 16.385000 137.300000 59.200000 137.370000 ;
      RECT 16.385000 137.300000 59.200000 137.370000 ;
      RECT 16.385000 148.015000 17.715000 148.085000 ;
      RECT 16.385000 183.185000 60.340000 183.255000 ;
      RECT 16.395000  56.025000 18.325000  56.095000 ;
      RECT 16.400000  36.395000 54.390000  36.465000 ;
      RECT 16.400000  36.395000 54.390000  36.465000 ;
      RECT 16.400000  43.430000 60.830000  43.500000 ;
      RECT 16.400000  43.430000 60.830000  43.500000 ;
      RECT 16.415000  28.500000 58.260000  28.570000 ;
      RECT 16.415000  28.500000 58.260000  28.570000 ;
      RECT 16.415000  91.125000 59.430000  91.195000 ;
      RECT 16.415000  91.125000 59.430000  91.195000 ;
      RECT 16.420000 114.160000 59.305000 114.230000 ;
      RECT 16.420000 114.160000 59.305000 114.230000 ;
      RECT 16.430000  79.085000 24.540000  79.155000 ;
      RECT 16.430000  79.085000 24.540000  79.155000 ;
      RECT 16.430000 102.085000 24.540000 102.155000 ;
      RECT 16.430000 102.085000 24.540000 102.155000 ;
      RECT 16.430000 124.990000 24.540000 125.060000 ;
      RECT 16.430000 124.990000 24.540000 125.060000 ;
      RECT 16.430000 171.065000 16.525000 171.135000 ;
      RECT 16.435000 160.160000 59.355000 160.230000 ;
      RECT 16.435000 160.160000 59.355000 160.230000 ;
      RECT 16.450000  68.090000 59.405000  68.160000 ;
      RECT 16.450000  68.090000 59.405000  68.160000 ;
      RECT 16.455000 137.230000 59.270000 137.300000 ;
      RECT 16.455000 137.230000 59.270000 137.300000 ;
      RECT 16.455000 148.085000 17.785000 148.155000 ;
      RECT 16.455000 183.115000 60.410000 183.185000 ;
      RECT 16.465000  56.095000 18.395000  56.165000 ;
      RECT 16.470000  36.465000 54.390000  36.535000 ;
      RECT 16.470000  36.465000 54.390000  36.535000 ;
      RECT 16.470000  43.360000 60.830000  43.430000 ;
      RECT 16.470000  43.360000 60.830000  43.430000 ;
      RECT 16.485000  28.430000 58.190000  28.500000 ;
      RECT 16.485000  28.430000 58.190000  28.500000 ;
      RECT 16.485000  91.055000 59.500000  91.125000 ;
      RECT 16.485000  91.055000 59.500000  91.125000 ;
      RECT 16.490000 114.090000 59.375000 114.160000 ;
      RECT 16.490000 114.090000 59.375000 114.160000 ;
      RECT 16.500000  79.155000 24.540000  79.225000 ;
      RECT 16.500000  79.155000 24.540000  79.225000 ;
      RECT 16.500000 102.155000 24.540000 102.225000 ;
      RECT 16.500000 102.155000 24.540000 102.225000 ;
      RECT 16.500000 125.060000 24.540000 125.130000 ;
      RECT 16.500000 125.060000 24.540000 125.130000 ;
      RECT 16.500000 171.135000 16.525000 171.205000 ;
      RECT 16.505000 160.090000 59.425000 160.160000 ;
      RECT 16.505000 160.090000 59.425000 160.160000 ;
      RECT 16.520000  68.020000 59.475000  68.090000 ;
      RECT 16.520000  68.020000 59.475000  68.090000 ;
      RECT 16.525000 137.160000 59.340000 137.230000 ;
      RECT 16.525000 137.160000 59.340000 137.230000 ;
      RECT 16.525000 148.155000 17.855000 148.225000 ;
      RECT 16.525000 183.045000 60.480000 183.115000 ;
      RECT 16.535000  56.165000 18.465000  56.235000 ;
      RECT 16.540000  36.535000 54.390000  36.605000 ;
      RECT 16.540000  36.535000 54.390000  36.605000 ;
      RECT 16.540000  43.290000 60.830000  43.360000 ;
      RECT 16.540000  43.290000 60.830000  43.360000 ;
      RECT 16.555000  28.360000 58.120000  28.430000 ;
      RECT 16.555000  28.360000 58.120000  28.430000 ;
      RECT 16.555000  90.985000 59.570000  91.055000 ;
      RECT 16.555000  90.985000 59.570000  91.055000 ;
      RECT 16.560000 114.020000 59.445000 114.090000 ;
      RECT 16.560000 114.020000 59.445000 114.090000 ;
      RECT 16.570000  79.225000 24.540000  79.295000 ;
      RECT 16.570000  79.225000 24.540000  79.295000 ;
      RECT 16.570000  79.295000 58.700000  80.500000 ;
      RECT 16.570000 102.225000 24.540000 102.295000 ;
      RECT 16.570000 102.225000 24.540000 102.295000 ;
      RECT 16.570000 102.295000 58.700000 103.500000 ;
      RECT 16.570000 125.130000 24.540000 125.200000 ;
      RECT 16.570000 125.130000 24.540000 125.200000 ;
      RECT 16.575000 160.020000 59.495000 160.090000 ;
      RECT 16.575000 160.020000 59.495000 160.090000 ;
      RECT 16.590000  67.950000 59.545000  68.020000 ;
      RECT 16.590000  67.950000 59.545000  68.020000 ;
      RECT 16.590000 171.295000 58.710000 172.500000 ;
      RECT 16.595000  56.295000 58.670000  57.500000 ;
      RECT 16.595000 137.090000 59.410000 137.160000 ;
      RECT 16.595000 137.090000 59.410000 137.160000 ;
      RECT 16.595000 148.225000 17.925000 148.295000 ;
      RECT 16.595000 148.295000 58.630000 149.500000 ;
      RECT 16.595000 182.975000 60.550000 183.045000 ;
      RECT 16.605000  56.235000 18.535000  56.305000 ;
      RECT 16.610000  36.605000 54.390000  36.675000 ;
      RECT 16.610000  36.605000 54.390000  36.675000 ;
      RECT 16.610000  43.220000 60.830000  43.290000 ;
      RECT 16.610000  43.220000 60.830000  43.290000 ;
      RECT 16.625000  28.290000 58.050000  28.360000 ;
      RECT 16.625000  28.290000 58.050000  28.360000 ;
      RECT 16.625000  90.915000 59.640000  90.985000 ;
      RECT 16.625000  90.915000 59.640000  90.985000 ;
      RECT 16.630000 113.950000 59.515000 114.020000 ;
      RECT 16.630000 113.950000 59.515000 114.020000 ;
      RECT 16.640000  79.295000 24.540000  79.365000 ;
      RECT 16.640000  79.295000 24.540000  79.365000 ;
      RECT 16.640000 102.295000 24.540000 102.365000 ;
      RECT 16.640000 102.295000 24.540000 102.365000 ;
      RECT 16.640000 125.200000 24.540000 125.270000 ;
      RECT 16.640000 125.200000 24.540000 125.270000 ;
      RECT 16.645000 159.950000 59.565000 160.020000 ;
      RECT 16.645000 159.950000 59.565000 160.020000 ;
      RECT 16.660000  67.880000 59.615000  67.950000 ;
      RECT 16.660000  67.880000 59.615000  67.950000 ;
      RECT 16.665000 125.295000 58.700000 126.500000 ;
      RECT 16.665000 137.020000 59.480000 137.090000 ;
      RECT 16.665000 137.020000 59.480000 137.090000 ;
      RECT 16.665000 148.295000 17.995000 148.365000 ;
      RECT 16.665000 182.905000 60.620000 182.975000 ;
      RECT 16.675000  56.305000 18.605000  56.375000 ;
      RECT 16.680000  36.675000 54.390000  36.745000 ;
      RECT 16.680000  36.675000 54.390000  36.745000 ;
      RECT 16.680000  43.150000 60.830000  43.220000 ;
      RECT 16.680000  43.150000 60.830000  43.220000 ;
      RECT 16.695000  28.220000 57.980000  28.290000 ;
      RECT 16.695000  28.220000 57.980000  28.290000 ;
      RECT 16.695000  90.845000 59.710000  90.915000 ;
      RECT 16.695000  90.845000 59.710000  90.915000 ;
      RECT 16.700000 113.880000 59.585000 113.950000 ;
      RECT 16.700000 113.880000 59.585000 113.950000 ;
      RECT 16.710000  79.365000 24.540000  79.435000 ;
      RECT 16.710000  79.365000 24.540000  79.435000 ;
      RECT 16.710000 102.365000 24.540000 102.435000 ;
      RECT 16.710000 102.365000 24.540000 102.435000 ;
      RECT 16.710000 125.270000 24.540000 125.340000 ;
      RECT 16.710000 125.270000 24.540000 125.340000 ;
      RECT 16.715000 159.880000 59.635000 159.950000 ;
      RECT 16.715000 159.880000 59.635000 159.950000 ;
      RECT 16.730000  67.810000 59.685000  67.880000 ;
      RECT 16.730000  67.810000 59.685000  67.880000 ;
      RECT 16.735000  56.375000 18.675000  56.435000 ;
      RECT 16.735000 136.950000 59.550000 137.020000 ;
      RECT 16.735000 136.950000 59.550000 137.020000 ;
      RECT 16.735000 148.365000 18.065000 148.435000 ;
      RECT 16.735000 182.835000 60.690000 182.905000 ;
      RECT 16.750000  36.745000 54.390000  36.815000 ;
      RECT 16.750000  36.745000 54.390000  36.815000 ;
      RECT 16.750000  43.080000 60.830000  43.150000 ;
      RECT 16.750000  43.080000 60.830000  43.150000 ;
      RECT 16.750000 182.820000 58.635000 185.155000 ;
      RECT 16.765000  28.150000 57.910000  28.220000 ;
      RECT 16.765000  28.150000 57.910000  28.220000 ;
      RECT 16.765000  90.775000 59.780000  90.845000 ;
      RECT 16.765000  90.775000 59.780000  90.845000 ;
      RECT 16.770000 113.810000 59.655000 113.880000 ;
      RECT 16.770000 113.810000 59.655000 113.880000 ;
      RECT 16.780000  79.435000 24.540000  79.505000 ;
      RECT 16.780000  79.435000 24.540000  79.505000 ;
      RECT 16.780000  79.435000 57.440000  79.505000 ;
      RECT 16.780000 102.435000 24.540000 102.505000 ;
      RECT 16.780000 102.435000 24.540000 102.505000 ;
      RECT 16.780000 102.435000 57.440000 102.505000 ;
      RECT 16.780000 125.340000 24.540000 125.410000 ;
      RECT 16.780000 125.340000 24.540000 125.410000 ;
      RECT 16.785000 159.810000 59.705000 159.880000 ;
      RECT 16.785000 159.810000 59.705000 159.880000 ;
      RECT 16.800000  67.740000 59.755000  67.810000 ;
      RECT 16.800000  67.740000 59.755000  67.810000 ;
      RECT 16.800000 171.435000 57.450000 171.505000 ;
      RECT 16.805000  56.435000 57.410000  56.505000 ;
      RECT 16.805000 125.410000 24.540000 125.435000 ;
      RECT 16.805000 125.410000 24.540000 125.435000 ;
      RECT 16.805000 136.880000 59.620000 136.950000 ;
      RECT 16.805000 136.880000 59.620000 136.950000 ;
      RECT 16.805000 148.435000 57.370000 148.505000 ;
      RECT 16.805000 182.765000 60.760000 182.835000 ;
      RECT 16.820000  36.815000 54.390000  36.885000 ;
      RECT 16.820000  36.815000 54.390000  36.885000 ;
      RECT 16.820000  43.010000 60.830000  43.080000 ;
      RECT 16.820000  43.010000 60.830000  43.080000 ;
      RECT 16.830000 182.740000 60.830000 182.765000 ;
      RECT 16.835000  28.080000 57.840000  28.150000 ;
      RECT 16.835000  28.080000 57.840000  28.150000 ;
      RECT 16.835000  90.705000 59.850000  90.775000 ;
      RECT 16.835000  90.705000 59.850000  90.775000 ;
      RECT 16.840000 113.740000 59.725000 113.810000 ;
      RECT 16.840000 113.740000 59.725000 113.810000 ;
      RECT 16.850000  79.505000 24.540000  79.575000 ;
      RECT 16.850000  79.505000 24.540000  79.575000 ;
      RECT 16.850000  79.505000 57.510000  79.575000 ;
      RECT 16.850000 102.505000 24.540000 102.575000 ;
      RECT 16.850000 102.505000 24.540000 102.575000 ;
      RECT 16.850000 102.505000 57.510000 102.575000 ;
      RECT 16.855000 159.740000 59.775000 159.810000 ;
      RECT 16.855000 159.740000 59.775000 159.810000 ;
      RECT 16.870000  67.670000 59.825000  67.740000 ;
      RECT 16.870000  67.670000 59.825000  67.740000 ;
      RECT 16.870000 171.505000 57.520000 171.575000 ;
      RECT 16.875000  56.505000 57.480000  56.575000 ;
      RECT 16.875000 125.435000 24.540000 125.505000 ;
      RECT 16.875000 125.435000 24.540000 125.505000 ;
      RECT 16.875000 125.435000 57.440000 125.505000 ;
      RECT 16.875000 136.810000 59.690000 136.880000 ;
      RECT 16.875000 136.810000 59.690000 136.880000 ;
      RECT 16.875000 148.505000 57.440000 148.575000 ;
      RECT 16.890000  36.885000 54.390000  36.955000 ;
      RECT 16.890000  36.885000 54.390000  36.955000 ;
      RECT 16.890000  42.940000 60.830000  43.010000 ;
      RECT 16.890000  42.940000 60.830000  43.010000 ;
      RECT 16.900000 182.670000 60.830000 182.740000 ;
      RECT 16.905000  28.010000 57.770000  28.080000 ;
      RECT 16.905000  28.010000 57.770000  28.080000 ;
      RECT 16.905000  90.635000 59.920000  90.705000 ;
      RECT 16.905000  90.635000 59.920000  90.705000 ;
      RECT 16.910000 113.670000 59.795000 113.740000 ;
      RECT 16.910000 113.670000 59.795000 113.740000 ;
      RECT 16.920000  79.575000 24.540000  79.645000 ;
      RECT 16.920000  79.575000 24.540000  79.645000 ;
      RECT 16.920000  79.575000 57.580000  79.645000 ;
      RECT 16.920000 102.575000 24.540000 102.645000 ;
      RECT 16.920000 102.575000 24.540000 102.645000 ;
      RECT 16.920000 102.575000 57.580000 102.645000 ;
      RECT 16.925000 159.670000 59.845000 159.740000 ;
      RECT 16.925000 159.670000 59.845000 159.740000 ;
      RECT 16.940000  67.600000 59.895000  67.670000 ;
      RECT 16.940000  67.600000 59.895000  67.670000 ;
      RECT 16.940000 171.575000 57.590000 171.645000 ;
      RECT 16.945000  56.575000 57.550000  56.645000 ;
      RECT 16.945000 125.505000 24.540000 125.575000 ;
      RECT 16.945000 125.505000 24.540000 125.575000 ;
      RECT 16.945000 125.505000 57.510000 125.575000 ;
      RECT 16.945000 136.740000 59.760000 136.810000 ;
      RECT 16.945000 136.740000 59.760000 136.810000 ;
      RECT 16.945000 148.575000 57.510000 148.645000 ;
      RECT 16.960000  36.955000 54.390000  37.025000 ;
      RECT 16.960000  36.955000 54.390000  37.025000 ;
      RECT 16.960000  42.870000 60.830000  42.940000 ;
      RECT 16.960000  42.870000 60.830000  42.940000 ;
      RECT 16.970000 182.600000 60.830000 182.670000 ;
      RECT 16.975000  27.940000 57.700000  28.010000 ;
      RECT 16.975000  27.940000 57.700000  28.010000 ;
      RECT 16.975000  90.565000 59.990000  90.635000 ;
      RECT 16.975000  90.565000 59.990000  90.635000 ;
      RECT 16.980000 113.600000 59.865000 113.670000 ;
      RECT 16.980000 113.600000 59.865000 113.670000 ;
      RECT 16.990000  79.645000 24.540000  79.715000 ;
      RECT 16.990000  79.645000 24.540000  79.715000 ;
      RECT 16.990000  79.645000 57.650000  79.715000 ;
      RECT 16.990000 102.645000 24.540000 102.715000 ;
      RECT 16.990000 102.645000 24.540000 102.715000 ;
      RECT 16.990000 102.645000 57.650000 102.715000 ;
      RECT 16.995000 159.600000 59.915000 159.670000 ;
      RECT 16.995000 159.600000 59.915000 159.670000 ;
      RECT 17.010000  67.530000 59.965000  67.600000 ;
      RECT 17.010000  67.530000 59.965000  67.600000 ;
      RECT 17.010000 171.645000 57.660000 171.715000 ;
      RECT 17.015000  56.645000 57.620000  56.715000 ;
      RECT 17.015000 125.575000 24.540000 125.645000 ;
      RECT 17.015000 125.575000 24.540000 125.645000 ;
      RECT 17.015000 125.575000 57.580000 125.645000 ;
      RECT 17.015000 136.670000 59.830000 136.740000 ;
      RECT 17.015000 136.670000 59.830000 136.740000 ;
      RECT 17.015000 148.645000 57.580000 148.715000 ;
      RECT 17.030000  37.025000 54.390000  37.095000 ;
      RECT 17.030000  37.025000 54.390000  37.095000 ;
      RECT 17.030000  42.800000 60.830000  42.870000 ;
      RECT 17.030000  42.800000 60.830000  42.870000 ;
      RECT 17.040000 182.530000 60.830000 182.600000 ;
      RECT 17.045000  27.870000 57.630000  27.940000 ;
      RECT 17.045000  27.870000 57.630000  27.940000 ;
      RECT 17.045000  90.495000 60.060000  90.565000 ;
      RECT 17.045000  90.495000 60.060000  90.565000 ;
      RECT 17.050000 113.530000 59.935000 113.600000 ;
      RECT 17.050000 113.530000 59.935000 113.600000 ;
      RECT 17.060000  79.715000 24.540000  79.785000 ;
      RECT 17.060000  79.715000 24.540000  79.785000 ;
      RECT 17.060000  79.715000 57.720000  79.785000 ;
      RECT 17.060000 102.715000 24.540000 102.785000 ;
      RECT 17.060000 102.715000 24.540000 102.785000 ;
      RECT 17.060000 102.715000 57.720000 102.785000 ;
      RECT 17.065000 159.530000 59.985000 159.600000 ;
      RECT 17.065000 159.530000 59.985000 159.600000 ;
      RECT 17.080000  67.460000 60.035000  67.530000 ;
      RECT 17.080000  67.460000 60.035000  67.530000 ;
      RECT 17.080000 171.715000 57.730000 171.785000 ;
      RECT 17.085000  56.715000 57.690000  56.785000 ;
      RECT 17.085000 125.645000 24.540000 125.715000 ;
      RECT 17.085000 125.645000 24.540000 125.715000 ;
      RECT 17.085000 125.645000 57.650000 125.715000 ;
      RECT 17.085000 136.600000 59.900000 136.670000 ;
      RECT 17.085000 136.600000 59.900000 136.670000 ;
      RECT 17.085000 148.715000 57.650000 148.785000 ;
      RECT 17.100000  37.095000 54.390000  37.165000 ;
      RECT 17.100000  37.095000 54.390000  37.165000 ;
      RECT 17.100000  42.730000 60.830000  42.800000 ;
      RECT 17.100000  42.730000 60.830000  42.800000 ;
      RECT 17.110000 182.460000 60.830000 182.530000 ;
      RECT 17.115000  27.800000 57.560000  27.870000 ;
      RECT 17.115000  27.800000 57.560000  27.870000 ;
      RECT 17.115000  90.425000 60.130000  90.495000 ;
      RECT 17.115000  90.425000 60.130000  90.495000 ;
      RECT 17.120000 113.460000 60.005000 113.530000 ;
      RECT 17.120000 113.460000 60.005000 113.530000 ;
      RECT 17.130000  79.785000 24.540000  79.855000 ;
      RECT 17.130000  79.785000 24.540000  79.855000 ;
      RECT 17.130000  79.785000 57.790000  79.855000 ;
      RECT 17.130000 102.785000 24.540000 102.855000 ;
      RECT 17.130000 102.785000 24.540000 102.855000 ;
      RECT 17.130000 102.785000 57.790000 102.855000 ;
      RECT 17.135000 159.460000 60.055000 159.530000 ;
      RECT 17.135000 159.460000 60.055000 159.530000 ;
      RECT 17.150000  67.390000 60.105000  67.460000 ;
      RECT 17.150000  67.390000 60.105000  67.460000 ;
      RECT 17.150000 171.785000 57.800000 171.855000 ;
      RECT 17.155000  56.785000 57.760000  56.855000 ;
      RECT 17.155000 125.715000 24.540000 125.785000 ;
      RECT 17.155000 125.715000 24.540000 125.785000 ;
      RECT 17.155000 125.715000 57.720000 125.785000 ;
      RECT 17.155000 136.530000 59.970000 136.600000 ;
      RECT 17.155000 136.530000 59.970000 136.600000 ;
      RECT 17.155000 148.785000 57.720000 148.855000 ;
      RECT 17.170000  37.165000 54.390000  37.235000 ;
      RECT 17.170000  37.165000 54.390000  37.235000 ;
      RECT 17.170000  42.660000 60.830000  42.730000 ;
      RECT 17.170000  42.660000 60.830000  42.730000 ;
      RECT 17.170000  42.660000 60.970000  43.760000 ;
      RECT 17.180000 182.390000 60.830000 182.460000 ;
      RECT 17.185000  27.730000 57.490000  27.800000 ;
      RECT 17.185000  27.730000 57.490000  27.800000 ;
      RECT 17.185000  90.355000 60.200000  90.425000 ;
      RECT 17.185000  90.355000 60.200000  90.425000 ;
      RECT 17.190000 113.390000 60.075000 113.460000 ;
      RECT 17.190000 113.390000 60.075000 113.460000 ;
      RECT 17.200000  79.855000 24.540000  79.925000 ;
      RECT 17.200000  79.855000 24.540000  79.925000 ;
      RECT 17.200000  79.855000 57.860000  79.925000 ;
      RECT 17.200000 102.855000 24.540000 102.925000 ;
      RECT 17.200000 102.855000 24.540000 102.925000 ;
      RECT 17.200000 102.855000 57.860000 102.925000 ;
      RECT 17.205000 159.390000 60.125000 159.460000 ;
      RECT 17.205000 159.390000 60.125000 159.460000 ;
      RECT 17.220000  67.320000 60.175000  67.390000 ;
      RECT 17.220000  67.320000 60.175000  67.390000 ;
      RECT 17.220000 171.855000 57.870000 171.925000 ;
      RECT 17.225000  56.855000 57.830000  56.925000 ;
      RECT 17.225000 125.785000 24.540000 125.855000 ;
      RECT 17.225000 125.785000 24.540000 125.855000 ;
      RECT 17.225000 125.785000 57.790000 125.855000 ;
      RECT 17.225000 136.460000 60.040000 136.530000 ;
      RECT 17.225000 136.460000 60.040000 136.530000 ;
      RECT 17.225000 148.855000 57.790000 148.925000 ;
      RECT 17.240000  37.235000 54.390000  37.305000 ;
      RECT 17.240000  37.235000 54.390000  37.305000 ;
      RECT 17.250000 182.320000 60.830000 182.390000 ;
      RECT 17.255000  27.660000 57.420000  27.730000 ;
      RECT 17.255000  27.660000 57.420000  27.730000 ;
      RECT 17.255000  90.285000 60.270000  90.355000 ;
      RECT 17.255000  90.285000 60.270000  90.355000 ;
      RECT 17.260000 113.320000 60.145000 113.390000 ;
      RECT 17.260000 113.320000 60.145000 113.390000 ;
      RECT 17.270000  79.925000 24.540000  79.995000 ;
      RECT 17.270000  79.925000 24.540000  79.995000 ;
      RECT 17.270000  79.925000 57.930000  79.995000 ;
      RECT 17.270000 102.925000 24.540000 102.995000 ;
      RECT 17.270000 102.925000 24.540000 102.995000 ;
      RECT 17.270000 102.925000 57.930000 102.995000 ;
      RECT 17.275000 159.320000 60.195000 159.390000 ;
      RECT 17.275000 159.320000 60.195000 159.390000 ;
      RECT 17.290000  67.250000 60.245000  67.320000 ;
      RECT 17.290000  67.250000 60.245000  67.320000 ;
      RECT 17.290000 171.925000 57.940000 171.995000 ;
      RECT 17.295000  56.925000 57.900000  56.995000 ;
      RECT 17.295000 125.855000 24.540000 125.925000 ;
      RECT 17.295000 125.855000 24.540000 125.925000 ;
      RECT 17.295000 125.855000 57.860000 125.925000 ;
      RECT 17.295000 136.390000 60.110000 136.460000 ;
      RECT 17.295000 136.390000 60.110000 136.460000 ;
      RECT 17.295000 148.925000 57.860000 148.995000 ;
      RECT 17.310000  37.305000 54.390000  37.375000 ;
      RECT 17.310000  37.305000 54.390000  37.375000 ;
      RECT 17.320000 182.250000 60.830000 182.320000 ;
      RECT 17.325000  27.590000 57.350000  27.660000 ;
      RECT 17.325000  27.590000 57.350000  27.660000 ;
      RECT 17.325000  90.215000 60.340000  90.285000 ;
      RECT 17.325000  90.215000 60.340000  90.285000 ;
      RECT 17.330000 113.250000 60.215000 113.320000 ;
      RECT 17.330000 113.250000 60.215000 113.320000 ;
      RECT 17.340000  79.995000 24.540000  80.065000 ;
      RECT 17.340000  79.995000 24.540000  80.065000 ;
      RECT 17.340000  79.995000 58.000000  80.065000 ;
      RECT 17.340000 102.995000 24.540000 103.065000 ;
      RECT 17.340000 102.995000 24.540000 103.065000 ;
      RECT 17.340000 102.995000 58.000000 103.065000 ;
      RECT 17.345000 159.250000 60.265000 159.320000 ;
      RECT 17.345000 159.250000 60.265000 159.320000 ;
      RECT 17.360000  67.180000 60.315000  67.250000 ;
      RECT 17.360000  67.180000 60.315000  67.250000 ;
      RECT 17.360000 171.995000 58.010000 172.065000 ;
      RECT 17.365000  56.995000 57.970000  57.065000 ;
      RECT 17.365000 125.925000 24.540000 125.995000 ;
      RECT 17.365000 125.925000 24.540000 125.995000 ;
      RECT 17.365000 125.925000 57.930000 125.995000 ;
      RECT 17.365000 136.320000 60.180000 136.390000 ;
      RECT 17.365000 136.320000 60.180000 136.390000 ;
      RECT 17.365000 148.995000 57.930000 149.065000 ;
      RECT 17.380000  37.375000 54.390000  37.445000 ;
      RECT 17.380000  37.375000 54.390000  37.445000 ;
      RECT 17.390000 182.180000 60.830000 182.250000 ;
      RECT 17.395000  27.520000 57.280000  27.590000 ;
      RECT 17.395000  27.520000 57.280000  27.590000 ;
      RECT 17.395000  90.145000 60.410000  90.215000 ;
      RECT 17.395000  90.145000 60.410000  90.215000 ;
      RECT 17.400000 113.180000 60.285000 113.250000 ;
      RECT 17.400000 113.180000 60.285000 113.250000 ;
      RECT 17.410000  80.065000 24.540000  80.135000 ;
      RECT 17.410000  80.065000 24.540000  80.135000 ;
      RECT 17.410000  80.065000 58.070000  80.135000 ;
      RECT 17.410000 103.065000 24.540000 103.135000 ;
      RECT 17.410000 103.065000 24.540000 103.135000 ;
      RECT 17.410000 103.065000 58.070000 103.135000 ;
      RECT 17.415000 159.180000 60.335000 159.250000 ;
      RECT 17.415000 159.180000 60.335000 159.250000 ;
      RECT 17.430000  67.110000 60.385000  67.180000 ;
      RECT 17.430000  67.110000 60.385000  67.180000 ;
      RECT 17.430000 172.065000 58.080000 172.135000 ;
      RECT 17.435000  57.065000 58.040000  57.135000 ;
      RECT 17.435000 125.995000 24.540000 126.065000 ;
      RECT 17.435000 125.995000 24.540000 126.065000 ;
      RECT 17.435000 125.995000 58.000000 126.065000 ;
      RECT 17.435000 136.250000 60.250000 136.320000 ;
      RECT 17.435000 136.250000 60.250000 136.320000 ;
      RECT 17.435000 149.065000 58.000000 149.135000 ;
      RECT 17.450000  37.445000 54.390000  37.515000 ;
      RECT 17.450000  37.445000 54.390000  37.515000 ;
      RECT 17.460000 182.110000 60.830000 182.180000 ;
      RECT 17.465000  27.450000 57.210000  27.520000 ;
      RECT 17.465000  27.450000 57.210000  27.520000 ;
      RECT 17.465000  90.075000 60.480000  90.145000 ;
      RECT 17.465000  90.075000 60.480000  90.145000 ;
      RECT 17.470000 113.110000 60.355000 113.180000 ;
      RECT 17.470000 113.110000 60.355000 113.180000 ;
      RECT 17.480000  80.135000 24.540000  80.205000 ;
      RECT 17.480000  80.135000 24.540000  80.205000 ;
      RECT 17.480000  80.135000 58.140000  80.205000 ;
      RECT 17.480000 103.135000 24.540000 103.205000 ;
      RECT 17.480000 103.135000 24.540000 103.205000 ;
      RECT 17.480000 103.135000 58.140000 103.205000 ;
      RECT 17.485000 159.110000 60.405000 159.180000 ;
      RECT 17.485000 159.110000 60.405000 159.180000 ;
      RECT 17.500000  67.040000 60.455000  67.110000 ;
      RECT 17.500000  67.040000 60.455000  67.110000 ;
      RECT 17.500000 172.135000 58.150000 172.205000 ;
      RECT 17.505000  57.135000 58.110000  57.205000 ;
      RECT 17.505000 126.065000 24.540000 126.135000 ;
      RECT 17.505000 126.065000 24.540000 126.135000 ;
      RECT 17.505000 126.065000 58.070000 126.135000 ;
      RECT 17.505000 136.180000 60.320000 136.250000 ;
      RECT 17.505000 136.180000 60.320000 136.250000 ;
      RECT 17.505000 149.135000 58.070000 149.205000 ;
      RECT 17.520000  37.515000 54.390000  37.585000 ;
      RECT 17.520000  37.515000 54.390000  37.585000 ;
      RECT 17.530000 182.040000 60.830000 182.110000 ;
      RECT 17.535000  27.380000 57.140000  27.450000 ;
      RECT 17.535000  27.380000 57.140000  27.450000 ;
      RECT 17.535000  90.005000 60.550000  90.075000 ;
      RECT 17.535000  90.005000 60.550000  90.075000 ;
      RECT 17.540000 113.040000 60.425000 113.110000 ;
      RECT 17.540000 113.040000 60.425000 113.110000 ;
      RECT 17.550000  80.205000 24.540000  80.275000 ;
      RECT 17.550000  80.205000 24.540000  80.275000 ;
      RECT 17.550000  80.205000 58.210000  80.275000 ;
      RECT 17.550000 103.205000 24.540000 103.275000 ;
      RECT 17.550000 103.205000 24.540000 103.275000 ;
      RECT 17.550000 103.205000 58.210000 103.275000 ;
      RECT 17.555000 159.040000 60.475000 159.110000 ;
      RECT 17.555000 159.040000 60.475000 159.110000 ;
      RECT 17.570000  66.970000 60.525000  67.040000 ;
      RECT 17.570000  66.970000 60.525000  67.040000 ;
      RECT 17.570000 172.205000 58.220000 172.275000 ;
      RECT 17.575000  57.205000 58.180000  57.275000 ;
      RECT 17.575000 126.135000 24.540000 126.205000 ;
      RECT 17.575000 126.135000 24.540000 126.205000 ;
      RECT 17.575000 126.135000 58.140000 126.205000 ;
      RECT 17.575000 136.110000 60.390000 136.180000 ;
      RECT 17.575000 136.110000 60.390000 136.180000 ;
      RECT 17.575000 149.205000 58.140000 149.275000 ;
      RECT 17.590000  37.585000 54.390000  37.655000 ;
      RECT 17.590000  37.585000 54.390000  37.655000 ;
      RECT 17.600000 181.970000 60.830000 182.040000 ;
      RECT 17.605000  27.310000 57.070000  27.380000 ;
      RECT 17.605000  27.310000 57.070000  27.380000 ;
      RECT 17.605000  89.935000 60.620000  90.005000 ;
      RECT 17.605000  89.935000 60.620000  90.005000 ;
      RECT 17.610000 112.970000 60.495000 113.040000 ;
      RECT 17.610000 112.970000 60.495000 113.040000 ;
      RECT 17.620000  80.275000 24.540000  80.345000 ;
      RECT 17.620000  80.275000 24.540000  80.345000 ;
      RECT 17.620000  80.275000 58.280000  80.345000 ;
      RECT 17.620000 103.275000 24.540000 103.345000 ;
      RECT 17.620000 103.275000 24.540000 103.345000 ;
      RECT 17.620000 103.275000 58.280000 103.345000 ;
      RECT 17.625000 158.970000 60.545000 159.040000 ;
      RECT 17.625000 158.970000 60.545000 159.040000 ;
      RECT 17.640000  66.900000 60.595000  66.970000 ;
      RECT 17.640000  66.900000 60.595000  66.970000 ;
      RECT 17.640000 172.275000 58.290000 172.345000 ;
      RECT 17.645000  57.275000 58.250000  57.345000 ;
      RECT 17.645000 126.205000 24.540000 126.275000 ;
      RECT 17.645000 126.205000 24.540000 126.275000 ;
      RECT 17.645000 126.205000 58.210000 126.275000 ;
      RECT 17.645000 136.040000 60.460000 136.110000 ;
      RECT 17.645000 136.040000 60.460000 136.110000 ;
      RECT 17.645000 149.275000 58.210000 149.345000 ;
      RECT 17.660000  37.655000 54.390000  37.725000 ;
      RECT 17.660000  37.655000 54.390000  37.725000 ;
      RECT 17.670000 181.900000 60.830000 181.970000 ;
      RECT 17.675000  27.240000 57.000000  27.310000 ;
      RECT 17.675000  27.240000 57.000000  27.310000 ;
      RECT 17.675000  89.865000 60.690000  89.935000 ;
      RECT 17.675000  89.865000 60.690000  89.935000 ;
      RECT 17.680000 112.900000 60.565000 112.970000 ;
      RECT 17.680000 112.900000 60.565000 112.970000 ;
      RECT 17.690000  80.345000 24.540000  80.415000 ;
      RECT 17.690000  80.345000 24.540000  80.415000 ;
      RECT 17.690000  80.345000 58.350000  80.415000 ;
      RECT 17.690000  89.850000 57.680000  93.140000 ;
      RECT 17.690000 103.345000 24.540000 103.415000 ;
      RECT 17.690000 103.345000 24.540000 103.415000 ;
      RECT 17.690000 103.345000 58.350000 103.415000 ;
      RECT 17.695000 158.900000 60.615000 158.970000 ;
      RECT 17.695000 158.900000 60.615000 158.970000 ;
      RECT 17.710000  66.830000 60.665000  66.900000 ;
      RECT 17.710000  66.830000 60.665000  66.900000 ;
      RECT 17.710000 172.345000 58.360000 172.415000 ;
      RECT 17.715000  57.345000 58.320000  57.415000 ;
      RECT 17.715000 126.275000 24.540000 126.345000 ;
      RECT 17.715000 126.275000 24.540000 126.345000 ;
      RECT 17.715000 126.275000 58.280000 126.345000 ;
      RECT 17.715000 135.970000 60.530000 136.040000 ;
      RECT 17.715000 135.970000 60.530000 136.040000 ;
      RECT 17.715000 149.345000 58.280000 149.415000 ;
      RECT 17.730000  37.725000 54.390000  37.795000 ;
      RECT 17.730000  37.725000 54.390000  37.795000 ;
      RECT 17.740000 181.830000 60.830000 181.900000 ;
      RECT 17.745000  27.170000 56.930000  27.240000 ;
      RECT 17.745000  27.170000 56.930000  27.240000 ;
      RECT 17.745000  89.795000 60.760000  89.865000 ;
      RECT 17.745000  89.795000 60.760000  89.865000 ;
      RECT 17.750000  66.790000 57.620000  70.140000 ;
      RECT 17.750000  89.790000 60.830000  89.795000 ;
      RECT 17.750000  89.790000 60.830000  89.795000 ;
      RECT 17.750000 112.830000 60.635000 112.900000 ;
      RECT 17.750000 112.830000 60.635000 112.900000 ;
      RECT 17.760000  80.415000 24.540000  80.485000 ;
      RECT 17.760000  80.415000 24.540000  80.485000 ;
      RECT 17.760000  80.415000 58.420000  80.485000 ;
      RECT 17.760000 103.415000 24.540000 103.485000 ;
      RECT 17.760000 103.415000 24.540000 103.485000 ;
      RECT 17.760000 103.415000 58.420000 103.485000 ;
      RECT 17.765000  89.775000 60.830000  89.790000 ;
      RECT 17.765000  89.775000 60.830000  89.790000 ;
      RECT 17.765000 158.830000 60.685000 158.900000 ;
      RECT 17.765000 158.830000 60.685000 158.900000 ;
      RECT 17.775000  80.485000 24.540000  80.500000 ;
      RECT 17.775000  80.485000 24.540000  80.500000 ;
      RECT 17.775000  80.485000 58.490000  80.500000 ;
      RECT 17.775000 103.485000 24.540000 103.500000 ;
      RECT 17.775000 103.485000 24.540000 103.500000 ;
      RECT 17.775000 103.485000 58.490000 103.500000 ;
      RECT 17.780000  66.760000 60.735000  66.830000 ;
      RECT 17.780000  66.760000 60.735000  66.830000 ;
      RECT 17.780000  66.760000 60.970000  66.790000 ;
      RECT 17.780000  89.760000 60.830000  89.775000 ;
      RECT 17.780000  89.760000 60.830000  89.775000 ;
      RECT 17.780000  89.760000 60.970000  89.850000 ;
      RECT 17.780000 172.415000 58.430000 172.485000 ;
      RECT 17.785000  57.415000 58.390000  57.485000 ;
      RECT 17.785000 126.345000 24.540000 126.415000 ;
      RECT 17.785000 126.345000 24.540000 126.415000 ;
      RECT 17.785000 126.345000 58.350000 126.415000 ;
      RECT 17.785000 135.900000 60.600000 135.970000 ;
      RECT 17.785000 135.900000 60.600000 135.970000 ;
      RECT 17.785000 149.415000 58.350000 149.485000 ;
      RECT 17.785000 158.810000 57.585000 162.195000 ;
      RECT 17.795000 172.485000 58.500000 172.500000 ;
      RECT 17.800000  37.795000 54.390000  37.865000 ;
      RECT 17.800000  37.795000 54.390000  37.865000 ;
      RECT 17.800000  57.485000 58.460000  57.500000 ;
      RECT 17.800000 149.485000 58.420000 149.500000 ;
      RECT 17.810000 181.760000 60.830000 181.830000 ;
      RECT 17.810000 181.760000 60.970000 182.820000 ;
      RECT 17.815000  27.100000 56.860000  27.170000 ;
      RECT 17.815000  27.100000 56.860000  27.170000 ;
      RECT 17.820000 112.760000 57.550000 116.180000 ;
      RECT 17.820000 112.760000 60.705000 112.830000 ;
      RECT 17.820000 112.760000 60.705000 112.830000 ;
      RECT 17.820000 112.760000 60.970000 112.760000 ;
      RECT 17.835000 158.760000 60.755000 158.830000 ;
      RECT 17.835000 158.760000 60.755000 158.830000 ;
      RECT 17.835000 158.760000 60.970000 158.810000 ;
      RECT 17.855000 126.415000 24.540000 126.485000 ;
      RECT 17.855000 126.415000 24.540000 126.485000 ;
      RECT 17.855000 126.415000 58.420000 126.485000 ;
      RECT 17.855000 135.830000 60.670000 135.900000 ;
      RECT 17.855000 135.830000 60.670000 135.900000 ;
      RECT 17.870000  37.865000 54.390000  37.935000 ;
      RECT 17.870000  37.865000 54.390000  37.935000 ;
      RECT 17.870000 126.485000 24.540000 126.500000 ;
      RECT 17.870000 126.485000 24.540000 126.500000 ;
      RECT 17.870000 126.485000 58.490000 126.500000 ;
      RECT 17.885000  27.030000 56.790000  27.100000 ;
      RECT 17.885000  27.030000 56.790000  27.100000 ;
      RECT 17.890000 135.795000 57.480000 139.285000 ;
      RECT 17.925000 135.760000 60.740000 135.830000 ;
      RECT 17.925000 135.760000 60.740000 135.830000 ;
      RECT 17.925000 135.760000 60.970000 135.795000 ;
      RECT 17.940000  37.935000 54.390000  38.005000 ;
      RECT 17.940000  37.935000 54.390000  38.005000 ;
      RECT 17.955000  26.960000 56.720000  27.030000 ;
      RECT 17.955000  26.960000 56.720000  27.030000 ;
      RECT 18.010000  38.005000 54.390000  38.075000 ;
      RECT 18.010000  38.005000 54.390000  38.075000 ;
      RECT 18.025000  26.890000 56.650000  26.960000 ;
      RECT 18.025000  26.890000 56.650000  26.960000 ;
      RECT 18.075000  38.075000 54.390000  38.140000 ;
      RECT 18.075000  38.075000 54.390000  38.140000 ;
      RECT 18.095000  26.820000 56.580000  26.890000 ;
      RECT 18.095000  26.820000 56.580000  26.890000 ;
      RECT 18.130000  38.195000 52.655000  40.070000 ;
      RECT 18.145000  38.140000 54.320000  38.210000 ;
      RECT 18.145000  38.140000 54.320000  38.210000 ;
      RECT 18.165000  26.750000 56.510000  26.820000 ;
      RECT 18.165000  26.750000 56.510000  26.820000 ;
      RECT 18.215000  38.210000 54.250000  38.280000 ;
      RECT 18.215000  38.210000 54.250000  38.280000 ;
      RECT 18.235000  26.680000 56.440000  26.750000 ;
      RECT 18.235000  26.680000 56.440000  26.750000 ;
      RECT 18.285000  38.280000 54.180000  38.350000 ;
      RECT 18.285000  38.280000 54.180000  38.350000 ;
      RECT 18.305000  26.610000 56.370000  26.680000 ;
      RECT 18.305000  26.610000 56.370000  26.680000 ;
      RECT 18.355000  38.350000 54.110000  38.420000 ;
      RECT 18.355000  38.350000 54.110000  38.420000 ;
      RECT 18.375000  26.540000 56.300000  26.610000 ;
      RECT 18.375000  26.540000 56.300000  26.610000 ;
      RECT 18.425000  38.420000 54.040000  38.490000 ;
      RECT 18.425000  38.420000 54.040000  38.490000 ;
      RECT 18.445000  26.470000 56.230000  26.540000 ;
      RECT 18.445000  26.470000 56.230000  26.540000 ;
      RECT 18.495000  38.490000 53.970000  38.560000 ;
      RECT 18.495000  38.490000 53.970000  38.560000 ;
      RECT 18.515000  26.400000 56.160000  26.470000 ;
      RECT 18.515000  26.400000 56.160000  26.470000 ;
      RECT 18.565000  38.560000 53.900000  38.630000 ;
      RECT 18.565000  38.560000 53.900000  38.630000 ;
      RECT 18.585000  26.330000 56.090000  26.400000 ;
      RECT 18.585000  26.330000 56.090000  26.400000 ;
      RECT 18.635000  38.630000 53.830000  38.700000 ;
      RECT 18.635000  38.630000 53.830000  38.700000 ;
      RECT 18.655000  26.260000 56.020000  26.330000 ;
      RECT 18.655000  26.260000 56.020000  26.330000 ;
      RECT 18.705000  38.700000 53.760000  38.770000 ;
      RECT 18.705000  38.700000 53.760000  38.770000 ;
      RECT 18.725000  26.190000 55.950000  26.260000 ;
      RECT 18.725000  26.190000 55.950000  26.260000 ;
      RECT 18.775000  38.770000 53.690000  38.840000 ;
      RECT 18.775000  38.770000 53.690000  38.840000 ;
      RECT 18.795000  26.120000 55.880000  26.190000 ;
      RECT 18.795000  26.120000 55.880000  26.190000 ;
      RECT 18.845000  38.840000 53.620000  38.910000 ;
      RECT 18.845000  38.840000 53.620000  38.910000 ;
      RECT 18.865000  26.050000 55.810000  26.120000 ;
      RECT 18.865000  26.050000 55.810000  26.120000 ;
      RECT 18.915000  38.910000 53.550000  38.980000 ;
      RECT 18.915000  38.910000 53.550000  38.980000 ;
      RECT 18.935000  25.980000 55.740000  26.050000 ;
      RECT 18.935000  25.980000 55.740000  26.050000 ;
      RECT 18.935000  25.980000 59.390000  29.430000 ;
      RECT 18.985000  38.980000 53.480000  39.050000 ;
      RECT 18.985000  38.980000 53.480000  39.050000 ;
      RECT 19.055000  39.050000 53.410000  39.120000 ;
      RECT 19.055000  39.050000 53.410000  39.120000 ;
      RECT 19.125000  39.120000 53.340000  39.190000 ;
      RECT 19.125000  39.120000 53.340000  39.190000 ;
      RECT 19.195000  39.190000 53.270000  39.260000 ;
      RECT 19.195000  39.190000 53.270000  39.260000 ;
      RECT 19.265000  39.260000 53.200000  39.330000 ;
      RECT 19.265000  39.260000 53.200000  39.330000 ;
      RECT 19.335000  39.330000 53.130000  39.400000 ;
      RECT 19.335000  39.330000 53.130000  39.400000 ;
      RECT 19.405000  39.400000 53.060000  39.470000 ;
      RECT 19.405000  39.400000 53.060000  39.470000 ;
      RECT 19.475000  39.470000 52.990000  39.540000 ;
      RECT 19.475000  39.470000 52.990000  39.540000 ;
      RECT 19.545000  39.540000 52.920000  39.610000 ;
      RECT 19.545000  39.540000 52.920000  39.610000 ;
      RECT 19.615000  39.610000 52.850000  39.680000 ;
      RECT 19.615000  39.610000 52.850000  39.680000 ;
      RECT 19.685000  39.680000 52.780000  39.750000 ;
      RECT 19.685000  39.680000 52.780000  39.750000 ;
      RECT 19.755000  39.750000 52.710000  39.820000 ;
      RECT 19.755000  39.750000 52.710000  39.820000 ;
      RECT 19.825000  39.820000 52.640000  39.890000 ;
      RECT 19.825000  39.820000 52.640000  39.890000 ;
      RECT 19.895000  39.890000 52.570000  39.960000 ;
      RECT 19.895000  39.890000 52.570000  39.960000 ;
      RECT 19.965000  39.960000 52.500000  40.030000 ;
      RECT 19.965000  39.960000 52.500000  40.030000 ;
      RECT 20.005000  40.030000 52.460000  40.070000 ;
      RECT 20.005000  40.030000 52.460000  40.070000 ;
      RECT 20.400000  40.070000 52.515000  40.210000 ;
      RECT 22.850000  42.520000 60.970000  42.660000 ;
      RECT 24.675000   0.000000 25.615000   0.815000 ;
      RECT 24.675000   0.000000 25.755000   0.675000 ;
      RECT 24.675000   0.675000 50.250000   8.480000 ;
      RECT 24.675000   0.815000 50.110000   8.480000 ;
      RECT 24.675000   8.480000 50.250000   8.565000 ;
      RECT 24.690000   8.480000 50.110000   8.495000 ;
      RECT 24.690000   8.480000 50.110000   8.495000 ;
      RECT 24.705000   8.495000 50.110000   8.510000 ;
      RECT 24.705000   8.495000 50.110000   8.510000 ;
      RECT 24.765000   8.565000 46.695000  12.120000 ;
      RECT 24.775000   8.510000 50.040000   8.580000 ;
      RECT 24.775000   8.510000 50.040000   8.580000 ;
      RECT 24.845000   8.580000 49.970000   8.650000 ;
      RECT 24.845000   8.580000 49.970000   8.650000 ;
      RECT 24.915000   8.650000 49.900000   8.720000 ;
      RECT 24.915000   8.650000 49.900000   8.720000 ;
      RECT 24.985000   8.720000 49.830000   8.790000 ;
      RECT 24.985000   8.720000 49.830000   8.790000 ;
      RECT 25.055000   8.790000 49.760000   8.860000 ;
      RECT 25.055000   8.790000 49.760000   8.860000 ;
      RECT 25.125000   8.860000 49.690000   8.930000 ;
      RECT 25.125000   8.860000 49.690000   8.930000 ;
      RECT 25.195000   8.930000 49.620000   9.000000 ;
      RECT 25.195000   8.930000 49.620000   9.000000 ;
      RECT 25.265000   9.000000 49.550000   9.070000 ;
      RECT 25.265000   9.000000 49.550000   9.070000 ;
      RECT 25.335000   9.070000 49.480000   9.140000 ;
      RECT 25.335000   9.070000 49.480000   9.140000 ;
      RECT 25.405000   9.140000 49.410000   9.210000 ;
      RECT 25.405000   9.140000 49.410000   9.210000 ;
      RECT 25.475000   9.210000 49.340000   9.280000 ;
      RECT 25.475000   9.210000 49.340000   9.280000 ;
      RECT 25.545000   9.280000 49.270000   9.350000 ;
      RECT 25.545000   9.280000 49.270000   9.350000 ;
      RECT 25.615000   9.350000 49.200000   9.420000 ;
      RECT 25.615000   9.350000 49.200000   9.420000 ;
      RECT 25.685000   9.420000 49.130000   9.490000 ;
      RECT 25.685000   9.420000 49.130000   9.490000 ;
      RECT 25.755000   9.490000 49.060000   9.560000 ;
      RECT 25.755000   9.490000 49.060000   9.560000 ;
      RECT 25.825000   9.560000 48.990000   9.630000 ;
      RECT 25.825000   9.560000 48.990000   9.630000 ;
      RECT 25.895000   9.630000 48.920000   9.700000 ;
      RECT 25.895000   9.630000 48.920000   9.700000 ;
      RECT 25.965000   9.700000 48.850000   9.770000 ;
      RECT 25.965000   9.700000 48.850000   9.770000 ;
      RECT 26.035000   9.770000 48.780000   9.840000 ;
      RECT 26.035000   9.770000 48.780000   9.840000 ;
      RECT 26.105000   9.840000 48.710000   9.910000 ;
      RECT 26.105000   9.840000 48.710000   9.910000 ;
      RECT 26.175000   9.910000 48.640000   9.980000 ;
      RECT 26.175000   9.910000 48.640000   9.980000 ;
      RECT 26.245000   9.980000 48.570000  10.050000 ;
      RECT 26.245000   9.980000 48.570000  10.050000 ;
      RECT 26.315000  10.050000 48.500000  10.120000 ;
      RECT 26.315000  10.050000 48.500000  10.120000 ;
      RECT 26.385000  10.120000 48.430000  10.190000 ;
      RECT 26.385000  10.120000 48.430000  10.190000 ;
      RECT 26.455000  10.190000 48.360000  10.260000 ;
      RECT 26.455000  10.190000 48.360000  10.260000 ;
      RECT 26.525000  10.260000 48.290000  10.330000 ;
      RECT 26.525000  10.260000 48.290000  10.330000 ;
      RECT 26.595000  10.330000 48.220000  10.400000 ;
      RECT 26.595000  10.330000 48.220000  10.400000 ;
      RECT 26.665000  10.400000 48.150000  10.470000 ;
      RECT 26.665000  10.400000 48.150000  10.470000 ;
      RECT 26.735000  10.470000 48.080000  10.540000 ;
      RECT 26.735000  10.470000 48.080000  10.540000 ;
      RECT 26.805000  10.540000 48.010000  10.610000 ;
      RECT 26.805000  10.540000 48.010000  10.610000 ;
      RECT 26.875000  10.610000 47.940000  10.680000 ;
      RECT 26.875000  10.610000 47.940000  10.680000 ;
      RECT 26.945000  10.680000 47.870000  10.750000 ;
      RECT 26.945000  10.680000 47.870000  10.750000 ;
      RECT 27.015000  10.750000 47.800000  10.820000 ;
      RECT 27.015000  10.750000 47.800000  10.820000 ;
      RECT 27.085000  10.820000 47.730000  10.890000 ;
      RECT 27.085000  10.820000 47.730000  10.890000 ;
      RECT 27.155000  10.890000 47.660000  10.960000 ;
      RECT 27.155000  10.890000 47.660000  10.960000 ;
      RECT 27.225000  10.960000 47.590000  11.030000 ;
      RECT 27.225000  10.960000 47.590000  11.030000 ;
      RECT 27.295000  11.030000 47.520000  11.100000 ;
      RECT 27.295000  11.030000 47.520000  11.100000 ;
      RECT 27.365000  11.100000 47.450000  11.170000 ;
      RECT 27.365000  11.100000 47.450000  11.170000 ;
      RECT 27.435000  11.170000 47.380000  11.240000 ;
      RECT 27.435000  11.170000 47.380000  11.240000 ;
      RECT 27.505000  11.240000 47.310000  11.310000 ;
      RECT 27.505000  11.240000 47.310000  11.310000 ;
      RECT 27.575000  11.310000 47.240000  11.380000 ;
      RECT 27.575000  11.310000 47.240000  11.380000 ;
      RECT 27.645000  11.380000 47.170000  11.450000 ;
      RECT 27.645000  11.380000 47.170000  11.450000 ;
      RECT 27.715000  11.450000 47.100000  11.520000 ;
      RECT 27.715000  11.450000 47.100000  11.520000 ;
      RECT 27.785000  11.520000 47.030000  11.590000 ;
      RECT 27.785000  11.520000 47.030000  11.590000 ;
      RECT 27.855000  11.590000 46.960000  11.660000 ;
      RECT 27.855000  11.590000 46.960000  11.660000 ;
      RECT 27.925000  11.660000 46.890000  11.730000 ;
      RECT 27.925000  11.660000 46.890000  11.730000 ;
      RECT 27.995000  11.730000 46.820000  11.800000 ;
      RECT 27.995000  11.730000 46.820000  11.800000 ;
      RECT 28.035000   0.000000 50.250000   0.675000 ;
      RECT 28.065000  11.800000 46.750000  11.870000 ;
      RECT 28.065000  11.800000 46.750000  11.870000 ;
      RECT 28.135000  11.870000 46.680000  11.940000 ;
      RECT 28.135000  11.870000 46.680000  11.940000 ;
      RECT 28.175000   0.000000 50.110000   0.815000 ;
      RECT 28.175000   0.000000 50.110000   8.480000 ;
      RECT 28.205000  11.940000 46.610000  12.010000 ;
      RECT 28.205000  11.940000 46.610000  12.010000 ;
      RECT 28.210000  12.010000 46.605000  12.015000 ;
      RECT 28.210000  12.010000 46.605000  12.015000 ;
      RECT 28.260000  12.015000 37.610000  12.065000 ;
      RECT 28.260000  12.015000 37.610000  12.065000 ;
      RECT 28.310000  12.065000 37.610000  12.115000 ;
      RECT 28.310000  12.065000 37.610000  12.115000 ;
      RECT 28.315000  12.115000 37.610000  12.120000 ;
      RECT 28.315000  12.115000 37.610000  12.120000 ;
      RECT 37.175000  12.120000 37.610000  25.940000 ;
      RECT 37.175000  12.120000 46.660000  12.155000 ;
      RECT 37.175000  12.155000 37.750000  25.800000 ;
      RECT 37.175000  25.800000 55.935000  25.980000 ;
      RECT 37.175000  25.940000 55.700000  25.960000 ;
      RECT 37.175000  25.940000 55.700000  25.960000 ;
      RECT 37.175000  25.960000 55.720000  25.980000 ;
      RECT 37.175000  25.960000 55.720000  25.980000 ;
      RECT 54.325000  42.650000 60.830000  42.660000 ;
      RECT 54.325000  42.650000 60.830000  42.660000 ;
      RECT 54.395000  42.580000 60.830000  42.650000 ;
      RECT 54.395000  42.580000 60.830000  42.650000 ;
      RECT 54.465000  42.510000 60.830000  42.580000 ;
      RECT 54.465000  42.510000 60.830000  42.580000 ;
      RECT 54.535000  42.440000 60.830000  42.510000 ;
      RECT 54.535000  42.440000 60.830000  42.510000 ;
      RECT 54.605000  42.370000 60.830000  42.440000 ;
      RECT 54.605000  42.370000 60.830000  42.440000 ;
      RECT 54.675000  42.300000 60.830000  42.370000 ;
      RECT 54.675000  42.300000 60.830000  42.370000 ;
      RECT 54.745000  42.230000 60.830000  42.300000 ;
      RECT 54.745000  42.230000 60.830000  42.300000 ;
      RECT 54.815000  42.160000 60.830000  42.230000 ;
      RECT 54.815000  42.160000 60.830000  42.230000 ;
      RECT 54.885000  42.090000 60.830000  42.160000 ;
      RECT 54.885000  42.090000 60.830000  42.160000 ;
      RECT 54.955000  42.020000 60.830000  42.090000 ;
      RECT 54.955000  42.020000 60.830000  42.090000 ;
      RECT 55.025000  41.950000 60.830000  42.020000 ;
      RECT 55.025000  41.950000 60.830000  42.020000 ;
      RECT 55.095000  41.880000 60.830000  41.950000 ;
      RECT 55.095000  41.880000 60.830000  41.950000 ;
      RECT 55.165000  41.810000 60.830000  41.880000 ;
      RECT 55.165000  41.810000 60.830000  41.880000 ;
      RECT 55.235000  41.740000 60.830000  41.810000 ;
      RECT 55.235000  41.740000 60.830000  41.810000 ;
      RECT 55.305000  41.670000 60.830000  41.740000 ;
      RECT 55.305000  41.670000 60.830000  41.740000 ;
      RECT 55.375000  41.600000 60.830000  41.670000 ;
      RECT 55.375000  41.600000 60.830000  41.670000 ;
      RECT 55.445000  41.530000 60.830000  41.600000 ;
      RECT 55.445000  41.530000 60.830000  41.600000 ;
      RECT 55.515000  41.460000 60.830000  41.530000 ;
      RECT 55.515000  41.460000 60.830000  41.530000 ;
      RECT 55.585000  41.390000 60.830000  41.460000 ;
      RECT 55.585000  41.390000 60.830000  41.460000 ;
      RECT 55.655000  41.320000 60.830000  41.390000 ;
      RECT 55.655000  41.320000 60.830000  41.390000 ;
      RECT 55.725000  41.250000 60.830000  41.320000 ;
      RECT 55.725000  41.250000 60.830000  41.320000 ;
      RECT 55.795000  41.180000 60.830000  41.250000 ;
      RECT 55.795000  41.180000 60.830000  41.250000 ;
      RECT 55.865000  41.110000 60.830000  41.180000 ;
      RECT 55.865000  41.110000 60.830000  41.180000 ;
      RECT 55.935000  41.040000 60.830000  41.110000 ;
      RECT 55.935000  41.040000 60.830000  41.110000 ;
      RECT 56.005000  40.970000 60.830000  41.040000 ;
      RECT 56.005000  40.970000 60.830000  41.040000 ;
      RECT 56.075000  40.900000 60.830000  40.970000 ;
      RECT 56.075000  40.900000 60.830000  40.970000 ;
      RECT 56.145000  40.830000 60.830000  40.900000 ;
      RECT 56.145000  40.830000 60.830000  40.900000 ;
      RECT 56.215000  40.760000 60.830000  40.830000 ;
      RECT 56.215000  40.760000 60.830000  40.830000 ;
      RECT 56.285000  40.690000 60.830000  40.760000 ;
      RECT 56.285000  40.690000 60.830000  40.760000 ;
      RECT 56.355000  40.620000 60.830000  40.690000 ;
      RECT 56.355000  40.620000 60.830000  40.690000 ;
      RECT 56.425000  40.550000 60.830000  40.620000 ;
      RECT 56.425000  40.550000 60.830000  40.620000 ;
      RECT 56.495000  40.480000 60.830000  40.550000 ;
      RECT 56.495000  40.480000 60.830000  40.550000 ;
      RECT 56.565000  40.410000 60.830000  40.480000 ;
      RECT 56.565000  40.410000 60.830000  40.480000 ;
      RECT 56.635000  40.340000 60.830000  40.410000 ;
      RECT 56.635000  40.340000 60.830000  40.410000 ;
      RECT 56.705000  40.270000 60.830000  40.340000 ;
      RECT 56.705000  40.270000 60.830000  40.340000 ;
      RECT 56.775000  40.200000 60.830000  40.270000 ;
      RECT 56.775000  40.200000 60.830000  40.270000 ;
      RECT 56.845000  40.130000 60.830000  40.200000 ;
      RECT 56.845000  40.130000 60.830000  40.200000 ;
      RECT 56.915000  40.060000 60.830000  40.130000 ;
      RECT 56.915000  40.060000 60.830000  40.130000 ;
      RECT 56.985000  39.990000 60.830000  40.060000 ;
      RECT 56.985000  39.990000 60.830000  40.060000 ;
      RECT 56.985000  79.435000 57.440000  79.505000 ;
      RECT 56.985000  79.435000 57.440000  79.505000 ;
      RECT 56.985000  79.505000 57.510000  79.575000 ;
      RECT 56.985000  79.505000 57.510000  79.575000 ;
      RECT 56.985000  79.575000 57.580000  79.645000 ;
      RECT 56.985000  79.575000 57.580000  79.645000 ;
      RECT 56.985000  79.645000 57.650000  79.715000 ;
      RECT 56.985000  79.645000 57.650000  79.715000 ;
      RECT 56.985000  79.715000 57.720000  79.785000 ;
      RECT 56.985000  79.715000 57.720000  79.785000 ;
      RECT 56.985000  79.785000 57.790000  79.855000 ;
      RECT 56.985000  79.785000 57.790000  79.855000 ;
      RECT 56.985000  79.855000 57.860000  79.925000 ;
      RECT 56.985000  79.855000 57.860000  79.925000 ;
      RECT 56.985000  79.925000 57.930000  79.995000 ;
      RECT 56.985000  79.925000 57.930000  79.995000 ;
      RECT 56.985000  79.995000 58.000000  80.065000 ;
      RECT 56.985000  79.995000 58.000000  80.065000 ;
      RECT 56.985000  80.065000 58.070000  80.135000 ;
      RECT 56.985000  80.065000 58.070000  80.135000 ;
      RECT 56.985000  80.135000 58.140000  80.205000 ;
      RECT 56.985000  80.135000 58.140000  80.205000 ;
      RECT 56.985000  80.205000 58.210000  80.275000 ;
      RECT 56.985000  80.205000 58.210000  80.275000 ;
      RECT 56.985000  80.275000 58.280000  80.345000 ;
      RECT 56.985000  80.275000 58.280000  80.345000 ;
      RECT 56.985000  80.345000 58.350000  80.415000 ;
      RECT 56.985000  80.345000 58.350000  80.415000 ;
      RECT 56.985000  80.415000 58.420000  80.485000 ;
      RECT 56.985000  80.415000 58.420000  80.485000 ;
      RECT 56.985000  80.485000 58.490000  80.500000 ;
      RECT 56.985000  80.485000 58.490000  80.500000 ;
      RECT 56.985000  80.500000 58.505000  80.570000 ;
      RECT 56.985000  80.500000 58.505000  80.570000 ;
      RECT 56.985000  80.500000 60.970000  82.770000 ;
      RECT 56.985000  80.570000 58.575000  80.640000 ;
      RECT 56.985000  80.570000 58.575000  80.640000 ;
      RECT 56.985000  80.640000 58.645000  80.710000 ;
      RECT 56.985000  80.640000 58.645000  80.710000 ;
      RECT 56.985000  80.710000 58.715000  80.780000 ;
      RECT 56.985000  80.710000 58.715000  80.780000 ;
      RECT 56.985000  80.780000 58.785000  80.850000 ;
      RECT 56.985000  80.780000 58.785000  80.850000 ;
      RECT 56.985000  80.850000 58.855000  80.920000 ;
      RECT 56.985000  80.850000 58.855000  80.920000 ;
      RECT 56.985000  80.920000 58.925000  80.990000 ;
      RECT 56.985000  80.920000 58.925000  80.990000 ;
      RECT 56.985000  80.990000 58.995000  81.060000 ;
      RECT 56.985000  80.990000 58.995000  81.060000 ;
      RECT 56.985000  81.060000 59.065000  81.130000 ;
      RECT 56.985000  81.060000 59.065000  81.130000 ;
      RECT 56.985000  81.130000 59.135000  81.200000 ;
      RECT 56.985000  81.130000 59.135000  81.200000 ;
      RECT 56.985000  81.200000 59.205000  81.270000 ;
      RECT 56.985000  81.200000 59.205000  81.270000 ;
      RECT 56.985000  81.270000 59.275000  81.340000 ;
      RECT 56.985000  81.270000 59.275000  81.340000 ;
      RECT 56.985000  81.340000 59.345000  81.410000 ;
      RECT 56.985000  81.340000 59.345000  81.410000 ;
      RECT 56.985000  81.410000 59.415000  81.480000 ;
      RECT 56.985000  81.410000 59.415000  81.480000 ;
      RECT 56.985000  81.480000 59.485000  81.550000 ;
      RECT 56.985000  81.480000 59.485000  81.550000 ;
      RECT 56.985000  81.550000 59.555000  81.620000 ;
      RECT 56.985000  81.550000 59.555000  81.620000 ;
      RECT 56.985000  81.620000 59.625000  81.690000 ;
      RECT 56.985000  81.620000 59.625000  81.690000 ;
      RECT 56.985000  81.690000 59.695000  81.760000 ;
      RECT 56.985000  81.690000 59.695000  81.760000 ;
      RECT 56.985000  81.760000 59.765000  81.830000 ;
      RECT 56.985000  81.760000 59.765000  81.830000 ;
      RECT 56.985000  81.830000 59.835000  81.900000 ;
      RECT 56.985000  81.830000 59.835000  81.900000 ;
      RECT 56.985000  81.900000 59.905000  81.970000 ;
      RECT 56.985000  81.900000 59.905000  81.970000 ;
      RECT 56.985000  81.970000 59.975000  82.040000 ;
      RECT 56.985000  81.970000 59.975000  82.040000 ;
      RECT 56.985000  82.040000 60.045000  82.110000 ;
      RECT 56.985000  82.040000 60.045000  82.110000 ;
      RECT 56.985000  82.110000 60.115000  82.180000 ;
      RECT 56.985000  82.110000 60.115000  82.180000 ;
      RECT 56.985000  82.180000 60.185000  82.250000 ;
      RECT 56.985000  82.180000 60.185000  82.250000 ;
      RECT 56.985000  82.250000 60.255000  82.320000 ;
      RECT 56.985000  82.250000 60.255000  82.320000 ;
      RECT 56.985000  82.320000 60.325000  82.390000 ;
      RECT 56.985000  82.320000 60.325000  82.390000 ;
      RECT 56.985000  82.390000 60.395000  82.460000 ;
      RECT 56.985000  82.390000 60.395000  82.460000 ;
      RECT 56.985000  82.460000 60.465000  82.530000 ;
      RECT 56.985000  82.460000 60.465000  82.530000 ;
      RECT 56.985000  82.530000 60.535000  82.600000 ;
      RECT 56.985000  82.530000 60.535000  82.600000 ;
      RECT 56.985000  82.600000 60.605000  82.670000 ;
      RECT 56.985000  82.600000 60.605000  82.670000 ;
      RECT 56.985000  82.670000 60.675000  82.740000 ;
      RECT 56.985000  82.670000 60.675000  82.740000 ;
      RECT 56.985000  82.740000 60.745000  82.810000 ;
      RECT 56.985000  82.740000 60.745000  82.810000 ;
      RECT 56.985000  82.770000 60.970000  89.760000 ;
      RECT 56.985000  82.810000 60.815000  82.825000 ;
      RECT 56.985000  82.810000 60.815000  82.825000 ;
      RECT 56.985000  82.825000 60.830000  89.760000 ;
      RECT 56.985000 102.435000 57.440000 102.505000 ;
      RECT 56.985000 102.435000 57.440000 102.505000 ;
      RECT 56.985000 102.505000 57.510000 102.575000 ;
      RECT 56.985000 102.505000 57.510000 102.575000 ;
      RECT 56.985000 102.575000 57.580000 102.645000 ;
      RECT 56.985000 102.575000 57.580000 102.645000 ;
      RECT 56.985000 102.645000 57.650000 102.715000 ;
      RECT 56.985000 102.645000 57.650000 102.715000 ;
      RECT 56.985000 102.715000 57.720000 102.785000 ;
      RECT 56.985000 102.715000 57.720000 102.785000 ;
      RECT 56.985000 102.785000 57.790000 102.855000 ;
      RECT 56.985000 102.785000 57.790000 102.855000 ;
      RECT 56.985000 102.855000 57.860000 102.925000 ;
      RECT 56.985000 102.855000 57.860000 102.925000 ;
      RECT 56.985000 102.925000 57.930000 102.995000 ;
      RECT 56.985000 102.925000 57.930000 102.995000 ;
      RECT 56.985000 102.995000 58.000000 103.065000 ;
      RECT 56.985000 102.995000 58.000000 103.065000 ;
      RECT 56.985000 103.065000 58.070000 103.135000 ;
      RECT 56.985000 103.065000 58.070000 103.135000 ;
      RECT 56.985000 103.135000 58.140000 103.205000 ;
      RECT 56.985000 103.135000 58.140000 103.205000 ;
      RECT 56.985000 103.205000 58.210000 103.275000 ;
      RECT 56.985000 103.205000 58.210000 103.275000 ;
      RECT 56.985000 103.275000 58.280000 103.345000 ;
      RECT 56.985000 103.275000 58.280000 103.345000 ;
      RECT 56.985000 103.345000 58.350000 103.415000 ;
      RECT 56.985000 103.345000 58.350000 103.415000 ;
      RECT 56.985000 103.415000 58.420000 103.485000 ;
      RECT 56.985000 103.415000 58.420000 103.485000 ;
      RECT 56.985000 103.485000 58.490000 103.500000 ;
      RECT 56.985000 103.485000 58.490000 103.500000 ;
      RECT 56.985000 103.500000 58.505000 103.570000 ;
      RECT 56.985000 103.500000 58.505000 103.570000 ;
      RECT 56.985000 103.500000 60.970000 105.770000 ;
      RECT 56.985000 103.570000 58.575000 103.640000 ;
      RECT 56.985000 103.570000 58.575000 103.640000 ;
      RECT 56.985000 103.640000 58.645000 103.710000 ;
      RECT 56.985000 103.640000 58.645000 103.710000 ;
      RECT 56.985000 103.710000 58.715000 103.780000 ;
      RECT 56.985000 103.710000 58.715000 103.780000 ;
      RECT 56.985000 103.780000 58.785000 103.850000 ;
      RECT 56.985000 103.780000 58.785000 103.850000 ;
      RECT 56.985000 103.850000 58.855000 103.920000 ;
      RECT 56.985000 103.850000 58.855000 103.920000 ;
      RECT 56.985000 103.920000 58.925000 103.990000 ;
      RECT 56.985000 103.920000 58.925000 103.990000 ;
      RECT 56.985000 103.990000 58.995000 104.060000 ;
      RECT 56.985000 103.990000 58.995000 104.060000 ;
      RECT 56.985000 104.060000 59.065000 104.130000 ;
      RECT 56.985000 104.060000 59.065000 104.130000 ;
      RECT 56.985000 104.130000 59.135000 104.200000 ;
      RECT 56.985000 104.130000 59.135000 104.200000 ;
      RECT 56.985000 104.200000 59.205000 104.270000 ;
      RECT 56.985000 104.200000 59.205000 104.270000 ;
      RECT 56.985000 104.270000 59.275000 104.340000 ;
      RECT 56.985000 104.270000 59.275000 104.340000 ;
      RECT 56.985000 104.340000 59.345000 104.410000 ;
      RECT 56.985000 104.340000 59.345000 104.410000 ;
      RECT 56.985000 104.410000 59.415000 104.480000 ;
      RECT 56.985000 104.410000 59.415000 104.480000 ;
      RECT 56.985000 104.480000 59.485000 104.550000 ;
      RECT 56.985000 104.480000 59.485000 104.550000 ;
      RECT 56.985000 104.550000 59.555000 104.620000 ;
      RECT 56.985000 104.550000 59.555000 104.620000 ;
      RECT 56.985000 104.620000 59.625000 104.690000 ;
      RECT 56.985000 104.620000 59.625000 104.690000 ;
      RECT 56.985000 104.690000 59.695000 104.760000 ;
      RECT 56.985000 104.690000 59.695000 104.760000 ;
      RECT 56.985000 104.760000 59.765000 104.830000 ;
      RECT 56.985000 104.760000 59.765000 104.830000 ;
      RECT 56.985000 104.830000 59.835000 104.900000 ;
      RECT 56.985000 104.830000 59.835000 104.900000 ;
      RECT 56.985000 104.900000 59.905000 104.970000 ;
      RECT 56.985000 104.900000 59.905000 104.970000 ;
      RECT 56.985000 104.970000 59.975000 105.040000 ;
      RECT 56.985000 104.970000 59.975000 105.040000 ;
      RECT 56.985000 105.040000 60.045000 105.110000 ;
      RECT 56.985000 105.040000 60.045000 105.110000 ;
      RECT 56.985000 105.110000 60.115000 105.180000 ;
      RECT 56.985000 105.110000 60.115000 105.180000 ;
      RECT 56.985000 105.180000 60.185000 105.250000 ;
      RECT 56.985000 105.180000 60.185000 105.250000 ;
      RECT 56.985000 105.250000 60.255000 105.320000 ;
      RECT 56.985000 105.250000 60.255000 105.320000 ;
      RECT 56.985000 105.320000 60.325000 105.390000 ;
      RECT 56.985000 105.320000 60.325000 105.390000 ;
      RECT 56.985000 105.390000 60.395000 105.460000 ;
      RECT 56.985000 105.390000 60.395000 105.460000 ;
      RECT 56.985000 105.460000 60.465000 105.530000 ;
      RECT 56.985000 105.460000 60.465000 105.530000 ;
      RECT 56.985000 105.530000 60.535000 105.600000 ;
      RECT 56.985000 105.530000 60.535000 105.600000 ;
      RECT 56.985000 105.600000 60.605000 105.670000 ;
      RECT 56.985000 105.600000 60.605000 105.670000 ;
      RECT 56.985000 105.670000 60.675000 105.740000 ;
      RECT 56.985000 105.670000 60.675000 105.740000 ;
      RECT 56.985000 105.740000 60.745000 105.810000 ;
      RECT 56.985000 105.740000 60.745000 105.810000 ;
      RECT 56.985000 105.770000 60.970000 112.760000 ;
      RECT 56.985000 105.810000 60.815000 105.825000 ;
      RECT 56.985000 105.810000 60.815000 105.825000 ;
      RECT 56.985000 105.825000 60.830000 112.705000 ;
      RECT 56.985000 112.705000 60.805000 112.730000 ;
      RECT 56.985000 112.705000 60.805000 112.730000 ;
      RECT 56.985000 112.730000 60.775000 112.760000 ;
      RECT 56.985000 112.730000 60.775000 112.760000 ;
      RECT 56.985000 125.435000 57.440000 125.505000 ;
      RECT 56.985000 125.435000 57.440000 125.505000 ;
      RECT 56.985000 125.505000 57.510000 125.575000 ;
      RECT 56.985000 125.505000 57.510000 125.575000 ;
      RECT 56.985000 125.575000 57.580000 125.645000 ;
      RECT 56.985000 125.575000 57.580000 125.645000 ;
      RECT 56.985000 125.645000 57.650000 125.715000 ;
      RECT 56.985000 125.645000 57.650000 125.715000 ;
      RECT 56.985000 125.715000 57.720000 125.785000 ;
      RECT 56.985000 125.715000 57.720000 125.785000 ;
      RECT 56.985000 125.785000 57.790000 125.855000 ;
      RECT 56.985000 125.785000 57.790000 125.855000 ;
      RECT 56.985000 125.855000 57.860000 125.925000 ;
      RECT 56.985000 125.855000 57.860000 125.925000 ;
      RECT 56.985000 125.925000 57.930000 125.995000 ;
      RECT 56.985000 125.925000 57.930000 125.995000 ;
      RECT 56.985000 125.995000 58.000000 126.065000 ;
      RECT 56.985000 125.995000 58.000000 126.065000 ;
      RECT 56.985000 126.065000 58.070000 126.135000 ;
      RECT 56.985000 126.065000 58.070000 126.135000 ;
      RECT 56.985000 126.135000 58.140000 126.205000 ;
      RECT 56.985000 126.135000 58.140000 126.205000 ;
      RECT 56.985000 126.205000 58.210000 126.275000 ;
      RECT 56.985000 126.205000 58.210000 126.275000 ;
      RECT 56.985000 126.275000 58.280000 126.345000 ;
      RECT 56.985000 126.275000 58.280000 126.345000 ;
      RECT 56.985000 126.345000 58.350000 126.415000 ;
      RECT 56.985000 126.345000 58.350000 126.415000 ;
      RECT 56.985000 126.415000 58.420000 126.485000 ;
      RECT 56.985000 126.415000 58.420000 126.485000 ;
      RECT 56.985000 126.485000 58.490000 126.500000 ;
      RECT 56.985000 126.485000 58.490000 126.500000 ;
      RECT 56.985000 126.500000 58.505000 126.570000 ;
      RECT 56.985000 126.500000 58.505000 126.570000 ;
      RECT 56.985000 126.500000 60.970000 128.770000 ;
      RECT 56.985000 126.570000 58.575000 126.640000 ;
      RECT 56.985000 126.570000 58.575000 126.640000 ;
      RECT 56.985000 126.640000 58.645000 126.710000 ;
      RECT 56.985000 126.640000 58.645000 126.710000 ;
      RECT 56.985000 126.710000 58.715000 126.780000 ;
      RECT 56.985000 126.710000 58.715000 126.780000 ;
      RECT 56.985000 126.780000 58.785000 126.850000 ;
      RECT 56.985000 126.780000 58.785000 126.850000 ;
      RECT 56.985000 126.850000 58.855000 126.920000 ;
      RECT 56.985000 126.850000 58.855000 126.920000 ;
      RECT 56.985000 126.920000 58.925000 126.990000 ;
      RECT 56.985000 126.920000 58.925000 126.990000 ;
      RECT 56.985000 126.990000 58.995000 127.060000 ;
      RECT 56.985000 126.990000 58.995000 127.060000 ;
      RECT 56.985000 127.060000 59.065000 127.130000 ;
      RECT 56.985000 127.060000 59.065000 127.130000 ;
      RECT 56.985000 127.130000 59.135000 127.200000 ;
      RECT 56.985000 127.130000 59.135000 127.200000 ;
      RECT 56.985000 127.200000 59.205000 127.270000 ;
      RECT 56.985000 127.200000 59.205000 127.270000 ;
      RECT 56.985000 127.270000 59.275000 127.340000 ;
      RECT 56.985000 127.270000 59.275000 127.340000 ;
      RECT 56.985000 127.340000 59.345000 127.410000 ;
      RECT 56.985000 127.340000 59.345000 127.410000 ;
      RECT 56.985000 127.410000 59.415000 127.480000 ;
      RECT 56.985000 127.410000 59.415000 127.480000 ;
      RECT 56.985000 127.480000 59.485000 127.550000 ;
      RECT 56.985000 127.480000 59.485000 127.550000 ;
      RECT 56.985000 127.550000 59.555000 127.620000 ;
      RECT 56.985000 127.550000 59.555000 127.620000 ;
      RECT 56.985000 127.620000 59.625000 127.690000 ;
      RECT 56.985000 127.620000 59.625000 127.690000 ;
      RECT 56.985000 127.690000 59.695000 127.760000 ;
      RECT 56.985000 127.690000 59.695000 127.760000 ;
      RECT 56.985000 127.760000 59.765000 127.830000 ;
      RECT 56.985000 127.760000 59.765000 127.830000 ;
      RECT 56.985000 127.830000 59.835000 127.900000 ;
      RECT 56.985000 127.830000 59.835000 127.900000 ;
      RECT 56.985000 127.900000 59.905000 127.970000 ;
      RECT 56.985000 127.900000 59.905000 127.970000 ;
      RECT 56.985000 127.970000 59.975000 128.040000 ;
      RECT 56.985000 127.970000 59.975000 128.040000 ;
      RECT 56.985000 128.040000 60.045000 128.110000 ;
      RECT 56.985000 128.040000 60.045000 128.110000 ;
      RECT 56.985000 128.110000 60.115000 128.180000 ;
      RECT 56.985000 128.110000 60.115000 128.180000 ;
      RECT 56.985000 128.180000 60.185000 128.250000 ;
      RECT 56.985000 128.180000 60.185000 128.250000 ;
      RECT 56.985000 128.250000 60.255000 128.320000 ;
      RECT 56.985000 128.250000 60.255000 128.320000 ;
      RECT 56.985000 128.320000 60.325000 128.390000 ;
      RECT 56.985000 128.320000 60.325000 128.390000 ;
      RECT 56.985000 128.390000 60.395000 128.460000 ;
      RECT 56.985000 128.390000 60.395000 128.460000 ;
      RECT 56.985000 128.460000 60.465000 128.530000 ;
      RECT 56.985000 128.460000 60.465000 128.530000 ;
      RECT 56.985000 128.530000 60.535000 128.600000 ;
      RECT 56.985000 128.530000 60.535000 128.600000 ;
      RECT 56.985000 128.600000 60.605000 128.670000 ;
      RECT 56.985000 128.600000 60.605000 128.670000 ;
      RECT 56.985000 128.670000 60.675000 128.740000 ;
      RECT 56.985000 128.670000 60.675000 128.740000 ;
      RECT 56.985000 128.740000 60.745000 128.810000 ;
      RECT 56.985000 128.740000 60.745000 128.810000 ;
      RECT 56.985000 128.770000 60.970000 135.760000 ;
      RECT 56.985000 128.810000 60.815000 128.825000 ;
      RECT 56.985000 128.810000 60.815000 128.825000 ;
      RECT 56.985000 128.825000 60.830000 135.740000 ;
      RECT 56.985000 135.740000 60.820000 135.750000 ;
      RECT 56.985000 135.740000 60.820000 135.750000 ;
      RECT 56.985000 135.750000 60.810000 135.760000 ;
      RECT 56.985000 135.750000 60.810000 135.760000 ;
      RECT 56.985000 148.435000 57.370000 148.505000 ;
      RECT 56.985000 148.435000 57.370000 148.505000 ;
      RECT 56.985000 148.505000 57.440000 148.575000 ;
      RECT 56.985000 148.505000 57.440000 148.575000 ;
      RECT 56.985000 148.575000 57.510000 148.645000 ;
      RECT 56.985000 148.575000 57.510000 148.645000 ;
      RECT 56.985000 148.645000 57.580000 148.715000 ;
      RECT 56.985000 148.645000 57.580000 148.715000 ;
      RECT 56.985000 148.715000 57.650000 148.785000 ;
      RECT 56.985000 148.715000 57.650000 148.785000 ;
      RECT 56.985000 148.785000 57.720000 148.855000 ;
      RECT 56.985000 148.785000 57.720000 148.855000 ;
      RECT 56.985000 148.855000 57.790000 148.925000 ;
      RECT 56.985000 148.855000 57.790000 148.925000 ;
      RECT 56.985000 148.925000 57.860000 148.995000 ;
      RECT 56.985000 148.925000 57.860000 148.995000 ;
      RECT 56.985000 148.995000 57.930000 149.065000 ;
      RECT 56.985000 148.995000 57.930000 149.065000 ;
      RECT 56.985000 149.065000 58.000000 149.135000 ;
      RECT 56.985000 149.065000 58.000000 149.135000 ;
      RECT 56.985000 149.135000 58.070000 149.205000 ;
      RECT 56.985000 149.135000 58.070000 149.205000 ;
      RECT 56.985000 149.205000 58.140000 149.275000 ;
      RECT 56.985000 149.205000 58.140000 149.275000 ;
      RECT 56.985000 149.275000 58.210000 149.345000 ;
      RECT 56.985000 149.275000 58.210000 149.345000 ;
      RECT 56.985000 149.345000 58.280000 149.415000 ;
      RECT 56.985000 149.345000 58.280000 149.415000 ;
      RECT 56.985000 149.415000 58.350000 149.485000 ;
      RECT 56.985000 149.415000 58.350000 149.485000 ;
      RECT 56.985000 149.485000 58.420000 149.500000 ;
      RECT 56.985000 149.485000 58.420000 149.500000 ;
      RECT 56.985000 149.500000 58.435000 149.570000 ;
      RECT 56.985000 149.500000 58.435000 149.570000 ;
      RECT 56.985000 149.500000 60.970000 151.840000 ;
      RECT 56.985000 149.570000 58.505000 149.640000 ;
      RECT 56.985000 149.570000 58.505000 149.640000 ;
      RECT 56.985000 149.640000 58.575000 149.710000 ;
      RECT 56.985000 149.640000 58.575000 149.710000 ;
      RECT 56.985000 149.710000 58.645000 149.780000 ;
      RECT 56.985000 149.710000 58.645000 149.780000 ;
      RECT 56.985000 149.780000 58.715000 149.850000 ;
      RECT 56.985000 149.780000 58.715000 149.850000 ;
      RECT 56.985000 149.850000 58.785000 149.920000 ;
      RECT 56.985000 149.850000 58.785000 149.920000 ;
      RECT 56.985000 149.920000 58.855000 149.990000 ;
      RECT 56.985000 149.920000 58.855000 149.990000 ;
      RECT 56.985000 149.990000 58.925000 150.060000 ;
      RECT 56.985000 149.990000 58.925000 150.060000 ;
      RECT 56.985000 150.060000 58.995000 150.130000 ;
      RECT 56.985000 150.060000 58.995000 150.130000 ;
      RECT 56.985000 150.130000 59.065000 150.200000 ;
      RECT 56.985000 150.130000 59.065000 150.200000 ;
      RECT 56.985000 150.200000 59.135000 150.270000 ;
      RECT 56.985000 150.200000 59.135000 150.270000 ;
      RECT 56.985000 150.270000 59.205000 150.340000 ;
      RECT 56.985000 150.270000 59.205000 150.340000 ;
      RECT 56.985000 150.340000 59.275000 150.410000 ;
      RECT 56.985000 150.340000 59.275000 150.410000 ;
      RECT 56.985000 150.410000 59.345000 150.480000 ;
      RECT 56.985000 150.410000 59.345000 150.480000 ;
      RECT 56.985000 150.480000 59.415000 150.550000 ;
      RECT 56.985000 150.480000 59.415000 150.550000 ;
      RECT 56.985000 150.550000 59.485000 150.620000 ;
      RECT 56.985000 150.550000 59.485000 150.620000 ;
      RECT 56.985000 150.620000 59.555000 150.690000 ;
      RECT 56.985000 150.620000 59.555000 150.690000 ;
      RECT 56.985000 150.690000 59.625000 150.760000 ;
      RECT 56.985000 150.690000 59.625000 150.760000 ;
      RECT 56.985000 150.760000 59.695000 150.830000 ;
      RECT 56.985000 150.760000 59.695000 150.830000 ;
      RECT 56.985000 150.830000 59.765000 150.900000 ;
      RECT 56.985000 150.830000 59.765000 150.900000 ;
      RECT 56.985000 150.900000 59.835000 150.970000 ;
      RECT 56.985000 150.900000 59.835000 150.970000 ;
      RECT 56.985000 150.970000 59.905000 151.040000 ;
      RECT 56.985000 150.970000 59.905000 151.040000 ;
      RECT 56.985000 151.040000 59.975000 151.110000 ;
      RECT 56.985000 151.040000 59.975000 151.110000 ;
      RECT 56.985000 151.110000 60.045000 151.180000 ;
      RECT 56.985000 151.110000 60.045000 151.180000 ;
      RECT 56.985000 151.180000 60.115000 151.250000 ;
      RECT 56.985000 151.180000 60.115000 151.250000 ;
      RECT 56.985000 151.250000 60.185000 151.320000 ;
      RECT 56.985000 151.250000 60.185000 151.320000 ;
      RECT 56.985000 151.320000 60.255000 151.390000 ;
      RECT 56.985000 151.320000 60.255000 151.390000 ;
      RECT 56.985000 151.390000 60.325000 151.460000 ;
      RECT 56.985000 151.390000 60.325000 151.460000 ;
      RECT 56.985000 151.460000 60.395000 151.530000 ;
      RECT 56.985000 151.460000 60.395000 151.530000 ;
      RECT 56.985000 151.530000 60.465000 151.600000 ;
      RECT 56.985000 151.530000 60.465000 151.600000 ;
      RECT 56.985000 151.600000 60.535000 151.670000 ;
      RECT 56.985000 151.600000 60.535000 151.670000 ;
      RECT 56.985000 151.670000 60.605000 151.740000 ;
      RECT 56.985000 151.670000 60.605000 151.740000 ;
      RECT 56.985000 151.740000 60.675000 151.810000 ;
      RECT 56.985000 151.740000 60.675000 151.810000 ;
      RECT 56.985000 151.810000 60.745000 151.880000 ;
      RECT 56.985000 151.810000 60.745000 151.880000 ;
      RECT 56.985000 151.840000 60.970000 158.760000 ;
      RECT 56.985000 151.880000 60.815000 151.895000 ;
      RECT 56.985000 151.880000 60.815000 151.895000 ;
      RECT 56.985000 151.895000 60.830000 158.755000 ;
      RECT 56.985000 158.755000 60.825000 158.760000 ;
      RECT 56.985000 158.755000 60.825000 158.760000 ;
      RECT 56.990000  56.435000 57.410000  56.505000 ;
      RECT 56.990000  56.435000 57.410000  56.505000 ;
      RECT 56.990000  56.505000 57.480000  56.575000 ;
      RECT 56.990000  56.505000 57.480000  56.575000 ;
      RECT 56.990000  56.575000 57.550000  56.645000 ;
      RECT 56.990000  56.575000 57.550000  56.645000 ;
      RECT 56.990000  56.645000 57.620000  56.715000 ;
      RECT 56.990000  56.645000 57.620000  56.715000 ;
      RECT 56.990000  56.715000 57.690000  56.785000 ;
      RECT 56.990000  56.715000 57.690000  56.785000 ;
      RECT 56.990000  56.785000 57.760000  56.855000 ;
      RECT 56.990000  56.785000 57.760000  56.855000 ;
      RECT 56.990000  56.855000 57.830000  56.925000 ;
      RECT 56.990000  56.855000 57.830000  56.925000 ;
      RECT 56.990000  56.925000 57.900000  56.995000 ;
      RECT 56.990000  56.925000 57.900000  56.995000 ;
      RECT 56.990000  56.995000 57.970000  57.065000 ;
      RECT 56.990000  56.995000 57.970000  57.065000 ;
      RECT 56.990000  57.065000 58.040000  57.135000 ;
      RECT 56.990000  57.065000 58.040000  57.135000 ;
      RECT 56.990000  57.135000 58.110000  57.205000 ;
      RECT 56.990000  57.135000 58.110000  57.205000 ;
      RECT 56.990000  57.205000 58.180000  57.275000 ;
      RECT 56.990000  57.205000 58.180000  57.275000 ;
      RECT 56.990000  57.275000 58.250000  57.345000 ;
      RECT 56.990000  57.275000 58.250000  57.345000 ;
      RECT 56.990000  57.345000 58.320000  57.415000 ;
      RECT 56.990000  57.345000 58.320000  57.415000 ;
      RECT 56.990000  57.415000 58.390000  57.485000 ;
      RECT 56.990000  57.415000 58.390000  57.485000 ;
      RECT 56.990000  57.485000 58.460000  57.500000 ;
      RECT 56.990000  57.485000 58.460000  57.500000 ;
      RECT 56.990000  57.500000 58.475000  57.570000 ;
      RECT 56.990000  57.500000 58.475000  57.570000 ;
      RECT 56.990000  57.500000 60.970000  59.800000 ;
      RECT 56.990000  57.570000 58.545000  57.640000 ;
      RECT 56.990000  57.570000 58.545000  57.640000 ;
      RECT 56.990000  57.640000 58.615000  57.710000 ;
      RECT 56.990000  57.640000 58.615000  57.710000 ;
      RECT 56.990000  57.710000 58.685000  57.780000 ;
      RECT 56.990000  57.710000 58.685000  57.780000 ;
      RECT 56.990000  57.780000 58.755000  57.850000 ;
      RECT 56.990000  57.780000 58.755000  57.850000 ;
      RECT 56.990000  57.850000 58.825000  57.920000 ;
      RECT 56.990000  57.850000 58.825000  57.920000 ;
      RECT 56.990000  57.920000 58.895000  57.990000 ;
      RECT 56.990000  57.920000 58.895000  57.990000 ;
      RECT 56.990000  57.990000 58.965000  58.060000 ;
      RECT 56.990000  57.990000 58.965000  58.060000 ;
      RECT 56.990000  58.060000 59.035000  58.130000 ;
      RECT 56.990000  58.060000 59.035000  58.130000 ;
      RECT 56.990000  58.130000 59.105000  58.200000 ;
      RECT 56.990000  58.130000 59.105000  58.200000 ;
      RECT 56.990000  58.200000 59.175000  58.270000 ;
      RECT 56.990000  58.200000 59.175000  58.270000 ;
      RECT 56.990000  58.270000 59.245000  58.340000 ;
      RECT 56.990000  58.270000 59.245000  58.340000 ;
      RECT 56.990000  58.340000 59.315000  58.410000 ;
      RECT 56.990000  58.340000 59.315000  58.410000 ;
      RECT 56.990000  58.410000 59.385000  58.480000 ;
      RECT 56.990000  58.410000 59.385000  58.480000 ;
      RECT 56.990000  58.480000 59.455000  58.550000 ;
      RECT 56.990000  58.480000 59.455000  58.550000 ;
      RECT 56.990000  58.550000 59.525000  58.620000 ;
      RECT 56.990000  58.550000 59.525000  58.620000 ;
      RECT 56.990000  58.620000 59.595000  58.690000 ;
      RECT 56.990000  58.620000 59.595000  58.690000 ;
      RECT 56.990000  58.690000 59.665000  58.760000 ;
      RECT 56.990000  58.690000 59.665000  58.760000 ;
      RECT 56.990000  58.760000 59.735000  58.830000 ;
      RECT 56.990000  58.760000 59.735000  58.830000 ;
      RECT 56.990000  58.830000 59.805000  58.900000 ;
      RECT 56.990000  58.830000 59.805000  58.900000 ;
      RECT 56.990000  58.900000 59.875000  58.970000 ;
      RECT 56.990000  58.900000 59.875000  58.970000 ;
      RECT 56.990000  58.970000 59.945000  59.040000 ;
      RECT 56.990000  58.970000 59.945000  59.040000 ;
      RECT 56.990000  59.040000 60.015000  59.110000 ;
      RECT 56.990000  59.040000 60.015000  59.110000 ;
      RECT 56.990000  59.110000 60.085000  59.180000 ;
      RECT 56.990000  59.110000 60.085000  59.180000 ;
      RECT 56.990000  59.180000 60.155000  59.250000 ;
      RECT 56.990000  59.180000 60.155000  59.250000 ;
      RECT 56.990000  59.250000 60.225000  59.320000 ;
      RECT 56.990000  59.250000 60.225000  59.320000 ;
      RECT 56.990000  59.320000 60.295000  59.390000 ;
      RECT 56.990000  59.320000 60.295000  59.390000 ;
      RECT 56.990000  59.390000 60.365000  59.460000 ;
      RECT 56.990000  59.390000 60.365000  59.460000 ;
      RECT 56.990000  59.460000 60.435000  59.530000 ;
      RECT 56.990000  59.460000 60.435000  59.530000 ;
      RECT 56.990000  59.530000 60.505000  59.600000 ;
      RECT 56.990000  59.530000 60.505000  59.600000 ;
      RECT 56.990000  59.600000 60.575000  59.670000 ;
      RECT 56.990000  59.600000 60.575000  59.670000 ;
      RECT 56.990000  59.670000 60.645000  59.740000 ;
      RECT 56.990000  59.670000 60.645000  59.740000 ;
      RECT 56.990000  59.740000 60.715000  59.810000 ;
      RECT 56.990000  59.740000 60.715000  59.810000 ;
      RECT 56.990000  59.800000 60.970000  66.760000 ;
      RECT 56.990000  59.810000 60.785000  59.855000 ;
      RECT 56.990000  59.810000 60.785000  59.855000 ;
      RECT 56.990000  59.855000 60.830000  66.735000 ;
      RECT 56.990000  66.735000 60.820000  66.745000 ;
      RECT 56.990000  66.735000 60.820000  66.745000 ;
      RECT 56.990000  66.745000 60.805000  66.760000 ;
      RECT 56.990000  66.745000 60.805000  66.760000 ;
      RECT 57.055000  35.975000 60.970000  39.725000 ;
      RECT 57.055000  39.725000 60.970000  42.520000 ;
      RECT 57.055000  39.920000 60.830000  39.990000 ;
      RECT 57.055000  39.920000 60.830000  39.990000 ;
      RECT 57.125000  39.850000 60.830000  39.920000 ;
      RECT 57.125000  39.850000 60.830000  39.920000 ;
      RECT 57.195000  35.835000 60.830000  39.780000 ;
      RECT 57.195000  39.780000 60.830000  39.850000 ;
      RECT 57.195000  39.780000 60.830000  39.850000 ;
      RECT 58.240000 172.500000 58.515000 172.570000 ;
      RECT 58.240000 172.500000 60.970000 174.760000 ;
      RECT 58.240000 172.570000 58.585000 172.640000 ;
      RECT 58.240000 172.640000 58.655000 172.710000 ;
      RECT 58.240000 172.710000 58.725000 172.780000 ;
      RECT 58.240000 172.780000 58.795000 172.850000 ;
      RECT 58.240000 172.850000 58.865000 172.920000 ;
      RECT 58.240000 172.920000 58.935000 172.990000 ;
      RECT 58.240000 172.990000 59.005000 173.060000 ;
      RECT 58.240000 173.060000 59.075000 173.130000 ;
      RECT 58.240000 173.130000 59.145000 173.200000 ;
      RECT 58.240000 173.200000 59.215000 173.270000 ;
      RECT 58.240000 173.270000 59.285000 173.340000 ;
      RECT 58.240000 173.340000 59.355000 173.410000 ;
      RECT 58.240000 173.410000 59.425000 173.480000 ;
      RECT 58.240000 173.480000 59.495000 173.550000 ;
      RECT 58.240000 173.550000 59.565000 173.620000 ;
      RECT 58.240000 173.620000 59.635000 173.690000 ;
      RECT 58.240000 173.690000 59.705000 173.760000 ;
      RECT 58.240000 173.760000 59.775000 173.830000 ;
      RECT 58.240000 173.830000 59.845000 173.900000 ;
      RECT 58.240000 173.900000 59.915000 173.970000 ;
      RECT 58.240000 173.970000 59.985000 174.040000 ;
      RECT 58.240000 174.040000 60.055000 174.110000 ;
      RECT 58.240000 174.110000 60.125000 174.180000 ;
      RECT 58.240000 174.180000 60.195000 174.250000 ;
      RECT 58.240000 174.250000 60.265000 174.320000 ;
      RECT 58.240000 174.320000 60.335000 174.390000 ;
      RECT 58.240000 174.390000 60.405000 174.460000 ;
      RECT 58.240000 174.460000 60.475000 174.530000 ;
      RECT 58.240000 174.530000 60.545000 174.600000 ;
      RECT 58.240000 174.600000 60.615000 174.670000 ;
      RECT 58.240000 174.670000 60.685000 174.740000 ;
      RECT 58.240000 174.740000 60.755000 174.810000 ;
      RECT 58.240000 174.760000 60.970000 181.760000 ;
      RECT 58.240000 174.810000 60.825000 174.815000 ;
      RECT 58.240000 174.815000 60.830000 181.760000 ;
      RECT 67.480000 190.280000 75.000000 195.355000 ;
      RECT 67.480000 190.295000 75.000000 200.000000 ;
      RECT 70.480000 193.295000 72.000000 197.000000 ;
      RECT 74.430000   0.000000 75.000000 190.155000 ;
      RECT 74.570000   0.000000 75.000000 190.295000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.195000  36.635000 ;
      RECT  0.000000  36.635000  0.670000  37.110000 ;
      RECT  0.000000  36.730000  0.150000  36.880000 ;
      RECT  0.000000  36.880000  0.300000  37.030000 ;
      RECT  0.000000  37.030000  0.450000  37.150000 ;
      RECT  0.000000  37.110000  0.670000  46.360000 ;
      RECT  0.000000  37.150000  0.570000  46.320000 ;
      RECT  0.000000  46.320000  0.420000  46.470000 ;
      RECT  0.000000  46.360000  0.195000  46.835000 ;
      RECT  0.000000  46.470000  0.270000  46.620000 ;
      RECT  0.000000  46.620000  0.120000  46.770000 ;
      RECT  0.000000  46.835000  0.195000 173.455000 ;
      RECT  0.000000 173.455000 13.650000 195.500000 ;
      RECT  0.000000 173.555000 13.650000 195.500000 ;
      RECT  0.000000 173.555000 13.650000 200.000000 ;
      RECT  0.000000 195.500000 75.000000 200.000000 ;
      RECT  0.000000 195.500000 75.000000 200.000000 ;
      RECT 13.800000 101.520000 15.100000 102.035000 ;
      RECT 13.800000 102.035000 15.100000 171.140000 ;
      RECT 13.900000 101.560000 15.425000 101.710000 ;
      RECT 13.900000 101.710000 15.275000 101.860000 ;
      RECT 13.900000 101.860000 15.125000 102.010000 ;
      RECT 13.900000 102.010000 15.100000 102.035000 ;
      RECT 13.900000 102.035000 15.100000 171.140000 ;
      RECT 13.900000 171.140000 14.950000 171.290000 ;
      RECT 13.900000 171.290000 14.800000 171.440000 ;
      RECT 13.900000 171.440000 14.650000 171.590000 ;
      RECT 13.900000 171.590000 14.500000 171.740000 ;
      RECT 13.900000 171.740000 14.350000 171.890000 ;
      RECT 13.900000 171.890000 14.200000 172.040000 ;
      RECT 13.900000 172.040000 14.050000 172.190000 ;
      RECT 14.020000 101.440000 15.575000 101.560000 ;
      RECT 14.170000 101.290000 15.695000 101.440000 ;
      RECT 14.320000 101.140000 15.845000 101.290000 ;
      RECT 14.470000 100.990000 15.995000 101.140000 ;
      RECT 14.620000 100.840000 16.145000 100.990000 ;
      RECT 14.770000 100.690000 16.295000 100.840000 ;
      RECT 14.920000 100.540000 16.445000 100.690000 ;
      RECT 15.070000 100.390000 16.595000 100.540000 ;
      RECT 15.220000 100.240000 16.745000 100.390000 ;
      RECT 15.370000 100.090000 16.895000 100.240000 ;
      RECT 15.520000  99.940000 17.045000 100.090000 ;
      RECT 15.670000  99.790000 17.195000  99.940000 ;
      RECT 15.820000  99.640000 17.345000  99.790000 ;
      RECT 15.970000  99.490000 17.495000  99.640000 ;
      RECT 16.120000  99.340000 17.645000  99.490000 ;
      RECT 16.270000  99.190000 17.795000  99.340000 ;
      RECT 16.420000  99.040000 17.945000  99.190000 ;
      RECT 16.570000  98.890000 18.095000  99.040000 ;
      RECT 16.720000  98.740000 18.245000  98.890000 ;
      RECT 16.870000  98.590000 18.395000  98.740000 ;
      RECT 17.020000  98.440000 18.545000  98.590000 ;
      RECT 17.170000  98.290000 18.695000  98.440000 ;
      RECT 17.320000  98.140000 18.845000  98.290000 ;
      RECT 17.470000  97.990000 18.995000  98.140000 ;
      RECT 17.620000  97.840000 19.145000  97.990000 ;
      RECT 17.770000  97.690000 19.295000  97.840000 ;
      RECT 17.920000  97.540000 19.445000  97.690000 ;
      RECT 18.070000  97.390000 19.595000  97.540000 ;
      RECT 18.220000  97.240000 19.745000  97.390000 ;
      RECT 18.370000  97.090000 19.895000  97.240000 ;
      RECT 18.520000  96.940000 20.045000  97.090000 ;
      RECT 18.670000  96.790000 20.195000  96.940000 ;
      RECT 18.820000  96.640000 20.345000  96.790000 ;
      RECT 18.970000  96.490000 20.495000  96.640000 ;
      RECT 19.120000  96.340000 20.645000  96.490000 ;
      RECT 19.270000  96.190000 20.795000  96.340000 ;
      RECT 19.420000  96.040000 20.945000  96.190000 ;
      RECT 19.570000  95.890000 21.095000  96.040000 ;
      RECT 19.720000  95.740000 21.245000  95.890000 ;
      RECT 19.870000  95.590000 21.395000  95.740000 ;
      RECT 20.020000  95.440000 21.545000  95.590000 ;
      RECT 20.170000  95.290000 21.695000  95.440000 ;
      RECT 20.320000  95.140000 21.845000  95.290000 ;
      RECT 20.470000  94.990000 21.995000  95.140000 ;
      RECT 20.620000  94.840000 22.145000  94.990000 ;
      RECT 20.770000  94.690000 22.295000  94.840000 ;
      RECT 20.920000  94.540000 22.445000  94.690000 ;
      RECT 21.070000  94.390000 22.595000  94.540000 ;
      RECT 21.220000  94.240000 22.745000  94.390000 ;
      RECT 21.370000  94.090000 22.895000  94.240000 ;
      RECT 21.520000  93.940000 23.045000  94.090000 ;
      RECT 21.670000  93.790000 23.195000  93.940000 ;
      RECT 21.695000  93.765000 23.345000  93.790000 ;
      RECT 21.845000  93.615000 23.345000  93.765000 ;
      RECT 21.900000 104.845000 25.530000 168.965000 ;
      RECT 21.900000 104.845000 25.530000 168.965000 ;
      RECT 21.900000 168.965000 25.530000 172.475000 ;
      RECT 21.970000 104.775000 25.530000 104.845000 ;
      RECT 21.995000  93.465000 23.345000  93.615000 ;
      RECT 22.050000 168.965000 25.530000 169.115000 ;
      RECT 22.120000 104.625000 25.530000 104.775000 ;
      RECT 22.145000  93.315000 23.345000  93.465000 ;
      RECT 22.200000 169.115000 25.530000 169.265000 ;
      RECT 22.270000 104.475000 25.530000 104.625000 ;
      RECT 22.295000  93.165000 23.345000  93.315000 ;
      RECT 22.350000 169.265000 25.530000 169.415000 ;
      RECT 22.420000 104.325000 25.530000 104.475000 ;
      RECT 22.445000  93.015000 23.345000  93.165000 ;
      RECT 22.500000 169.415000 25.530000 169.565000 ;
      RECT 22.570000 104.175000 25.530000 104.325000 ;
      RECT 22.595000  92.865000 23.345000  93.015000 ;
      RECT 22.650000 169.565000 25.530000 169.715000 ;
      RECT 22.720000 104.025000 25.530000 104.175000 ;
      RECT 22.745000  92.715000 23.345000  92.865000 ;
      RECT 22.800000 169.715000 25.530000 169.865000 ;
      RECT 22.870000 103.875000 25.530000 104.025000 ;
      RECT 22.895000  92.565000 23.345000  92.715000 ;
      RECT 22.945000  92.375000 23.345000  93.790000 ;
      RECT 22.950000 169.865000 25.530000 170.015000 ;
      RECT 23.020000 103.725000 25.530000 103.875000 ;
      RECT 23.045000  92.415000 23.345000  92.565000 ;
      RECT 23.100000 170.015000 25.530000 170.165000 ;
      RECT 23.170000 103.575000 25.530000 103.725000 ;
      RECT 23.195000  92.265000 23.345000  92.415000 ;
      RECT 23.250000 170.165000 25.530000 170.315000 ;
      RECT 23.320000 103.425000 25.530000 103.575000 ;
      RECT 23.400000 170.315000 25.530000 170.465000 ;
      RECT 23.470000 103.275000 25.530000 103.425000 ;
      RECT 23.550000 170.465000 25.530000 170.615000 ;
      RECT 23.620000 103.125000 25.530000 103.275000 ;
      RECT 23.700000 170.615000 25.530000 170.765000 ;
      RECT 23.770000 102.975000 25.530000 103.125000 ;
      RECT 23.850000 170.765000 25.530000 170.915000 ;
      RECT 23.920000 102.825000 25.530000 102.975000 ;
      RECT 24.000000 170.915000 25.530000 171.065000 ;
      RECT 24.070000 102.675000 25.530000 102.825000 ;
      RECT 24.150000 171.065000 25.530000 171.215000 ;
      RECT 24.220000 102.525000 25.530000 102.675000 ;
      RECT 24.300000 171.215000 25.530000 171.365000 ;
      RECT 24.370000 102.375000 25.530000 102.525000 ;
      RECT 24.450000 171.365000 25.530000 171.515000 ;
      RECT 24.520000 102.225000 25.530000 102.375000 ;
      RECT 24.520000 102.225000 25.530000 104.845000 ;
      RECT 24.525000 102.220000 25.530000 102.225000 ;
      RECT 24.600000 171.515000 25.530000 171.665000 ;
      RECT 24.675000 102.070000 25.535000 102.220000 ;
      RECT 24.695000   0.000000 25.495000  90.225000 ;
      RECT 24.695000  90.225000 25.095000  90.625000 ;
      RECT 24.750000 171.665000 25.530000 171.815000 ;
      RECT 24.795000   0.000000 25.495000  90.225000 ;
      RECT 24.795000  90.225000 25.345000  90.375000 ;
      RECT 24.795000  90.375000 25.195000  90.525000 ;
      RECT 24.795000  90.525000 25.045000  90.675000 ;
      RECT 24.795000  90.675000 24.895000  90.825000 ;
      RECT 24.825000 101.920000 25.685000 102.070000 ;
      RECT 24.900000 171.815000 25.530000 171.965000 ;
      RECT 24.975000 101.770000 25.835000 101.920000 ;
      RECT 25.050000 171.965000 25.530000 172.115000 ;
      RECT 25.125000 101.620000 25.985000 101.770000 ;
      RECT 25.200000 172.115000 25.530000 172.265000 ;
      RECT 25.275000 101.470000 26.135000 101.620000 ;
      RECT 25.350000 172.265000 25.530000 172.415000 ;
      RECT 25.410000 172.475000 25.530000 195.500000 ;
      RECT 25.425000 101.320000 26.285000 101.470000 ;
      RECT 25.500000 172.415000 25.530000 172.565000 ;
      RECT 25.575000 101.170000 26.435000 101.320000 ;
      RECT 25.725000 101.020000 26.585000 101.170000 ;
      RECT 25.875000 100.870000 26.735000 101.020000 ;
      RECT 26.025000 100.720000 26.885000 100.870000 ;
      RECT 26.175000 100.570000 27.035000 100.720000 ;
      RECT 26.325000 100.420000 27.185000 100.570000 ;
      RECT 26.475000 100.270000 27.335000 100.420000 ;
      RECT 26.625000 100.120000 27.485000 100.270000 ;
      RECT 26.775000  99.970000 27.635000 100.120000 ;
      RECT 26.925000  99.820000 27.785000  99.970000 ;
      RECT 27.075000  99.670000 27.935000  99.820000 ;
      RECT 27.225000  99.520000 28.085000  99.670000 ;
      RECT 27.375000  99.370000 28.235000  99.520000 ;
      RECT 27.525000  99.220000 28.385000  99.370000 ;
      RECT 27.675000  99.070000 28.535000  99.220000 ;
      RECT 27.825000  98.920000 28.685000  99.070000 ;
      RECT 27.975000  98.770000 28.835000  98.920000 ;
      RECT 28.125000  98.620000 28.985000  98.770000 ;
      RECT 28.275000  98.470000 29.135000  98.620000 ;
      RECT 28.425000  98.320000 29.285000  98.470000 ;
      RECT 28.575000  98.170000 29.435000  98.320000 ;
      RECT 28.725000  98.020000 29.585000  98.170000 ;
      RECT 28.875000  97.870000 29.735000  98.020000 ;
      RECT 29.025000  97.720000 29.885000  97.870000 ;
      RECT 29.175000  97.570000 30.035000  97.720000 ;
      RECT 29.325000  97.420000 30.185000  97.570000 ;
      RECT 29.475000  97.270000 30.335000  97.420000 ;
      RECT 29.625000  97.120000 30.485000  97.270000 ;
      RECT 29.775000  96.970000 30.635000  97.120000 ;
      RECT 29.925000  93.265000 31.545000  96.210000 ;
      RECT 29.925000  93.265000 31.545000  96.210000 ;
      RECT 29.925000  96.210000 30.935000  96.820000 ;
      RECT 29.925000  96.210000 31.395000  96.360000 ;
      RECT 29.925000  96.360000 31.245000  96.510000 ;
      RECT 29.925000  96.510000 31.095000  96.660000 ;
      RECT 29.925000  96.660000 30.945000  96.810000 ;
      RECT 29.925000  96.810000 30.935000  96.820000 ;
      RECT 29.925000  96.820000 30.785000  96.970000 ;
      RECT 29.950000  93.240000 31.520000  93.265000 ;
      RECT 30.100000  93.090000 31.370000  93.240000 ;
      RECT 30.250000  92.940000 31.220000  93.090000 ;
      RECT 30.400000  92.790000 31.070000  92.940000 ;
      RECT 30.400000  92.790000 31.545000  93.265000 ;
      RECT 32.330000  99.865000 37.490000 110.785000 ;
      RECT 32.330000 105.025000 37.490000 105.820000 ;
      RECT 32.330000 105.025000 37.490000 105.820000 ;
      RECT 32.330000 105.820000 37.490000 105.970000 ;
      RECT 32.330000 105.820000 37.490000 105.970000 ;
      RECT 32.330000 105.820000 42.455000 110.785000 ;
      RECT 32.330000 105.820000 42.455000 175.185000 ;
      RECT 32.330000 105.970000 37.640000 106.120000 ;
      RECT 32.330000 105.970000 37.640000 106.120000 ;
      RECT 32.330000 106.120000 37.790000 106.270000 ;
      RECT 32.330000 106.120000 37.790000 106.270000 ;
      RECT 32.330000 106.270000 37.940000 106.420000 ;
      RECT 32.330000 106.270000 37.940000 106.420000 ;
      RECT 32.330000 106.420000 38.090000 106.570000 ;
      RECT 32.330000 106.420000 38.090000 106.570000 ;
      RECT 32.330000 106.570000 38.240000 106.720000 ;
      RECT 32.330000 106.570000 38.240000 106.720000 ;
      RECT 32.330000 106.720000 38.390000 106.870000 ;
      RECT 32.330000 106.720000 38.390000 106.870000 ;
      RECT 32.330000 106.870000 38.540000 107.020000 ;
      RECT 32.330000 106.870000 38.540000 107.020000 ;
      RECT 32.330000 107.020000 38.690000 107.170000 ;
      RECT 32.330000 107.020000 38.690000 107.170000 ;
      RECT 32.330000 107.170000 38.840000 107.320000 ;
      RECT 32.330000 107.170000 38.840000 107.320000 ;
      RECT 32.330000 107.320000 38.990000 107.470000 ;
      RECT 32.330000 107.320000 38.990000 107.470000 ;
      RECT 32.330000 107.470000 39.140000 107.620000 ;
      RECT 32.330000 107.470000 39.140000 107.620000 ;
      RECT 32.330000 107.620000 39.290000 107.770000 ;
      RECT 32.330000 107.620000 39.290000 107.770000 ;
      RECT 32.330000 107.770000 39.440000 107.920000 ;
      RECT 32.330000 107.770000 39.440000 107.920000 ;
      RECT 32.330000 107.920000 39.590000 108.070000 ;
      RECT 32.330000 107.920000 39.590000 108.070000 ;
      RECT 32.330000 108.070000 39.740000 108.220000 ;
      RECT 32.330000 108.070000 39.740000 108.220000 ;
      RECT 32.330000 108.220000 39.890000 108.370000 ;
      RECT 32.330000 108.220000 39.890000 108.370000 ;
      RECT 32.330000 108.370000 40.040000 108.520000 ;
      RECT 32.330000 108.370000 40.040000 108.520000 ;
      RECT 32.330000 108.520000 40.190000 108.670000 ;
      RECT 32.330000 108.520000 40.190000 108.670000 ;
      RECT 32.330000 108.670000 40.340000 108.820000 ;
      RECT 32.330000 108.670000 40.340000 108.820000 ;
      RECT 32.330000 108.820000 40.490000 108.970000 ;
      RECT 32.330000 108.820000 40.490000 108.970000 ;
      RECT 32.330000 108.970000 40.640000 109.120000 ;
      RECT 32.330000 108.970000 40.640000 109.120000 ;
      RECT 32.330000 109.120000 40.790000 109.270000 ;
      RECT 32.330000 109.120000 40.790000 109.270000 ;
      RECT 32.330000 109.270000 40.940000 109.420000 ;
      RECT 32.330000 109.270000 40.940000 109.420000 ;
      RECT 32.330000 109.420000 41.090000 109.570000 ;
      RECT 32.330000 109.420000 41.090000 109.570000 ;
      RECT 32.330000 109.570000 41.240000 109.720000 ;
      RECT 32.330000 109.570000 41.240000 109.720000 ;
      RECT 32.330000 109.720000 41.390000 109.870000 ;
      RECT 32.330000 109.720000 41.390000 109.870000 ;
      RECT 32.330000 109.870000 41.540000 110.020000 ;
      RECT 32.330000 109.870000 41.540000 110.020000 ;
      RECT 32.330000 110.020000 41.690000 110.170000 ;
      RECT 32.330000 110.020000 41.690000 110.170000 ;
      RECT 32.330000 110.170000 41.840000 110.320000 ;
      RECT 32.330000 110.170000 41.840000 110.320000 ;
      RECT 32.330000 110.320000 41.990000 110.470000 ;
      RECT 32.330000 110.320000 41.990000 110.470000 ;
      RECT 32.330000 110.470000 42.140000 110.620000 ;
      RECT 32.330000 110.470000 42.140000 110.620000 ;
      RECT 32.330000 110.620000 42.290000 110.770000 ;
      RECT 32.330000 110.620000 42.290000 110.770000 ;
      RECT 32.330000 110.770000 42.440000 110.785000 ;
      RECT 32.330000 110.770000 42.440000 110.785000 ;
      RECT 32.330000 110.785000 42.455000 170.295000 ;
      RECT 32.330000 110.785000 42.455000 170.295000 ;
      RECT 32.330000 170.295000 37.565000 175.185000 ;
      RECT 32.390000 104.965000 37.490000 105.025000 ;
      RECT 32.390000 104.965000 37.490000 105.025000 ;
      RECT 32.480000 170.295000 42.305000 170.445000 ;
      RECT 32.480000 170.295000 42.305000 170.445000 ;
      RECT 32.540000 104.815000 37.490000 104.965000 ;
      RECT 32.540000 104.815000 37.490000 104.965000 ;
      RECT 32.630000 170.445000 42.155000 170.595000 ;
      RECT 32.630000 170.445000 42.155000 170.595000 ;
      RECT 32.690000 104.665000 37.490000 104.815000 ;
      RECT 32.690000 104.665000 37.490000 104.815000 ;
      RECT 32.780000 170.595000 42.005000 170.745000 ;
      RECT 32.780000 170.595000 42.005000 170.745000 ;
      RECT 32.840000 104.515000 37.490000 104.665000 ;
      RECT 32.840000 104.515000 37.490000 104.665000 ;
      RECT 32.930000 170.745000 41.855000 170.895000 ;
      RECT 32.930000 170.745000 41.855000 170.895000 ;
      RECT 32.990000 104.365000 37.490000 104.515000 ;
      RECT 32.990000 104.365000 37.490000 104.515000 ;
      RECT 33.080000 170.895000 41.705000 171.045000 ;
      RECT 33.080000 170.895000 41.705000 171.045000 ;
      RECT 33.140000 104.215000 37.490000 104.365000 ;
      RECT 33.140000 104.215000 37.490000 104.365000 ;
      RECT 33.230000 171.045000 41.555000 171.195000 ;
      RECT 33.230000 171.045000 41.555000 171.195000 ;
      RECT 33.290000 104.065000 37.490000 104.215000 ;
      RECT 33.290000 104.065000 37.490000 104.215000 ;
      RECT 33.380000 171.195000 41.405000 171.345000 ;
      RECT 33.380000 171.195000 41.405000 171.345000 ;
      RECT 33.440000 103.915000 37.490000 104.065000 ;
      RECT 33.440000 103.915000 37.490000 104.065000 ;
      RECT 33.530000 171.345000 41.255000 171.495000 ;
      RECT 33.530000 171.345000 41.255000 171.495000 ;
      RECT 33.590000 103.765000 37.490000 103.915000 ;
      RECT 33.590000 103.765000 37.490000 103.915000 ;
      RECT 33.680000 171.495000 41.105000 171.645000 ;
      RECT 33.680000 171.495000 41.105000 171.645000 ;
      RECT 33.740000 103.615000 37.490000 103.765000 ;
      RECT 33.740000 103.615000 37.490000 103.765000 ;
      RECT 33.830000 171.645000 40.955000 171.795000 ;
      RECT 33.830000 171.645000 40.955000 171.795000 ;
      RECT 33.890000 103.465000 37.490000 103.615000 ;
      RECT 33.890000 103.465000 37.490000 103.615000 ;
      RECT 33.980000 171.795000 40.805000 171.945000 ;
      RECT 33.980000 171.795000 40.805000 171.945000 ;
      RECT 34.040000 103.315000 37.490000 103.465000 ;
      RECT 34.040000 103.315000 37.490000 103.465000 ;
      RECT 34.130000 171.945000 40.655000 172.095000 ;
      RECT 34.130000 171.945000 40.655000 172.095000 ;
      RECT 34.190000 103.165000 37.490000 103.315000 ;
      RECT 34.190000 103.165000 37.490000 103.315000 ;
      RECT 34.280000 172.095000 40.505000 172.245000 ;
      RECT 34.280000 172.095000 40.505000 172.245000 ;
      RECT 34.340000 103.015000 37.490000 103.165000 ;
      RECT 34.340000 103.015000 37.490000 103.165000 ;
      RECT 34.430000 172.245000 40.355000 172.395000 ;
      RECT 34.430000 172.245000 40.355000 172.395000 ;
      RECT 34.490000 102.865000 37.490000 103.015000 ;
      RECT 34.490000 102.865000 37.490000 103.015000 ;
      RECT 34.580000 172.395000 40.205000 172.545000 ;
      RECT 34.580000 172.395000 40.205000 172.545000 ;
      RECT 34.640000 102.715000 37.490000 102.865000 ;
      RECT 34.640000 102.715000 37.490000 102.865000 ;
      RECT 34.730000 172.545000 40.055000 172.695000 ;
      RECT 34.730000 172.545000 40.055000 172.695000 ;
      RECT 34.790000 102.565000 37.490000 102.715000 ;
      RECT 34.790000 102.565000 37.490000 102.715000 ;
      RECT 34.880000 172.695000 39.905000 172.845000 ;
      RECT 34.880000 172.695000 39.905000 172.845000 ;
      RECT 34.940000 102.415000 37.490000 102.565000 ;
      RECT 34.940000 102.415000 37.490000 102.565000 ;
      RECT 35.030000 172.845000 39.755000 172.995000 ;
      RECT 35.030000 172.845000 39.755000 172.995000 ;
      RECT 35.090000 102.265000 37.490000 102.415000 ;
      RECT 35.090000 102.265000 37.490000 102.415000 ;
      RECT 35.180000 172.995000 39.605000 173.145000 ;
      RECT 35.180000 172.995000 39.605000 173.145000 ;
      RECT 35.240000 102.115000 37.490000 102.265000 ;
      RECT 35.240000 102.115000 37.490000 102.265000 ;
      RECT 35.330000 173.145000 39.455000 173.295000 ;
      RECT 35.330000 173.145000 39.455000 173.295000 ;
      RECT 35.390000 101.965000 37.490000 102.115000 ;
      RECT 35.390000 101.965000 37.490000 102.115000 ;
      RECT 35.480000 173.295000 39.305000 173.445000 ;
      RECT 35.480000 173.295000 39.305000 173.445000 ;
      RECT 35.540000 101.815000 37.490000 101.965000 ;
      RECT 35.540000 101.815000 37.490000 101.965000 ;
      RECT 35.630000 173.445000 39.155000 173.595000 ;
      RECT 35.630000 173.445000 39.155000 173.595000 ;
      RECT 35.690000 101.665000 37.490000 101.815000 ;
      RECT 35.690000 101.665000 37.490000 101.815000 ;
      RECT 35.780000 173.595000 39.005000 173.745000 ;
      RECT 35.780000 173.595000 39.005000 173.745000 ;
      RECT 35.840000 101.515000 37.490000 101.665000 ;
      RECT 35.840000 101.515000 37.490000 101.665000 ;
      RECT 35.930000 173.745000 38.855000 173.895000 ;
      RECT 35.930000 173.745000 38.855000 173.895000 ;
      RECT 35.990000 101.365000 37.490000 101.515000 ;
      RECT 35.990000 101.365000 37.490000 101.515000 ;
      RECT 36.080000 173.895000 38.705000 174.045000 ;
      RECT 36.080000 173.895000 38.705000 174.045000 ;
      RECT 36.140000 101.215000 37.490000 101.365000 ;
      RECT 36.140000 101.215000 37.490000 101.365000 ;
      RECT 36.230000 174.045000 38.555000 174.195000 ;
      RECT 36.230000 174.045000 38.555000 174.195000 ;
      RECT 36.290000 101.065000 37.490000 101.215000 ;
      RECT 36.290000 101.065000 37.490000 101.215000 ;
      RECT 36.380000 174.195000 38.405000 174.345000 ;
      RECT 36.380000 174.195000 38.405000 174.345000 ;
      RECT 36.440000 100.915000 37.490000 101.065000 ;
      RECT 36.440000 100.915000 37.490000 101.065000 ;
      RECT 36.530000 174.345000 38.255000 174.495000 ;
      RECT 36.530000 174.345000 38.255000 174.495000 ;
      RECT 36.590000 100.765000 37.490000 100.915000 ;
      RECT 36.590000 100.765000 37.490000 100.915000 ;
      RECT 36.680000 174.495000 38.105000 174.645000 ;
      RECT 36.680000 174.495000 38.105000 174.645000 ;
      RECT 36.740000 100.615000 37.490000 100.765000 ;
      RECT 36.740000 100.615000 37.490000 100.765000 ;
      RECT 36.830000 174.645000 37.955000 174.795000 ;
      RECT 36.830000 174.645000 37.955000 174.795000 ;
      RECT 36.890000 100.465000 37.490000 100.615000 ;
      RECT 36.890000 100.465000 37.490000 100.615000 ;
      RECT 36.980000 174.795000 37.805000 174.945000 ;
      RECT 36.980000 174.795000 37.805000 174.945000 ;
      RECT 37.040000 100.315000 37.490000 100.465000 ;
      RECT 37.040000 100.315000 37.490000 100.465000 ;
      RECT 37.130000 174.945000 37.655000 175.095000 ;
      RECT 37.130000 174.945000 37.655000 175.095000 ;
      RECT 37.190000 100.165000 37.490000 100.315000 ;
      RECT 37.190000 100.165000 37.490000 100.315000 ;
      RECT 37.220000 175.185000 37.565000 190.420000 ;
      RECT 37.220000 175.270000 37.305000 175.355000 ;
      RECT 37.220000 175.355000 37.565000 190.420000 ;
      RECT 37.220000 190.420000 49.375000 190.440000 ;
      RECT 37.220000 190.420000 49.375000 190.440000 ;
      RECT 37.220000 190.420000 49.375000 200.000000 ;
      RECT 37.220000 190.440000 75.000000 195.500000 ;
      RECT 37.220000 190.440000 75.000000 195.500000 ;
      RECT 37.220000 190.440000 75.000000 200.000000 ;
      RECT 37.280000 175.095000 37.505000 175.245000 ;
      RECT 37.280000 175.095000 37.505000 175.245000 ;
      RECT 37.295000   0.000000 37.490000 100.060000 ;
      RECT 37.295000 100.060000 37.490000 105.025000 ;
      RECT 37.340000 100.015000 37.490000 100.165000 ;
      RECT 37.340000 100.015000 37.490000 100.165000 ;
      RECT 37.390000 175.245000 37.395000 175.355000 ;
      RECT 37.390000 175.245000 37.395000 175.355000 ;
      RECT 37.480000 175.270000 37.565000 175.355000 ;
      RECT 43.240000 100.380000 44.860000 101.970000 ;
      RECT 43.240000 100.380000 44.860000 101.970000 ;
      RECT 43.240000 101.970000 44.860000 102.580000 ;
      RECT 43.265000 100.355000 44.835000 100.380000 ;
      RECT 43.390000 101.970000 44.860000 102.120000 ;
      RECT 43.415000 100.205000 44.685000 100.355000 ;
      RECT 43.540000 102.120000 44.860000 102.270000 ;
      RECT 43.565000 100.055000 44.535000 100.205000 ;
      RECT 43.690000 102.270000 44.860000 102.420000 ;
      RECT 43.715000  99.905000 44.385000 100.055000 ;
      RECT 43.715000  99.905000 44.860000 100.380000 ;
      RECT 43.840000 102.420000 44.860000 102.570000 ;
      RECT 43.850000 102.570000 44.860000 102.580000 ;
      RECT 43.850000 102.580000 50.265000 107.985000 ;
      RECT 44.000000 102.580000 44.860000 102.730000 ;
      RECT 44.150000 102.730000 45.010000 102.880000 ;
      RECT 44.300000 102.880000 45.160000 103.030000 ;
      RECT 44.450000 103.030000 45.310000 103.180000 ;
      RECT 44.600000 103.180000 45.460000 103.330000 ;
      RECT 44.750000 103.330000 45.610000 103.480000 ;
      RECT 44.900000 103.480000 45.760000 103.630000 ;
      RECT 45.050000 103.630000 45.910000 103.780000 ;
      RECT 45.200000 103.780000 46.060000 103.930000 ;
      RECT 45.350000 103.930000 46.210000 104.080000 ;
      RECT 45.500000 104.080000 46.360000 104.230000 ;
      RECT 45.650000 104.230000 46.510000 104.380000 ;
      RECT 45.800000 104.380000 46.660000 104.530000 ;
      RECT 45.950000 104.530000 46.810000 104.680000 ;
      RECT 46.100000 104.680000 46.960000 104.830000 ;
      RECT 46.250000 104.830000 47.110000 104.980000 ;
      RECT 46.400000 104.980000 47.260000 105.130000 ;
      RECT 46.550000 105.130000 47.410000 105.280000 ;
      RECT 46.700000 105.280000 47.560000 105.430000 ;
      RECT 46.850000 105.430000 47.710000 105.580000 ;
      RECT 47.000000 105.580000 47.860000 105.730000 ;
      RECT 47.150000 105.730000 48.010000 105.880000 ;
      RECT 47.300000 105.880000 48.160000 106.030000 ;
      RECT 47.450000 106.030000 48.310000 106.180000 ;
      RECT 47.600000 106.180000 48.460000 106.330000 ;
      RECT 47.750000 106.330000 48.610000 106.480000 ;
      RECT 47.900000 106.480000 48.760000 106.630000 ;
      RECT 48.050000 106.630000 48.910000 106.780000 ;
      RECT 48.200000 106.780000 49.060000 106.930000 ;
      RECT 48.350000 106.930000 49.210000 107.080000 ;
      RECT 48.500000 107.080000 49.360000 107.230000 ;
      RECT 48.650000 107.230000 49.510000 107.380000 ;
      RECT 48.800000 107.380000 49.660000 107.530000 ;
      RECT 48.950000 107.530000 49.810000 107.680000 ;
      RECT 49.100000 107.680000 49.960000 107.830000 ;
      RECT 49.250000 107.830000 50.110000 107.980000 ;
      RECT 49.255000 107.980000 50.260000 107.985000 ;
      RECT 49.255000 107.985000 50.265000 108.135000 ;
      RECT 49.255000 107.985000 52.885000 110.605000 ;
      RECT 49.255000 108.135000 50.415000 108.285000 ;
      RECT 49.255000 108.285000 50.565000 108.435000 ;
      RECT 49.255000 108.435000 50.715000 108.585000 ;
      RECT 49.255000 108.585000 50.865000 108.735000 ;
      RECT 49.255000 108.735000 51.015000 108.885000 ;
      RECT 49.255000 108.885000 51.165000 109.035000 ;
      RECT 49.255000 109.035000 51.315000 109.185000 ;
      RECT 49.255000 109.185000 51.465000 109.335000 ;
      RECT 49.255000 109.335000 51.615000 109.485000 ;
      RECT 49.255000 109.485000 51.765000 109.635000 ;
      RECT 49.255000 109.635000 51.915000 109.785000 ;
      RECT 49.255000 109.785000 52.065000 109.935000 ;
      RECT 49.255000 109.935000 52.215000 110.085000 ;
      RECT 49.255000 110.085000 52.365000 110.235000 ;
      RECT 49.255000 110.235000 52.515000 110.385000 ;
      RECT 49.255000 110.385000 52.665000 110.535000 ;
      RECT 49.255000 110.535000 52.815000 110.605000 ;
      RECT 49.255000 110.605000 52.885000 168.970000 ;
      RECT 49.255000 110.605000 52.885000 168.970000 ;
      RECT 49.255000 168.970000 49.375000 172.480000 ;
      RECT 49.255000 168.970000 52.735000 169.120000 ;
      RECT 49.255000 169.120000 52.585000 169.270000 ;
      RECT 49.255000 169.270000 52.435000 169.420000 ;
      RECT 49.255000 169.420000 52.285000 169.570000 ;
      RECT 49.255000 169.570000 52.135000 169.720000 ;
      RECT 49.255000 169.720000 51.985000 169.870000 ;
      RECT 49.255000 169.870000 51.835000 170.020000 ;
      RECT 49.255000 170.020000 51.685000 170.170000 ;
      RECT 49.255000 170.170000 51.535000 170.320000 ;
      RECT 49.255000 170.320000 51.385000 170.470000 ;
      RECT 49.255000 170.470000 51.235000 170.620000 ;
      RECT 49.255000 170.620000 51.085000 170.770000 ;
      RECT 49.255000 170.770000 50.935000 170.920000 ;
      RECT 49.255000 170.920000 50.785000 171.070000 ;
      RECT 49.255000 171.070000 50.635000 171.220000 ;
      RECT 49.255000 171.220000 50.485000 171.370000 ;
      RECT 49.255000 171.370000 50.335000 171.520000 ;
      RECT 49.255000 171.520000 50.185000 171.670000 ;
      RECT 49.255000 171.670000 50.035000 171.820000 ;
      RECT 49.255000 171.820000 49.885000 171.970000 ;
      RECT 49.255000 171.970000 49.735000 172.120000 ;
      RECT 49.255000 172.120000 49.585000 172.270000 ;
      RECT 49.255000 172.270000 49.435000 172.420000 ;
      RECT 49.255000 172.420000 49.285000 172.570000 ;
      RECT 49.255000 172.480000 49.375000 190.420000 ;
      RECT 49.290000   0.000000 49.990000  89.650000 ;
      RECT 49.290000   0.000000 50.090000  90.310000 ;
      RECT 49.290000  89.800000 49.440000  89.950000 ;
      RECT 49.290000  89.800000 49.440000  89.950000 ;
      RECT 49.290000  89.950000 49.590000  90.100000 ;
      RECT 49.290000  89.950000 49.590000  90.100000 ;
      RECT 49.290000  90.100000 49.740000  90.250000 ;
      RECT 49.290000  90.100000 49.740000  90.250000 ;
      RECT 49.290000  90.250000 49.890000  90.400000 ;
      RECT 49.290000  90.250000 49.890000  90.400000 ;
      RECT 49.290000  90.310000 55.765000  95.985000 ;
      RECT 49.290000  90.400000 50.040000  90.550000 ;
      RECT 49.290000  90.400000 50.040000  90.550000 ;
      RECT 49.290000  90.550000 50.190000  90.700000 ;
      RECT 49.290000  90.550000 50.190000  90.700000 ;
      RECT 49.290000  90.700000 50.340000  90.850000 ;
      RECT 49.290000  90.700000 50.340000  90.850000 ;
      RECT 49.290000  90.850000 50.490000  91.000000 ;
      RECT 49.290000  90.850000 50.490000  91.000000 ;
      RECT 49.290000  91.000000 50.640000  91.150000 ;
      RECT 49.290000  91.000000 50.640000  91.150000 ;
      RECT 49.290000  91.150000 50.790000  91.300000 ;
      RECT 49.290000  91.150000 50.790000  91.300000 ;
      RECT 49.290000  91.300000 50.940000  91.450000 ;
      RECT 49.290000  91.300000 50.940000  91.450000 ;
      RECT 49.290000  91.450000 51.090000  91.600000 ;
      RECT 49.290000  91.450000 51.090000  91.600000 ;
      RECT 49.290000  91.600000 51.240000  91.750000 ;
      RECT 49.290000  91.600000 51.240000  91.750000 ;
      RECT 49.290000  91.750000 51.390000  91.900000 ;
      RECT 49.290000  91.750000 51.390000  91.900000 ;
      RECT 49.290000  91.900000 51.540000  92.050000 ;
      RECT 49.290000  91.900000 51.540000  92.050000 ;
      RECT 49.290000  92.050000 51.690000  92.200000 ;
      RECT 49.290000  92.050000 51.690000  92.200000 ;
      RECT 49.290000  92.200000 51.840000  92.350000 ;
      RECT 49.290000  92.200000 51.840000  92.350000 ;
      RECT 49.290000  92.350000 51.990000  92.500000 ;
      RECT 49.290000  92.350000 51.990000  92.500000 ;
      RECT 49.290000  92.500000 52.140000  92.650000 ;
      RECT 49.290000  92.500000 52.140000  92.650000 ;
      RECT 49.290000  92.650000 52.290000  92.800000 ;
      RECT 49.290000  92.650000 52.290000  92.800000 ;
      RECT 49.290000  92.800000 52.440000  92.950000 ;
      RECT 49.290000  92.800000 52.440000  92.950000 ;
      RECT 49.290000  92.950000 52.590000  93.100000 ;
      RECT 49.290000  92.950000 52.590000  93.100000 ;
      RECT 49.290000  93.100000 52.740000  93.250000 ;
      RECT 49.290000  93.100000 52.740000  93.250000 ;
      RECT 49.290000  93.250000 52.890000  93.400000 ;
      RECT 49.290000  93.250000 52.890000  93.400000 ;
      RECT 49.290000  93.400000 53.040000  93.550000 ;
      RECT 49.290000  93.400000 53.040000  93.550000 ;
      RECT 49.290000  93.550000 53.190000  93.700000 ;
      RECT 49.290000  93.550000 53.190000  93.700000 ;
      RECT 49.290000  93.700000 53.340000  93.850000 ;
      RECT 49.290000  93.700000 53.340000  93.850000 ;
      RECT 49.290000  93.850000 53.490000  94.000000 ;
      RECT 49.290000  93.850000 53.490000  94.000000 ;
      RECT 49.290000  94.000000 53.640000  94.150000 ;
      RECT 49.290000  94.000000 53.640000  94.150000 ;
      RECT 49.290000  94.150000 53.790000  94.300000 ;
      RECT 49.290000  94.150000 53.790000  94.300000 ;
      RECT 49.290000  94.300000 53.940000  94.450000 ;
      RECT 49.290000  94.300000 53.940000  94.450000 ;
      RECT 49.290000  94.450000 54.090000  94.600000 ;
      RECT 49.290000  94.450000 54.090000  94.600000 ;
      RECT 49.290000  94.600000 54.240000  94.750000 ;
      RECT 49.290000  94.600000 54.240000  94.750000 ;
      RECT 49.290000  94.750000 54.390000  94.900000 ;
      RECT 49.290000  94.750000 54.390000  94.900000 ;
      RECT 49.290000  94.900000 54.540000  95.050000 ;
      RECT 49.290000  94.900000 54.540000  95.050000 ;
      RECT 49.290000  95.050000 54.690000  95.200000 ;
      RECT 49.290000  95.050000 54.690000  95.200000 ;
      RECT 49.290000  95.200000 54.840000  95.350000 ;
      RECT 49.290000  95.200000 54.840000  95.350000 ;
      RECT 49.290000  95.350000 54.990000  95.500000 ;
      RECT 49.290000  95.350000 54.990000  95.500000 ;
      RECT 49.290000  95.500000 55.140000  95.650000 ;
      RECT 49.290000  95.500000 55.140000  95.650000 ;
      RECT 49.290000  95.650000 55.290000  95.800000 ;
      RECT 49.290000  95.650000 55.290000  95.800000 ;
      RECT 49.290000  95.800000 55.440000  95.950000 ;
      RECT 49.290000  95.800000 55.440000  95.950000 ;
      RECT 49.290000  95.950000 55.590000  95.985000 ;
      RECT 49.290000  95.950000 55.590000  95.985000 ;
      RECT 49.290000  95.985000 57.915000  98.135000 ;
      RECT 49.440000  95.985000 55.625000  96.135000 ;
      RECT 49.440000  95.985000 55.625000  96.135000 ;
      RECT 49.590000  96.135000 55.775000  96.285000 ;
      RECT 49.590000  96.135000 55.775000  96.285000 ;
      RECT 49.740000  96.285000 55.925000  96.435000 ;
      RECT 49.740000  96.285000 55.925000  96.435000 ;
      RECT 49.890000  96.435000 56.075000  96.585000 ;
      RECT 49.890000  96.435000 56.075000  96.585000 ;
      RECT 50.040000  96.585000 56.225000  96.735000 ;
      RECT 50.040000  96.585000 56.225000  96.735000 ;
      RECT 50.190000  96.735000 56.375000  96.885000 ;
      RECT 50.190000  96.735000 56.375000  96.885000 ;
      RECT 50.340000  96.885000 56.525000  97.035000 ;
      RECT 50.340000  96.885000 56.525000  97.035000 ;
      RECT 50.490000  97.035000 56.675000  97.185000 ;
      RECT 50.490000  97.035000 56.675000  97.185000 ;
      RECT 50.640000  97.185000 56.825000  97.335000 ;
      RECT 50.640000  97.185000 56.825000  97.335000 ;
      RECT 50.790000  97.335000 56.975000  97.485000 ;
      RECT 50.790000  97.335000 56.975000  97.485000 ;
      RECT 50.940000  97.485000 57.125000  97.635000 ;
      RECT 50.940000  97.485000 57.125000  97.635000 ;
      RECT 51.090000  97.635000 57.275000  97.785000 ;
      RECT 51.090000  97.635000 57.275000  97.785000 ;
      RECT 51.240000  97.785000 57.425000  97.935000 ;
      RECT 51.240000  97.785000 57.425000  97.935000 ;
      RECT 51.390000  97.935000 57.575000  98.085000 ;
      RECT 51.390000  97.935000 57.575000  98.085000 ;
      RECT 51.440000  98.085000 57.725000  98.135000 ;
      RECT 51.440000  98.085000 57.725000  98.135000 ;
      RECT 51.440000  98.135000 57.775000  98.285000 ;
      RECT 51.440000  98.135000 57.775000  98.285000 ;
      RECT 51.440000  98.135000 59.330000  99.550000 ;
      RECT 51.440000  98.285000 57.925000  98.435000 ;
      RECT 51.440000  98.285000 57.925000  98.435000 ;
      RECT 51.440000  98.435000 58.075000  98.585000 ;
      RECT 51.440000  98.435000 58.075000  98.585000 ;
      RECT 51.440000  98.585000 58.225000  98.735000 ;
      RECT 51.440000  98.585000 58.225000  98.735000 ;
      RECT 51.440000  98.735000 58.375000  98.885000 ;
      RECT 51.440000  98.735000 58.375000  98.885000 ;
      RECT 51.440000  98.885000 58.525000  99.035000 ;
      RECT 51.440000  98.885000 58.525000  99.035000 ;
      RECT 51.440000  99.035000 58.675000  99.185000 ;
      RECT 51.440000  99.035000 58.675000  99.185000 ;
      RECT 51.440000  99.185000 58.825000  99.335000 ;
      RECT 51.440000  99.185000 58.825000  99.335000 ;
      RECT 51.440000  99.335000 58.975000  99.485000 ;
      RECT 51.440000  99.335000 58.975000  99.485000 ;
      RECT 51.440000  99.485000 59.125000  99.550000 ;
      RECT 51.440000  99.485000 59.125000  99.550000 ;
      RECT 51.440000  99.550000 61.200000 101.420000 ;
      RECT 51.590000  99.550000 59.190000  99.700000 ;
      RECT 51.590000  99.550000 59.190000  99.700000 ;
      RECT 51.740000  99.700000 59.340000  99.850000 ;
      RECT 51.740000  99.700000 59.340000  99.850000 ;
      RECT 51.890000  99.850000 59.490000 100.000000 ;
      RECT 51.890000  99.850000 59.490000 100.000000 ;
      RECT 52.040000 100.000000 59.640000 100.150000 ;
      RECT 52.040000 100.000000 59.640000 100.150000 ;
      RECT 52.190000 100.150000 59.790000 100.300000 ;
      RECT 52.190000 100.150000 59.790000 100.300000 ;
      RECT 52.340000 100.300000 59.940000 100.450000 ;
      RECT 52.340000 100.300000 59.940000 100.450000 ;
      RECT 52.490000 100.450000 60.090000 100.600000 ;
      RECT 52.490000 100.450000 60.090000 100.600000 ;
      RECT 52.640000 100.600000 60.240000 100.750000 ;
      RECT 52.640000 100.600000 60.240000 100.750000 ;
      RECT 52.790000 100.750000 60.390000 100.900000 ;
      RECT 52.790000 100.750000 60.390000 100.900000 ;
      RECT 52.940000 100.900000 60.540000 101.050000 ;
      RECT 52.940000 100.900000 60.540000 101.050000 ;
      RECT 53.090000 101.050000 60.690000 101.200000 ;
      RECT 53.090000 101.050000 60.690000 101.200000 ;
      RECT 53.240000 101.200000 60.840000 101.350000 ;
      RECT 53.240000 101.200000 60.840000 101.350000 ;
      RECT 53.310000 101.420000 61.200000 107.795000 ;
      RECT 53.350000 101.350000 60.990000 101.460000 ;
      RECT 53.350000 101.350000 60.990000 101.460000 ;
      RECT 53.500000 101.460000 61.100000 101.610000 ;
      RECT 53.500000 101.460000 61.100000 101.610000 ;
      RECT 53.650000 101.610000 61.100000 101.760000 ;
      RECT 53.650000 101.610000 61.100000 101.760000 ;
      RECT 53.800000 101.760000 61.100000 101.910000 ;
      RECT 53.800000 101.760000 61.100000 101.910000 ;
      RECT 53.950000 101.910000 61.100000 102.060000 ;
      RECT 53.950000 101.910000 61.100000 102.060000 ;
      RECT 54.100000 102.060000 61.100000 102.210000 ;
      RECT 54.100000 102.060000 61.100000 102.210000 ;
      RECT 54.250000 102.210000 61.100000 102.360000 ;
      RECT 54.250000 102.210000 61.100000 102.360000 ;
      RECT 54.400000 102.360000 61.100000 102.510000 ;
      RECT 54.400000 102.360000 61.100000 102.510000 ;
      RECT 54.550000 102.510000 61.100000 102.660000 ;
      RECT 54.550000 102.510000 61.100000 102.660000 ;
      RECT 54.700000 102.660000 61.100000 102.810000 ;
      RECT 54.700000 102.660000 61.100000 102.810000 ;
      RECT 54.850000 102.810000 61.100000 102.960000 ;
      RECT 54.850000 102.810000 61.100000 102.960000 ;
      RECT 55.000000 102.960000 61.100000 103.110000 ;
      RECT 55.000000 102.960000 61.100000 103.110000 ;
      RECT 55.150000 103.110000 61.100000 103.260000 ;
      RECT 55.150000 103.110000 61.100000 103.260000 ;
      RECT 55.300000 103.260000 61.100000 103.410000 ;
      RECT 55.300000 103.260000 61.100000 103.410000 ;
      RECT 55.450000 103.410000 61.100000 103.560000 ;
      RECT 55.450000 103.410000 61.100000 103.560000 ;
      RECT 55.600000 103.560000 61.100000 103.710000 ;
      RECT 55.600000 103.560000 61.100000 103.710000 ;
      RECT 55.750000 103.710000 61.100000 103.860000 ;
      RECT 55.750000 103.710000 61.100000 103.860000 ;
      RECT 55.900000 103.860000 61.100000 104.010000 ;
      RECT 55.900000 103.860000 61.100000 104.010000 ;
      RECT 56.050000 104.010000 61.100000 104.160000 ;
      RECT 56.050000 104.010000 61.100000 104.160000 ;
      RECT 56.200000 104.160000 61.100000 104.310000 ;
      RECT 56.200000 104.160000 61.100000 104.310000 ;
      RECT 56.350000 104.310000 61.100000 104.460000 ;
      RECT 56.350000 104.310000 61.100000 104.460000 ;
      RECT 56.500000 104.460000 61.100000 104.610000 ;
      RECT 56.500000 104.460000 61.100000 104.610000 ;
      RECT 56.650000 104.610000 61.100000 104.760000 ;
      RECT 56.650000 104.610000 61.100000 104.760000 ;
      RECT 56.800000 104.760000 61.100000 104.910000 ;
      RECT 56.800000 104.760000 61.100000 104.910000 ;
      RECT 56.950000 104.910000 61.100000 105.060000 ;
      RECT 56.950000 104.910000 61.100000 105.060000 ;
      RECT 57.100000 105.060000 61.100000 105.210000 ;
      RECT 57.100000 105.060000 61.100000 105.210000 ;
      RECT 57.250000 105.210000 61.100000 105.360000 ;
      RECT 57.250000 105.210000 61.100000 105.360000 ;
      RECT 57.400000 105.360000 61.100000 105.510000 ;
      RECT 57.400000 105.360000 61.100000 105.510000 ;
      RECT 57.550000 105.510000 61.100000 105.660000 ;
      RECT 57.550000 105.510000 61.100000 105.660000 ;
      RECT 57.700000 105.660000 61.100000 105.810000 ;
      RECT 57.700000 105.660000 61.100000 105.810000 ;
      RECT 57.850000 105.810000 61.100000 105.960000 ;
      RECT 57.850000 105.810000 61.100000 105.960000 ;
      RECT 58.000000 105.960000 61.100000 106.110000 ;
      RECT 58.000000 105.960000 61.100000 106.110000 ;
      RECT 58.150000 106.110000 61.100000 106.260000 ;
      RECT 58.150000 106.110000 61.100000 106.260000 ;
      RECT 58.300000 106.260000 61.100000 106.410000 ;
      RECT 58.300000 106.260000 61.100000 106.410000 ;
      RECT 58.450000 106.410000 61.100000 106.560000 ;
      RECT 58.450000 106.410000 61.100000 106.560000 ;
      RECT 58.600000 106.560000 61.100000 106.710000 ;
      RECT 58.600000 106.560000 61.100000 106.710000 ;
      RECT 58.750000 106.710000 61.100000 106.860000 ;
      RECT 58.750000 106.710000 61.100000 106.860000 ;
      RECT 58.900000 106.860000 61.100000 107.010000 ;
      RECT 58.900000 106.860000 61.100000 107.010000 ;
      RECT 59.050000 107.010000 61.100000 107.160000 ;
      RECT 59.050000 107.010000 61.100000 107.160000 ;
      RECT 59.200000 107.160000 61.100000 107.310000 ;
      RECT 59.200000 107.160000 61.100000 107.310000 ;
      RECT 59.350000 107.310000 61.100000 107.460000 ;
      RECT 59.350000 107.310000 61.100000 107.460000 ;
      RECT 59.500000 107.460000 61.100000 107.610000 ;
      RECT 59.500000 107.460000 61.100000 107.610000 ;
      RECT 59.650000 107.610000 61.100000 107.760000 ;
      RECT 59.650000 107.610000 61.100000 107.760000 ;
      RECT 59.685000 107.795000 61.200000 172.855000 ;
      RECT 59.685000 107.945000 59.835000 108.095000 ;
      RECT 59.685000 108.095000 59.985000 108.245000 ;
      RECT 59.685000 108.245000 60.135000 108.395000 ;
      RECT 59.685000 108.395000 60.285000 108.545000 ;
      RECT 59.685000 108.545000 60.435000 108.695000 ;
      RECT 59.685000 108.695000 60.585000 108.845000 ;
      RECT 59.685000 108.845000 60.735000 108.995000 ;
      RECT 59.685000 108.995000 60.885000 109.145000 ;
      RECT 59.685000 109.145000 61.035000 109.210000 ;
      RECT 59.685000 109.210000 61.100000 172.855000 ;
      RECT 59.685000 172.855000 61.200000 173.620000 ;
      RECT 59.800000 107.760000 61.100000 107.910000 ;
      RECT 59.800000 107.760000 61.100000 107.910000 ;
      RECT 59.835000 172.855000 61.100000 173.005000 ;
      RECT 59.950000 107.910000 61.100000 108.060000 ;
      RECT 59.950000 107.910000 61.100000 108.060000 ;
      RECT 59.985000 173.005000 61.100000 173.155000 ;
      RECT 60.100000 108.060000 61.100000 108.210000 ;
      RECT 60.100000 108.060000 61.100000 108.210000 ;
      RECT 60.135000 173.155000 61.100000 173.305000 ;
      RECT 60.250000 108.210000 61.100000 108.360000 ;
      RECT 60.250000 108.210000 61.100000 108.360000 ;
      RECT 60.285000 173.305000 61.100000 173.455000 ;
      RECT 60.400000 108.360000 61.100000 108.510000 ;
      RECT 60.400000 108.360000 61.100000 108.510000 ;
      RECT 60.435000 173.455000 61.100000 173.605000 ;
      RECT 60.450000 173.620000 75.000000 174.515000 ;
      RECT 60.550000 108.510000 61.100000 108.660000 ;
      RECT 60.550000 108.510000 61.100000 108.660000 ;
      RECT 60.550000 173.605000 61.100000 173.720000 ;
      RECT 60.700000 108.660000 61.100000 108.810000 ;
      RECT 60.700000 108.660000 61.100000 108.810000 ;
      RECT 60.700000 173.720000 75.000000 173.870000 ;
      RECT 60.850000 108.810000 61.100000 108.960000 ;
      RECT 60.850000 108.810000 61.100000 108.960000 ;
      RECT 60.850000 173.870000 75.000000 174.020000 ;
      RECT 61.000000 108.960000 61.100000 109.110000 ;
      RECT 61.000000 108.960000 61.100000 109.110000 ;
      RECT 61.000000 174.020000 75.000000 174.170000 ;
      RECT 61.150000 174.170000 75.000000 174.320000 ;
      RECT 61.300000 174.320000 75.000000 174.470000 ;
      RECT 61.345000 173.720000 75.000000 190.440000 ;
      RECT 61.345000 173.720000 75.000000 200.000000 ;
      RECT 61.345000 174.470000 75.000000 174.515000 ;
      RECT 61.345000 174.515000 75.000000 190.440000 ;
      RECT 74.590000   0.000000 75.000000 173.620000 ;
      RECT 74.690000   0.000000 75.000000 173.720000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   0.000000 75.000000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000   7.885000 75.000000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  13.935000 75.000000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  18.785000 75.000000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  24.835000 75.000000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  30.885000 75.000000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  35.735000 75.000000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  40.585000 75.000000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  46.635000 75.000000  47.435000 ;
      RECT  0.000000  57.035000 75.000000  57.835000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  63.085000 75.000000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  68.935000 75.000000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.570000  47.435000 73.430000  57.035000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000  19.385000 73.330000  95.400000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000 75.000000   0.535000 ;
      RECT  0.000000  96.585000 75.000000 137.725000 ;
      RECT  0.000000 137.725000 35.045000 147.535000 ;
      RECT  0.000000 147.535000 75.000000 174.185000 ;
      RECT  2.565000  15.035000 72.435000  18.285000 ;
      RECT  2.870000   0.000000 72.130000  15.035000 ;
      RECT  2.870000  18.285000 72.130000  96.585000 ;
      RECT  2.870000 174.185000 72.130000 200.000000 ;
      RECT 39.570000 137.725000 75.000000 147.535000 ;
  END
END sky130_fd_io__top_ground_hvc_wpad


MACRO sky130_fd_io__overlay_vccd_lvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.600000 6.890000 24.500000 11.530000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 6.890000 74.655000 11.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 24.475000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.690000  6.960000  0.890000  7.160000 ;
        RECT  0.690000  7.390000  0.890000  7.590000 ;
        RECT  0.690000  7.820000  0.890000  8.020000 ;
        RECT  0.690000  8.250000  0.890000  8.450000 ;
        RECT  0.690000  8.680000  0.890000  8.880000 ;
        RECT  0.690000  9.110000  0.890000  9.310000 ;
        RECT  0.690000  9.540000  0.890000  9.740000 ;
        RECT  0.690000  9.970000  0.890000 10.170000 ;
        RECT  0.690000 10.400000  0.890000 10.600000 ;
        RECT  0.690000 10.830000  0.890000 11.030000 ;
        RECT  0.690000 11.260000  0.890000 11.460000 ;
        RECT  1.100000  6.960000  1.300000  7.160000 ;
        RECT  1.100000  7.390000  1.300000  7.590000 ;
        RECT  1.100000  7.820000  1.300000  8.020000 ;
        RECT  1.100000  8.250000  1.300000  8.450000 ;
        RECT  1.100000  8.680000  1.300000  8.880000 ;
        RECT  1.100000  9.110000  1.300000  9.310000 ;
        RECT  1.100000  9.540000  1.300000  9.740000 ;
        RECT  1.100000  9.970000  1.300000 10.170000 ;
        RECT  1.100000 10.400000  1.300000 10.600000 ;
        RECT  1.100000 10.830000  1.300000 11.030000 ;
        RECT  1.100000 11.260000  1.300000 11.460000 ;
        RECT  1.510000  6.960000  1.710000  7.160000 ;
        RECT  1.510000  7.390000  1.710000  7.590000 ;
        RECT  1.510000  7.820000  1.710000  8.020000 ;
        RECT  1.510000  8.250000  1.710000  8.450000 ;
        RECT  1.510000  8.680000  1.710000  8.880000 ;
        RECT  1.510000  9.110000  1.710000  9.310000 ;
        RECT  1.510000  9.540000  1.710000  9.740000 ;
        RECT  1.510000  9.970000  1.710000 10.170000 ;
        RECT  1.510000 10.400000  1.710000 10.600000 ;
        RECT  1.510000 10.830000  1.710000 11.030000 ;
        RECT  1.510000 11.260000  1.710000 11.460000 ;
        RECT  1.920000  6.960000  2.120000  7.160000 ;
        RECT  1.920000  7.390000  2.120000  7.590000 ;
        RECT  1.920000  7.820000  2.120000  8.020000 ;
        RECT  1.920000  8.250000  2.120000  8.450000 ;
        RECT  1.920000  8.680000  2.120000  8.880000 ;
        RECT  1.920000  9.110000  2.120000  9.310000 ;
        RECT  1.920000  9.540000  2.120000  9.740000 ;
        RECT  1.920000  9.970000  2.120000 10.170000 ;
        RECT  1.920000 10.400000  2.120000 10.600000 ;
        RECT  1.920000 10.830000  2.120000 11.030000 ;
        RECT  1.920000 11.260000  2.120000 11.460000 ;
        RECT  2.330000  6.960000  2.530000  7.160000 ;
        RECT  2.330000  7.390000  2.530000  7.590000 ;
        RECT  2.330000  7.820000  2.530000  8.020000 ;
        RECT  2.330000  8.250000  2.530000  8.450000 ;
        RECT  2.330000  8.680000  2.530000  8.880000 ;
        RECT  2.330000  9.110000  2.530000  9.310000 ;
        RECT  2.330000  9.540000  2.530000  9.740000 ;
        RECT  2.330000  9.970000  2.530000 10.170000 ;
        RECT  2.330000 10.400000  2.530000 10.600000 ;
        RECT  2.330000 10.830000  2.530000 11.030000 ;
        RECT  2.330000 11.260000  2.530000 11.460000 ;
        RECT  2.740000  6.960000  2.940000  7.160000 ;
        RECT  2.740000  7.390000  2.940000  7.590000 ;
        RECT  2.740000  7.820000  2.940000  8.020000 ;
        RECT  2.740000  8.250000  2.940000  8.450000 ;
        RECT  2.740000  8.680000  2.940000  8.880000 ;
        RECT  2.740000  9.110000  2.940000  9.310000 ;
        RECT  2.740000  9.540000  2.940000  9.740000 ;
        RECT  2.740000  9.970000  2.940000 10.170000 ;
        RECT  2.740000 10.400000  2.940000 10.600000 ;
        RECT  2.740000 10.830000  2.940000 11.030000 ;
        RECT  2.740000 11.260000  2.940000 11.460000 ;
        RECT  3.150000  6.960000  3.350000  7.160000 ;
        RECT  3.150000  7.390000  3.350000  7.590000 ;
        RECT  3.150000  7.820000  3.350000  8.020000 ;
        RECT  3.150000  8.250000  3.350000  8.450000 ;
        RECT  3.150000  8.680000  3.350000  8.880000 ;
        RECT  3.150000  9.110000  3.350000  9.310000 ;
        RECT  3.150000  9.540000  3.350000  9.740000 ;
        RECT  3.150000  9.970000  3.350000 10.170000 ;
        RECT  3.150000 10.400000  3.350000 10.600000 ;
        RECT  3.150000 10.830000  3.350000 11.030000 ;
        RECT  3.150000 11.260000  3.350000 11.460000 ;
        RECT  3.555000  6.960000  3.755000  7.160000 ;
        RECT  3.555000  7.390000  3.755000  7.590000 ;
        RECT  3.555000  7.820000  3.755000  8.020000 ;
        RECT  3.555000  8.250000  3.755000  8.450000 ;
        RECT  3.555000  8.680000  3.755000  8.880000 ;
        RECT  3.555000  9.110000  3.755000  9.310000 ;
        RECT  3.555000  9.540000  3.755000  9.740000 ;
        RECT  3.555000  9.970000  3.755000 10.170000 ;
        RECT  3.555000 10.400000  3.755000 10.600000 ;
        RECT  3.555000 10.830000  3.755000 11.030000 ;
        RECT  3.555000 11.260000  3.755000 11.460000 ;
        RECT  3.960000  6.960000  4.160000  7.160000 ;
        RECT  3.960000  7.390000  4.160000  7.590000 ;
        RECT  3.960000  7.820000  4.160000  8.020000 ;
        RECT  3.960000  8.250000  4.160000  8.450000 ;
        RECT  3.960000  8.680000  4.160000  8.880000 ;
        RECT  3.960000  9.110000  4.160000  9.310000 ;
        RECT  3.960000  9.540000  4.160000  9.740000 ;
        RECT  3.960000  9.970000  4.160000 10.170000 ;
        RECT  3.960000 10.400000  4.160000 10.600000 ;
        RECT  3.960000 10.830000  4.160000 11.030000 ;
        RECT  3.960000 11.260000  4.160000 11.460000 ;
        RECT  4.365000  6.960000  4.565000  7.160000 ;
        RECT  4.365000  7.390000  4.565000  7.590000 ;
        RECT  4.365000  7.820000  4.565000  8.020000 ;
        RECT  4.365000  8.250000  4.565000  8.450000 ;
        RECT  4.365000  8.680000  4.565000  8.880000 ;
        RECT  4.365000  9.110000  4.565000  9.310000 ;
        RECT  4.365000  9.540000  4.565000  9.740000 ;
        RECT  4.365000  9.970000  4.565000 10.170000 ;
        RECT  4.365000 10.400000  4.565000 10.600000 ;
        RECT  4.365000 10.830000  4.565000 11.030000 ;
        RECT  4.365000 11.260000  4.565000 11.460000 ;
        RECT  4.770000  6.960000  4.970000  7.160000 ;
        RECT  4.770000  7.390000  4.970000  7.590000 ;
        RECT  4.770000  7.820000  4.970000  8.020000 ;
        RECT  4.770000  8.250000  4.970000  8.450000 ;
        RECT  4.770000  8.680000  4.970000  8.880000 ;
        RECT  4.770000  9.110000  4.970000  9.310000 ;
        RECT  4.770000  9.540000  4.970000  9.740000 ;
        RECT  4.770000  9.970000  4.970000 10.170000 ;
        RECT  4.770000 10.400000  4.970000 10.600000 ;
        RECT  4.770000 10.830000  4.970000 11.030000 ;
        RECT  4.770000 11.260000  4.970000 11.460000 ;
        RECT  5.175000  6.960000  5.375000  7.160000 ;
        RECT  5.175000  7.390000  5.375000  7.590000 ;
        RECT  5.175000  7.820000  5.375000  8.020000 ;
        RECT  5.175000  8.250000  5.375000  8.450000 ;
        RECT  5.175000  8.680000  5.375000  8.880000 ;
        RECT  5.175000  9.110000  5.375000  9.310000 ;
        RECT  5.175000  9.540000  5.375000  9.740000 ;
        RECT  5.175000  9.970000  5.375000 10.170000 ;
        RECT  5.175000 10.400000  5.375000 10.600000 ;
        RECT  5.175000 10.830000  5.375000 11.030000 ;
        RECT  5.175000 11.260000  5.375000 11.460000 ;
        RECT  5.580000  6.960000  5.780000  7.160000 ;
        RECT  5.580000  7.390000  5.780000  7.590000 ;
        RECT  5.580000  7.820000  5.780000  8.020000 ;
        RECT  5.580000  8.250000  5.780000  8.450000 ;
        RECT  5.580000  8.680000  5.780000  8.880000 ;
        RECT  5.580000  9.110000  5.780000  9.310000 ;
        RECT  5.580000  9.540000  5.780000  9.740000 ;
        RECT  5.580000  9.970000  5.780000 10.170000 ;
        RECT  5.580000 10.400000  5.780000 10.600000 ;
        RECT  5.580000 10.830000  5.780000 11.030000 ;
        RECT  5.580000 11.260000  5.780000 11.460000 ;
        RECT  5.985000  6.960000  6.185000  7.160000 ;
        RECT  5.985000  7.390000  6.185000  7.590000 ;
        RECT  5.985000  7.820000  6.185000  8.020000 ;
        RECT  5.985000  8.250000  6.185000  8.450000 ;
        RECT  5.985000  8.680000  6.185000  8.880000 ;
        RECT  5.985000  9.110000  6.185000  9.310000 ;
        RECT  5.985000  9.540000  6.185000  9.740000 ;
        RECT  5.985000  9.970000  6.185000 10.170000 ;
        RECT  5.985000 10.400000  6.185000 10.600000 ;
        RECT  5.985000 10.830000  6.185000 11.030000 ;
        RECT  5.985000 11.260000  6.185000 11.460000 ;
        RECT  6.390000  6.960000  6.590000  7.160000 ;
        RECT  6.390000  7.390000  6.590000  7.590000 ;
        RECT  6.390000  7.820000  6.590000  8.020000 ;
        RECT  6.390000  8.250000  6.590000  8.450000 ;
        RECT  6.390000  8.680000  6.590000  8.880000 ;
        RECT  6.390000  9.110000  6.590000  9.310000 ;
        RECT  6.390000  9.540000  6.590000  9.740000 ;
        RECT  6.390000  9.970000  6.590000 10.170000 ;
        RECT  6.390000 10.400000  6.590000 10.600000 ;
        RECT  6.390000 10.830000  6.590000 11.030000 ;
        RECT  6.390000 11.260000  6.590000 11.460000 ;
        RECT  6.795000  6.960000  6.995000  7.160000 ;
        RECT  6.795000  7.390000  6.995000  7.590000 ;
        RECT  6.795000  7.820000  6.995000  8.020000 ;
        RECT  6.795000  8.250000  6.995000  8.450000 ;
        RECT  6.795000  8.680000  6.995000  8.880000 ;
        RECT  6.795000  9.110000  6.995000  9.310000 ;
        RECT  6.795000  9.540000  6.995000  9.740000 ;
        RECT  6.795000  9.970000  6.995000 10.170000 ;
        RECT  6.795000 10.400000  6.995000 10.600000 ;
        RECT  6.795000 10.830000  6.995000 11.030000 ;
        RECT  6.795000 11.260000  6.995000 11.460000 ;
        RECT  7.200000  6.960000  7.400000  7.160000 ;
        RECT  7.200000  7.390000  7.400000  7.590000 ;
        RECT  7.200000  7.820000  7.400000  8.020000 ;
        RECT  7.200000  8.250000  7.400000  8.450000 ;
        RECT  7.200000  8.680000  7.400000  8.880000 ;
        RECT  7.200000  9.110000  7.400000  9.310000 ;
        RECT  7.200000  9.540000  7.400000  9.740000 ;
        RECT  7.200000  9.970000  7.400000 10.170000 ;
        RECT  7.200000 10.400000  7.400000 10.600000 ;
        RECT  7.200000 10.830000  7.400000 11.030000 ;
        RECT  7.200000 11.260000  7.400000 11.460000 ;
        RECT  7.605000  6.960000  7.805000  7.160000 ;
        RECT  7.605000  7.390000  7.805000  7.590000 ;
        RECT  7.605000  7.820000  7.805000  8.020000 ;
        RECT  7.605000  8.250000  7.805000  8.450000 ;
        RECT  7.605000  8.680000  7.805000  8.880000 ;
        RECT  7.605000  9.110000  7.805000  9.310000 ;
        RECT  7.605000  9.540000  7.805000  9.740000 ;
        RECT  7.605000  9.970000  7.805000 10.170000 ;
        RECT  7.605000 10.400000  7.805000 10.600000 ;
        RECT  7.605000 10.830000  7.805000 11.030000 ;
        RECT  7.605000 11.260000  7.805000 11.460000 ;
        RECT  8.010000  6.960000  8.210000  7.160000 ;
        RECT  8.010000  7.390000  8.210000  7.590000 ;
        RECT  8.010000  7.820000  8.210000  8.020000 ;
        RECT  8.010000  8.250000  8.210000  8.450000 ;
        RECT  8.010000  8.680000  8.210000  8.880000 ;
        RECT  8.010000  9.110000  8.210000  9.310000 ;
        RECT  8.010000  9.540000  8.210000  9.740000 ;
        RECT  8.010000  9.970000  8.210000 10.170000 ;
        RECT  8.010000 10.400000  8.210000 10.600000 ;
        RECT  8.010000 10.830000  8.210000 11.030000 ;
        RECT  8.010000 11.260000  8.210000 11.460000 ;
        RECT  8.415000  6.960000  8.615000  7.160000 ;
        RECT  8.415000  7.390000  8.615000  7.590000 ;
        RECT  8.415000  7.820000  8.615000  8.020000 ;
        RECT  8.415000  8.250000  8.615000  8.450000 ;
        RECT  8.415000  8.680000  8.615000  8.880000 ;
        RECT  8.415000  9.110000  8.615000  9.310000 ;
        RECT  8.415000  9.540000  8.615000  9.740000 ;
        RECT  8.415000  9.970000  8.615000 10.170000 ;
        RECT  8.415000 10.400000  8.615000 10.600000 ;
        RECT  8.415000 10.830000  8.615000 11.030000 ;
        RECT  8.415000 11.260000  8.615000 11.460000 ;
        RECT  8.820000  6.960000  9.020000  7.160000 ;
        RECT  8.820000  7.390000  9.020000  7.590000 ;
        RECT  8.820000  7.820000  9.020000  8.020000 ;
        RECT  8.820000  8.250000  9.020000  8.450000 ;
        RECT  8.820000  8.680000  9.020000  8.880000 ;
        RECT  8.820000  9.110000  9.020000  9.310000 ;
        RECT  8.820000  9.540000  9.020000  9.740000 ;
        RECT  8.820000  9.970000  9.020000 10.170000 ;
        RECT  8.820000 10.400000  9.020000 10.600000 ;
        RECT  8.820000 10.830000  9.020000 11.030000 ;
        RECT  8.820000 11.260000  9.020000 11.460000 ;
        RECT  9.225000  6.960000  9.425000  7.160000 ;
        RECT  9.225000  7.390000  9.425000  7.590000 ;
        RECT  9.225000  7.820000  9.425000  8.020000 ;
        RECT  9.225000  8.250000  9.425000  8.450000 ;
        RECT  9.225000  8.680000  9.425000  8.880000 ;
        RECT  9.225000  9.110000  9.425000  9.310000 ;
        RECT  9.225000  9.540000  9.425000  9.740000 ;
        RECT  9.225000  9.970000  9.425000 10.170000 ;
        RECT  9.225000 10.400000  9.425000 10.600000 ;
        RECT  9.225000 10.830000  9.425000 11.030000 ;
        RECT  9.225000 11.260000  9.425000 11.460000 ;
        RECT  9.630000  6.960000  9.830000  7.160000 ;
        RECT  9.630000  7.390000  9.830000  7.590000 ;
        RECT  9.630000  7.820000  9.830000  8.020000 ;
        RECT  9.630000  8.250000  9.830000  8.450000 ;
        RECT  9.630000  8.680000  9.830000  8.880000 ;
        RECT  9.630000  9.110000  9.830000  9.310000 ;
        RECT  9.630000  9.540000  9.830000  9.740000 ;
        RECT  9.630000  9.970000  9.830000 10.170000 ;
        RECT  9.630000 10.400000  9.830000 10.600000 ;
        RECT  9.630000 10.830000  9.830000 11.030000 ;
        RECT  9.630000 11.260000  9.830000 11.460000 ;
        RECT 10.035000  6.960000 10.235000  7.160000 ;
        RECT 10.035000  7.390000 10.235000  7.590000 ;
        RECT 10.035000  7.820000 10.235000  8.020000 ;
        RECT 10.035000  8.250000 10.235000  8.450000 ;
        RECT 10.035000  8.680000 10.235000  8.880000 ;
        RECT 10.035000  9.110000 10.235000  9.310000 ;
        RECT 10.035000  9.540000 10.235000  9.740000 ;
        RECT 10.035000  9.970000 10.235000 10.170000 ;
        RECT 10.035000 10.400000 10.235000 10.600000 ;
        RECT 10.035000 10.830000 10.235000 11.030000 ;
        RECT 10.035000 11.260000 10.235000 11.460000 ;
        RECT 10.440000  6.960000 10.640000  7.160000 ;
        RECT 10.440000  7.390000 10.640000  7.590000 ;
        RECT 10.440000  7.820000 10.640000  8.020000 ;
        RECT 10.440000  8.250000 10.640000  8.450000 ;
        RECT 10.440000  8.680000 10.640000  8.880000 ;
        RECT 10.440000  9.110000 10.640000  9.310000 ;
        RECT 10.440000  9.540000 10.640000  9.740000 ;
        RECT 10.440000  9.970000 10.640000 10.170000 ;
        RECT 10.440000 10.400000 10.640000 10.600000 ;
        RECT 10.440000 10.830000 10.640000 11.030000 ;
        RECT 10.440000 11.260000 10.640000 11.460000 ;
        RECT 10.845000  6.960000 11.045000  7.160000 ;
        RECT 10.845000  7.390000 11.045000  7.590000 ;
        RECT 10.845000  7.820000 11.045000  8.020000 ;
        RECT 10.845000  8.250000 11.045000  8.450000 ;
        RECT 10.845000  8.680000 11.045000  8.880000 ;
        RECT 10.845000  9.110000 11.045000  9.310000 ;
        RECT 10.845000  9.540000 11.045000  9.740000 ;
        RECT 10.845000  9.970000 11.045000 10.170000 ;
        RECT 10.845000 10.400000 11.045000 10.600000 ;
        RECT 10.845000 10.830000 11.045000 11.030000 ;
        RECT 10.845000 11.260000 11.045000 11.460000 ;
        RECT 11.250000  6.960000 11.450000  7.160000 ;
        RECT 11.250000  7.390000 11.450000  7.590000 ;
        RECT 11.250000  7.820000 11.450000  8.020000 ;
        RECT 11.250000  8.250000 11.450000  8.450000 ;
        RECT 11.250000  8.680000 11.450000  8.880000 ;
        RECT 11.250000  9.110000 11.450000  9.310000 ;
        RECT 11.250000  9.540000 11.450000  9.740000 ;
        RECT 11.250000  9.970000 11.450000 10.170000 ;
        RECT 11.250000 10.400000 11.450000 10.600000 ;
        RECT 11.250000 10.830000 11.450000 11.030000 ;
        RECT 11.250000 11.260000 11.450000 11.460000 ;
        RECT 11.655000  6.960000 11.855000  7.160000 ;
        RECT 11.655000  7.390000 11.855000  7.590000 ;
        RECT 11.655000  7.820000 11.855000  8.020000 ;
        RECT 11.655000  8.250000 11.855000  8.450000 ;
        RECT 11.655000  8.680000 11.855000  8.880000 ;
        RECT 11.655000  9.110000 11.855000  9.310000 ;
        RECT 11.655000  9.540000 11.855000  9.740000 ;
        RECT 11.655000  9.970000 11.855000 10.170000 ;
        RECT 11.655000 10.400000 11.855000 10.600000 ;
        RECT 11.655000 10.830000 11.855000 11.030000 ;
        RECT 11.655000 11.260000 11.855000 11.460000 ;
        RECT 12.060000  6.960000 12.260000  7.160000 ;
        RECT 12.060000  7.390000 12.260000  7.590000 ;
        RECT 12.060000  7.820000 12.260000  8.020000 ;
        RECT 12.060000  8.250000 12.260000  8.450000 ;
        RECT 12.060000  8.680000 12.260000  8.880000 ;
        RECT 12.060000  9.110000 12.260000  9.310000 ;
        RECT 12.060000  9.540000 12.260000  9.740000 ;
        RECT 12.060000  9.970000 12.260000 10.170000 ;
        RECT 12.060000 10.400000 12.260000 10.600000 ;
        RECT 12.060000 10.830000 12.260000 11.030000 ;
        RECT 12.060000 11.260000 12.260000 11.460000 ;
        RECT 12.465000  6.960000 12.665000  7.160000 ;
        RECT 12.465000  7.390000 12.665000  7.590000 ;
        RECT 12.465000  7.820000 12.665000  8.020000 ;
        RECT 12.465000  8.250000 12.665000  8.450000 ;
        RECT 12.465000  8.680000 12.665000  8.880000 ;
        RECT 12.465000  9.110000 12.665000  9.310000 ;
        RECT 12.465000  9.540000 12.665000  9.740000 ;
        RECT 12.465000  9.970000 12.665000 10.170000 ;
        RECT 12.465000 10.400000 12.665000 10.600000 ;
        RECT 12.465000 10.830000 12.665000 11.030000 ;
        RECT 12.465000 11.260000 12.665000 11.460000 ;
        RECT 12.870000  6.960000 13.070000  7.160000 ;
        RECT 12.870000  7.390000 13.070000  7.590000 ;
        RECT 12.870000  7.820000 13.070000  8.020000 ;
        RECT 12.870000  8.250000 13.070000  8.450000 ;
        RECT 12.870000  8.680000 13.070000  8.880000 ;
        RECT 12.870000  9.110000 13.070000  9.310000 ;
        RECT 12.870000  9.540000 13.070000  9.740000 ;
        RECT 12.870000  9.970000 13.070000 10.170000 ;
        RECT 12.870000 10.400000 13.070000 10.600000 ;
        RECT 12.870000 10.830000 13.070000 11.030000 ;
        RECT 12.870000 11.260000 13.070000 11.460000 ;
        RECT 13.275000  6.960000 13.475000  7.160000 ;
        RECT 13.275000  7.390000 13.475000  7.590000 ;
        RECT 13.275000  7.820000 13.475000  8.020000 ;
        RECT 13.275000  8.250000 13.475000  8.450000 ;
        RECT 13.275000  8.680000 13.475000  8.880000 ;
        RECT 13.275000  9.110000 13.475000  9.310000 ;
        RECT 13.275000  9.540000 13.475000  9.740000 ;
        RECT 13.275000  9.970000 13.475000 10.170000 ;
        RECT 13.275000 10.400000 13.475000 10.600000 ;
        RECT 13.275000 10.830000 13.475000 11.030000 ;
        RECT 13.275000 11.260000 13.475000 11.460000 ;
        RECT 13.680000  6.960000 13.880000  7.160000 ;
        RECT 13.680000  7.390000 13.880000  7.590000 ;
        RECT 13.680000  7.820000 13.880000  8.020000 ;
        RECT 13.680000  8.250000 13.880000  8.450000 ;
        RECT 13.680000  8.680000 13.880000  8.880000 ;
        RECT 13.680000  9.110000 13.880000  9.310000 ;
        RECT 13.680000  9.540000 13.880000  9.740000 ;
        RECT 13.680000  9.970000 13.880000 10.170000 ;
        RECT 13.680000 10.400000 13.880000 10.600000 ;
        RECT 13.680000 10.830000 13.880000 11.030000 ;
        RECT 13.680000 11.260000 13.880000 11.460000 ;
        RECT 14.085000  6.960000 14.285000  7.160000 ;
        RECT 14.085000  7.390000 14.285000  7.590000 ;
        RECT 14.085000  7.820000 14.285000  8.020000 ;
        RECT 14.085000  8.250000 14.285000  8.450000 ;
        RECT 14.085000  8.680000 14.285000  8.880000 ;
        RECT 14.085000  9.110000 14.285000  9.310000 ;
        RECT 14.085000  9.540000 14.285000  9.740000 ;
        RECT 14.085000  9.970000 14.285000 10.170000 ;
        RECT 14.085000 10.400000 14.285000 10.600000 ;
        RECT 14.085000 10.830000 14.285000 11.030000 ;
        RECT 14.085000 11.260000 14.285000 11.460000 ;
        RECT 14.490000  6.960000 14.690000  7.160000 ;
        RECT 14.490000  7.390000 14.690000  7.590000 ;
        RECT 14.490000  7.820000 14.690000  8.020000 ;
        RECT 14.490000  8.250000 14.690000  8.450000 ;
        RECT 14.490000  8.680000 14.690000  8.880000 ;
        RECT 14.490000  9.110000 14.690000  9.310000 ;
        RECT 14.490000  9.540000 14.690000  9.740000 ;
        RECT 14.490000  9.970000 14.690000 10.170000 ;
        RECT 14.490000 10.400000 14.690000 10.600000 ;
        RECT 14.490000 10.830000 14.690000 11.030000 ;
        RECT 14.490000 11.260000 14.690000 11.460000 ;
        RECT 14.895000  6.960000 15.095000  7.160000 ;
        RECT 14.895000  7.390000 15.095000  7.590000 ;
        RECT 14.895000  7.820000 15.095000  8.020000 ;
        RECT 14.895000  8.250000 15.095000  8.450000 ;
        RECT 14.895000  8.680000 15.095000  8.880000 ;
        RECT 14.895000  9.110000 15.095000  9.310000 ;
        RECT 14.895000  9.540000 15.095000  9.740000 ;
        RECT 14.895000  9.970000 15.095000 10.170000 ;
        RECT 14.895000 10.400000 15.095000 10.600000 ;
        RECT 14.895000 10.830000 15.095000 11.030000 ;
        RECT 14.895000 11.260000 15.095000 11.460000 ;
        RECT 15.300000  6.960000 15.500000  7.160000 ;
        RECT 15.300000  7.390000 15.500000  7.590000 ;
        RECT 15.300000  7.820000 15.500000  8.020000 ;
        RECT 15.300000  8.250000 15.500000  8.450000 ;
        RECT 15.300000  8.680000 15.500000  8.880000 ;
        RECT 15.300000  9.110000 15.500000  9.310000 ;
        RECT 15.300000  9.540000 15.500000  9.740000 ;
        RECT 15.300000  9.970000 15.500000 10.170000 ;
        RECT 15.300000 10.400000 15.500000 10.600000 ;
        RECT 15.300000 10.830000 15.500000 11.030000 ;
        RECT 15.300000 11.260000 15.500000 11.460000 ;
        RECT 15.705000  6.960000 15.905000  7.160000 ;
        RECT 15.705000  7.390000 15.905000  7.590000 ;
        RECT 15.705000  7.820000 15.905000  8.020000 ;
        RECT 15.705000  8.250000 15.905000  8.450000 ;
        RECT 15.705000  8.680000 15.905000  8.880000 ;
        RECT 15.705000  9.110000 15.905000  9.310000 ;
        RECT 15.705000  9.540000 15.905000  9.740000 ;
        RECT 15.705000  9.970000 15.905000 10.170000 ;
        RECT 15.705000 10.400000 15.905000 10.600000 ;
        RECT 15.705000 10.830000 15.905000 11.030000 ;
        RECT 15.705000 11.260000 15.905000 11.460000 ;
        RECT 16.110000  6.960000 16.310000  7.160000 ;
        RECT 16.110000  7.390000 16.310000  7.590000 ;
        RECT 16.110000  7.820000 16.310000  8.020000 ;
        RECT 16.110000  8.250000 16.310000  8.450000 ;
        RECT 16.110000  8.680000 16.310000  8.880000 ;
        RECT 16.110000  9.110000 16.310000  9.310000 ;
        RECT 16.110000  9.540000 16.310000  9.740000 ;
        RECT 16.110000  9.970000 16.310000 10.170000 ;
        RECT 16.110000 10.400000 16.310000 10.600000 ;
        RECT 16.110000 10.830000 16.310000 11.030000 ;
        RECT 16.110000 11.260000 16.310000 11.460000 ;
        RECT 16.515000  6.960000 16.715000  7.160000 ;
        RECT 16.515000  7.390000 16.715000  7.590000 ;
        RECT 16.515000  7.820000 16.715000  8.020000 ;
        RECT 16.515000  8.250000 16.715000  8.450000 ;
        RECT 16.515000  8.680000 16.715000  8.880000 ;
        RECT 16.515000  9.110000 16.715000  9.310000 ;
        RECT 16.515000  9.540000 16.715000  9.740000 ;
        RECT 16.515000  9.970000 16.715000 10.170000 ;
        RECT 16.515000 10.400000 16.715000 10.600000 ;
        RECT 16.515000 10.830000 16.715000 11.030000 ;
        RECT 16.515000 11.260000 16.715000 11.460000 ;
        RECT 16.920000  6.960000 17.120000  7.160000 ;
        RECT 16.920000  7.390000 17.120000  7.590000 ;
        RECT 16.920000  7.820000 17.120000  8.020000 ;
        RECT 16.920000  8.250000 17.120000  8.450000 ;
        RECT 16.920000  8.680000 17.120000  8.880000 ;
        RECT 16.920000  9.110000 17.120000  9.310000 ;
        RECT 16.920000  9.540000 17.120000  9.740000 ;
        RECT 16.920000  9.970000 17.120000 10.170000 ;
        RECT 16.920000 10.400000 17.120000 10.600000 ;
        RECT 16.920000 10.830000 17.120000 11.030000 ;
        RECT 16.920000 11.260000 17.120000 11.460000 ;
        RECT 17.325000  6.960000 17.525000  7.160000 ;
        RECT 17.325000  7.390000 17.525000  7.590000 ;
        RECT 17.325000  7.820000 17.525000  8.020000 ;
        RECT 17.325000  8.250000 17.525000  8.450000 ;
        RECT 17.325000  8.680000 17.525000  8.880000 ;
        RECT 17.325000  9.110000 17.525000  9.310000 ;
        RECT 17.325000  9.540000 17.525000  9.740000 ;
        RECT 17.325000  9.970000 17.525000 10.170000 ;
        RECT 17.325000 10.400000 17.525000 10.600000 ;
        RECT 17.325000 10.830000 17.525000 11.030000 ;
        RECT 17.325000 11.260000 17.525000 11.460000 ;
        RECT 17.730000  6.960000 17.930000  7.160000 ;
        RECT 17.730000  7.390000 17.930000  7.590000 ;
        RECT 17.730000  7.820000 17.930000  8.020000 ;
        RECT 17.730000  8.250000 17.930000  8.450000 ;
        RECT 17.730000  8.680000 17.930000  8.880000 ;
        RECT 17.730000  9.110000 17.930000  9.310000 ;
        RECT 17.730000  9.540000 17.930000  9.740000 ;
        RECT 17.730000  9.970000 17.930000 10.170000 ;
        RECT 17.730000 10.400000 17.930000 10.600000 ;
        RECT 17.730000 10.830000 17.930000 11.030000 ;
        RECT 17.730000 11.260000 17.930000 11.460000 ;
        RECT 18.135000  6.960000 18.335000  7.160000 ;
        RECT 18.135000  7.390000 18.335000  7.590000 ;
        RECT 18.135000  7.820000 18.335000  8.020000 ;
        RECT 18.135000  8.250000 18.335000  8.450000 ;
        RECT 18.135000  8.680000 18.335000  8.880000 ;
        RECT 18.135000  9.110000 18.335000  9.310000 ;
        RECT 18.135000  9.540000 18.335000  9.740000 ;
        RECT 18.135000  9.970000 18.335000 10.170000 ;
        RECT 18.135000 10.400000 18.335000 10.600000 ;
        RECT 18.135000 10.830000 18.335000 11.030000 ;
        RECT 18.135000 11.260000 18.335000 11.460000 ;
        RECT 18.540000  6.960000 18.740000  7.160000 ;
        RECT 18.540000  7.390000 18.740000  7.590000 ;
        RECT 18.540000  7.820000 18.740000  8.020000 ;
        RECT 18.540000  8.250000 18.740000  8.450000 ;
        RECT 18.540000  8.680000 18.740000  8.880000 ;
        RECT 18.540000  9.110000 18.740000  9.310000 ;
        RECT 18.540000  9.540000 18.740000  9.740000 ;
        RECT 18.540000  9.970000 18.740000 10.170000 ;
        RECT 18.540000 10.400000 18.740000 10.600000 ;
        RECT 18.540000 10.830000 18.740000 11.030000 ;
        RECT 18.540000 11.260000 18.740000 11.460000 ;
        RECT 18.945000  6.960000 19.145000  7.160000 ;
        RECT 18.945000  7.390000 19.145000  7.590000 ;
        RECT 18.945000  7.820000 19.145000  8.020000 ;
        RECT 18.945000  8.250000 19.145000  8.450000 ;
        RECT 18.945000  8.680000 19.145000  8.880000 ;
        RECT 18.945000  9.110000 19.145000  9.310000 ;
        RECT 18.945000  9.540000 19.145000  9.740000 ;
        RECT 18.945000  9.970000 19.145000 10.170000 ;
        RECT 18.945000 10.400000 19.145000 10.600000 ;
        RECT 18.945000 10.830000 19.145000 11.030000 ;
        RECT 18.945000 11.260000 19.145000 11.460000 ;
        RECT 19.350000  6.960000 19.550000  7.160000 ;
        RECT 19.350000  7.390000 19.550000  7.590000 ;
        RECT 19.350000  7.820000 19.550000  8.020000 ;
        RECT 19.350000  8.250000 19.550000  8.450000 ;
        RECT 19.350000  8.680000 19.550000  8.880000 ;
        RECT 19.350000  9.110000 19.550000  9.310000 ;
        RECT 19.350000  9.540000 19.550000  9.740000 ;
        RECT 19.350000  9.970000 19.550000 10.170000 ;
        RECT 19.350000 10.400000 19.550000 10.600000 ;
        RECT 19.350000 10.830000 19.550000 11.030000 ;
        RECT 19.350000 11.260000 19.550000 11.460000 ;
        RECT 19.755000  6.960000 19.955000  7.160000 ;
        RECT 19.755000  7.390000 19.955000  7.590000 ;
        RECT 19.755000  7.820000 19.955000  8.020000 ;
        RECT 19.755000  8.250000 19.955000  8.450000 ;
        RECT 19.755000  8.680000 19.955000  8.880000 ;
        RECT 19.755000  9.110000 19.955000  9.310000 ;
        RECT 19.755000  9.540000 19.955000  9.740000 ;
        RECT 19.755000  9.970000 19.955000 10.170000 ;
        RECT 19.755000 10.400000 19.955000 10.600000 ;
        RECT 19.755000 10.830000 19.955000 11.030000 ;
        RECT 19.755000 11.260000 19.955000 11.460000 ;
        RECT 20.160000  6.960000 20.360000  7.160000 ;
        RECT 20.160000  7.390000 20.360000  7.590000 ;
        RECT 20.160000  7.820000 20.360000  8.020000 ;
        RECT 20.160000  8.250000 20.360000  8.450000 ;
        RECT 20.160000  8.680000 20.360000  8.880000 ;
        RECT 20.160000  9.110000 20.360000  9.310000 ;
        RECT 20.160000  9.540000 20.360000  9.740000 ;
        RECT 20.160000  9.970000 20.360000 10.170000 ;
        RECT 20.160000 10.400000 20.360000 10.600000 ;
        RECT 20.160000 10.830000 20.360000 11.030000 ;
        RECT 20.160000 11.260000 20.360000 11.460000 ;
        RECT 20.565000  6.960000 20.765000  7.160000 ;
        RECT 20.565000  7.390000 20.765000  7.590000 ;
        RECT 20.565000  7.820000 20.765000  8.020000 ;
        RECT 20.565000  8.250000 20.765000  8.450000 ;
        RECT 20.565000  8.680000 20.765000  8.880000 ;
        RECT 20.565000  9.110000 20.765000  9.310000 ;
        RECT 20.565000  9.540000 20.765000  9.740000 ;
        RECT 20.565000  9.970000 20.765000 10.170000 ;
        RECT 20.565000 10.400000 20.765000 10.600000 ;
        RECT 20.565000 10.830000 20.765000 11.030000 ;
        RECT 20.565000 11.260000 20.765000 11.460000 ;
        RECT 20.970000  6.960000 21.170000  7.160000 ;
        RECT 20.970000  7.390000 21.170000  7.590000 ;
        RECT 20.970000  7.820000 21.170000  8.020000 ;
        RECT 20.970000  8.250000 21.170000  8.450000 ;
        RECT 20.970000  8.680000 21.170000  8.880000 ;
        RECT 20.970000  9.110000 21.170000  9.310000 ;
        RECT 20.970000  9.540000 21.170000  9.740000 ;
        RECT 20.970000  9.970000 21.170000 10.170000 ;
        RECT 20.970000 10.400000 21.170000 10.600000 ;
        RECT 20.970000 10.830000 21.170000 11.030000 ;
        RECT 20.970000 11.260000 21.170000 11.460000 ;
        RECT 21.375000  6.960000 21.575000  7.160000 ;
        RECT 21.375000  7.390000 21.575000  7.590000 ;
        RECT 21.375000  7.820000 21.575000  8.020000 ;
        RECT 21.375000  8.250000 21.575000  8.450000 ;
        RECT 21.375000  8.680000 21.575000  8.880000 ;
        RECT 21.375000  9.110000 21.575000  9.310000 ;
        RECT 21.375000  9.540000 21.575000  9.740000 ;
        RECT 21.375000  9.970000 21.575000 10.170000 ;
        RECT 21.375000 10.400000 21.575000 10.600000 ;
        RECT 21.375000 10.830000 21.575000 11.030000 ;
        RECT 21.375000 11.260000 21.575000 11.460000 ;
        RECT 21.780000  6.960000 21.980000  7.160000 ;
        RECT 21.780000  7.390000 21.980000  7.590000 ;
        RECT 21.780000  7.820000 21.980000  8.020000 ;
        RECT 21.780000  8.250000 21.980000  8.450000 ;
        RECT 21.780000  8.680000 21.980000  8.880000 ;
        RECT 21.780000  9.110000 21.980000  9.310000 ;
        RECT 21.780000  9.540000 21.980000  9.740000 ;
        RECT 21.780000  9.970000 21.980000 10.170000 ;
        RECT 21.780000 10.400000 21.980000 10.600000 ;
        RECT 21.780000 10.830000 21.980000 11.030000 ;
        RECT 21.780000 11.260000 21.980000 11.460000 ;
        RECT 22.185000  6.960000 22.385000  7.160000 ;
        RECT 22.185000  7.390000 22.385000  7.590000 ;
        RECT 22.185000  7.820000 22.385000  8.020000 ;
        RECT 22.185000  8.250000 22.385000  8.450000 ;
        RECT 22.185000  8.680000 22.385000  8.880000 ;
        RECT 22.185000  9.110000 22.385000  9.310000 ;
        RECT 22.185000  9.540000 22.385000  9.740000 ;
        RECT 22.185000  9.970000 22.385000 10.170000 ;
        RECT 22.185000 10.400000 22.385000 10.600000 ;
        RECT 22.185000 10.830000 22.385000 11.030000 ;
        RECT 22.185000 11.260000 22.385000 11.460000 ;
        RECT 22.590000  6.960000 22.790000  7.160000 ;
        RECT 22.590000  7.390000 22.790000  7.590000 ;
        RECT 22.590000  7.820000 22.790000  8.020000 ;
        RECT 22.590000  8.250000 22.790000  8.450000 ;
        RECT 22.590000  8.680000 22.790000  8.880000 ;
        RECT 22.590000  9.110000 22.790000  9.310000 ;
        RECT 22.590000  9.540000 22.790000  9.740000 ;
        RECT 22.590000  9.970000 22.790000 10.170000 ;
        RECT 22.590000 10.400000 22.790000 10.600000 ;
        RECT 22.590000 10.830000 22.790000 11.030000 ;
        RECT 22.590000 11.260000 22.790000 11.460000 ;
        RECT 22.995000  6.960000 23.195000  7.160000 ;
        RECT 22.995000  7.390000 23.195000  7.590000 ;
        RECT 22.995000  7.820000 23.195000  8.020000 ;
        RECT 22.995000  8.250000 23.195000  8.450000 ;
        RECT 22.995000  8.680000 23.195000  8.880000 ;
        RECT 22.995000  9.110000 23.195000  9.310000 ;
        RECT 22.995000  9.540000 23.195000  9.740000 ;
        RECT 22.995000  9.970000 23.195000 10.170000 ;
        RECT 22.995000 10.400000 23.195000 10.600000 ;
        RECT 22.995000 10.830000 23.195000 11.030000 ;
        RECT 22.995000 11.260000 23.195000 11.460000 ;
        RECT 23.400000  6.960000 23.600000  7.160000 ;
        RECT 23.400000  7.390000 23.600000  7.590000 ;
        RECT 23.400000  7.820000 23.600000  8.020000 ;
        RECT 23.400000  8.250000 23.600000  8.450000 ;
        RECT 23.400000  8.680000 23.600000  8.880000 ;
        RECT 23.400000  9.110000 23.600000  9.310000 ;
        RECT 23.400000  9.540000 23.600000  9.740000 ;
        RECT 23.400000  9.970000 23.600000 10.170000 ;
        RECT 23.400000 10.400000 23.600000 10.600000 ;
        RECT 23.400000 10.830000 23.600000 11.030000 ;
        RECT 23.400000 11.260000 23.600000 11.460000 ;
        RECT 23.805000  6.960000 24.005000  7.160000 ;
        RECT 23.805000  7.390000 24.005000  7.590000 ;
        RECT 23.805000  7.820000 24.005000  8.020000 ;
        RECT 23.805000  8.250000 24.005000  8.450000 ;
        RECT 23.805000  8.680000 24.005000  8.880000 ;
        RECT 23.805000  9.110000 24.005000  9.310000 ;
        RECT 23.805000  9.540000 24.005000  9.740000 ;
        RECT 23.805000  9.970000 24.005000 10.170000 ;
        RECT 23.805000 10.400000 24.005000 10.600000 ;
        RECT 23.805000 10.830000 24.005000 11.030000 ;
        RECT 23.805000 11.260000 24.005000 11.460000 ;
        RECT 24.210000  6.960000 24.410000  7.160000 ;
        RECT 24.210000  7.390000 24.410000  7.590000 ;
        RECT 24.210000  7.820000 24.410000  8.020000 ;
        RECT 24.210000  8.250000 24.410000  8.450000 ;
        RECT 24.210000  8.680000 24.410000  8.880000 ;
        RECT 24.210000  9.110000 24.410000  9.310000 ;
        RECT 24.210000  9.540000 24.410000  9.740000 ;
        RECT 24.210000  9.970000 24.410000 10.170000 ;
        RECT 24.210000 10.400000 24.410000 10.600000 ;
        RECT 24.210000 10.830000 24.410000 11.030000 ;
        RECT 24.210000 11.260000 24.410000 11.460000 ;
        RECT 50.845000  6.960000 51.045000  7.160000 ;
        RECT 50.845000  7.390000 51.045000  7.590000 ;
        RECT 50.845000  7.820000 51.045000  8.020000 ;
        RECT 50.845000  8.250000 51.045000  8.450000 ;
        RECT 50.845000  8.680000 51.045000  8.880000 ;
        RECT 50.845000  9.110000 51.045000  9.310000 ;
        RECT 50.845000  9.540000 51.045000  9.740000 ;
        RECT 50.845000  9.970000 51.045000 10.170000 ;
        RECT 50.845000 10.400000 51.045000 10.600000 ;
        RECT 50.845000 10.830000 51.045000 11.030000 ;
        RECT 50.845000 11.260000 51.045000 11.460000 ;
        RECT 51.255000  6.960000 51.455000  7.160000 ;
        RECT 51.255000  7.390000 51.455000  7.590000 ;
        RECT 51.255000  7.820000 51.455000  8.020000 ;
        RECT 51.255000  8.250000 51.455000  8.450000 ;
        RECT 51.255000  8.680000 51.455000  8.880000 ;
        RECT 51.255000  9.110000 51.455000  9.310000 ;
        RECT 51.255000  9.540000 51.455000  9.740000 ;
        RECT 51.255000  9.970000 51.455000 10.170000 ;
        RECT 51.255000 10.400000 51.455000 10.600000 ;
        RECT 51.255000 10.830000 51.455000 11.030000 ;
        RECT 51.255000 11.260000 51.455000 11.460000 ;
        RECT 51.665000  6.960000 51.865000  7.160000 ;
        RECT 51.665000  7.390000 51.865000  7.590000 ;
        RECT 51.665000  7.820000 51.865000  8.020000 ;
        RECT 51.665000  8.250000 51.865000  8.450000 ;
        RECT 51.665000  8.680000 51.865000  8.880000 ;
        RECT 51.665000  9.110000 51.865000  9.310000 ;
        RECT 51.665000  9.540000 51.865000  9.740000 ;
        RECT 51.665000  9.970000 51.865000 10.170000 ;
        RECT 51.665000 10.400000 51.865000 10.600000 ;
        RECT 51.665000 10.830000 51.865000 11.030000 ;
        RECT 51.665000 11.260000 51.865000 11.460000 ;
        RECT 52.075000  6.960000 52.275000  7.160000 ;
        RECT 52.075000  7.390000 52.275000  7.590000 ;
        RECT 52.075000  7.820000 52.275000  8.020000 ;
        RECT 52.075000  8.250000 52.275000  8.450000 ;
        RECT 52.075000  8.680000 52.275000  8.880000 ;
        RECT 52.075000  9.110000 52.275000  9.310000 ;
        RECT 52.075000  9.540000 52.275000  9.740000 ;
        RECT 52.075000  9.970000 52.275000 10.170000 ;
        RECT 52.075000 10.400000 52.275000 10.600000 ;
        RECT 52.075000 10.830000 52.275000 11.030000 ;
        RECT 52.075000 11.260000 52.275000 11.460000 ;
        RECT 52.485000  6.960000 52.685000  7.160000 ;
        RECT 52.485000  7.390000 52.685000  7.590000 ;
        RECT 52.485000  7.820000 52.685000  8.020000 ;
        RECT 52.485000  8.250000 52.685000  8.450000 ;
        RECT 52.485000  8.680000 52.685000  8.880000 ;
        RECT 52.485000  9.110000 52.685000  9.310000 ;
        RECT 52.485000  9.540000 52.685000  9.740000 ;
        RECT 52.485000  9.970000 52.685000 10.170000 ;
        RECT 52.485000 10.400000 52.685000 10.600000 ;
        RECT 52.485000 10.830000 52.685000 11.030000 ;
        RECT 52.485000 11.260000 52.685000 11.460000 ;
        RECT 52.895000  6.960000 53.095000  7.160000 ;
        RECT 52.895000  7.390000 53.095000  7.590000 ;
        RECT 52.895000  7.820000 53.095000  8.020000 ;
        RECT 52.895000  8.250000 53.095000  8.450000 ;
        RECT 52.895000  8.680000 53.095000  8.880000 ;
        RECT 52.895000  9.110000 53.095000  9.310000 ;
        RECT 52.895000  9.540000 53.095000  9.740000 ;
        RECT 52.895000  9.970000 53.095000 10.170000 ;
        RECT 52.895000 10.400000 53.095000 10.600000 ;
        RECT 52.895000 10.830000 53.095000 11.030000 ;
        RECT 52.895000 11.260000 53.095000 11.460000 ;
        RECT 53.305000  6.960000 53.505000  7.160000 ;
        RECT 53.305000  7.390000 53.505000  7.590000 ;
        RECT 53.305000  7.820000 53.505000  8.020000 ;
        RECT 53.305000  8.250000 53.505000  8.450000 ;
        RECT 53.305000  8.680000 53.505000  8.880000 ;
        RECT 53.305000  9.110000 53.505000  9.310000 ;
        RECT 53.305000  9.540000 53.505000  9.740000 ;
        RECT 53.305000  9.970000 53.505000 10.170000 ;
        RECT 53.305000 10.400000 53.505000 10.600000 ;
        RECT 53.305000 10.830000 53.505000 11.030000 ;
        RECT 53.305000 11.260000 53.505000 11.460000 ;
        RECT 53.710000  6.960000 53.910000  7.160000 ;
        RECT 53.710000  7.390000 53.910000  7.590000 ;
        RECT 53.710000  7.820000 53.910000  8.020000 ;
        RECT 53.710000  8.250000 53.910000  8.450000 ;
        RECT 53.710000  8.680000 53.910000  8.880000 ;
        RECT 53.710000  9.110000 53.910000  9.310000 ;
        RECT 53.710000  9.540000 53.910000  9.740000 ;
        RECT 53.710000  9.970000 53.910000 10.170000 ;
        RECT 53.710000 10.400000 53.910000 10.600000 ;
        RECT 53.710000 10.830000 53.910000 11.030000 ;
        RECT 53.710000 11.260000 53.910000 11.460000 ;
        RECT 54.115000  6.960000 54.315000  7.160000 ;
        RECT 54.115000  7.390000 54.315000  7.590000 ;
        RECT 54.115000  7.820000 54.315000  8.020000 ;
        RECT 54.115000  8.250000 54.315000  8.450000 ;
        RECT 54.115000  8.680000 54.315000  8.880000 ;
        RECT 54.115000  9.110000 54.315000  9.310000 ;
        RECT 54.115000  9.540000 54.315000  9.740000 ;
        RECT 54.115000  9.970000 54.315000 10.170000 ;
        RECT 54.115000 10.400000 54.315000 10.600000 ;
        RECT 54.115000 10.830000 54.315000 11.030000 ;
        RECT 54.115000 11.260000 54.315000 11.460000 ;
        RECT 54.520000  6.960000 54.720000  7.160000 ;
        RECT 54.520000  7.390000 54.720000  7.590000 ;
        RECT 54.520000  7.820000 54.720000  8.020000 ;
        RECT 54.520000  8.250000 54.720000  8.450000 ;
        RECT 54.520000  8.680000 54.720000  8.880000 ;
        RECT 54.520000  9.110000 54.720000  9.310000 ;
        RECT 54.520000  9.540000 54.720000  9.740000 ;
        RECT 54.520000  9.970000 54.720000 10.170000 ;
        RECT 54.520000 10.400000 54.720000 10.600000 ;
        RECT 54.520000 10.830000 54.720000 11.030000 ;
        RECT 54.520000 11.260000 54.720000 11.460000 ;
        RECT 54.925000  6.960000 55.125000  7.160000 ;
        RECT 54.925000  7.390000 55.125000  7.590000 ;
        RECT 54.925000  7.820000 55.125000  8.020000 ;
        RECT 54.925000  8.250000 55.125000  8.450000 ;
        RECT 54.925000  8.680000 55.125000  8.880000 ;
        RECT 54.925000  9.110000 55.125000  9.310000 ;
        RECT 54.925000  9.540000 55.125000  9.740000 ;
        RECT 54.925000  9.970000 55.125000 10.170000 ;
        RECT 54.925000 10.400000 55.125000 10.600000 ;
        RECT 54.925000 10.830000 55.125000 11.030000 ;
        RECT 54.925000 11.260000 55.125000 11.460000 ;
        RECT 55.330000  6.960000 55.530000  7.160000 ;
        RECT 55.330000  7.390000 55.530000  7.590000 ;
        RECT 55.330000  7.820000 55.530000  8.020000 ;
        RECT 55.330000  8.250000 55.530000  8.450000 ;
        RECT 55.330000  8.680000 55.530000  8.880000 ;
        RECT 55.330000  9.110000 55.530000  9.310000 ;
        RECT 55.330000  9.540000 55.530000  9.740000 ;
        RECT 55.330000  9.970000 55.530000 10.170000 ;
        RECT 55.330000 10.400000 55.530000 10.600000 ;
        RECT 55.330000 10.830000 55.530000 11.030000 ;
        RECT 55.330000 11.260000 55.530000 11.460000 ;
        RECT 55.735000  6.960000 55.935000  7.160000 ;
        RECT 55.735000  7.390000 55.935000  7.590000 ;
        RECT 55.735000  7.820000 55.935000  8.020000 ;
        RECT 55.735000  8.250000 55.935000  8.450000 ;
        RECT 55.735000  8.680000 55.935000  8.880000 ;
        RECT 55.735000  9.110000 55.935000  9.310000 ;
        RECT 55.735000  9.540000 55.935000  9.740000 ;
        RECT 55.735000  9.970000 55.935000 10.170000 ;
        RECT 55.735000 10.400000 55.935000 10.600000 ;
        RECT 55.735000 10.830000 55.935000 11.030000 ;
        RECT 55.735000 11.260000 55.935000 11.460000 ;
        RECT 56.140000  6.960000 56.340000  7.160000 ;
        RECT 56.140000  7.390000 56.340000  7.590000 ;
        RECT 56.140000  7.820000 56.340000  8.020000 ;
        RECT 56.140000  8.250000 56.340000  8.450000 ;
        RECT 56.140000  8.680000 56.340000  8.880000 ;
        RECT 56.140000  9.110000 56.340000  9.310000 ;
        RECT 56.140000  9.540000 56.340000  9.740000 ;
        RECT 56.140000  9.970000 56.340000 10.170000 ;
        RECT 56.140000 10.400000 56.340000 10.600000 ;
        RECT 56.140000 10.830000 56.340000 11.030000 ;
        RECT 56.140000 11.260000 56.340000 11.460000 ;
        RECT 56.545000  6.960000 56.745000  7.160000 ;
        RECT 56.545000  7.390000 56.745000  7.590000 ;
        RECT 56.545000  7.820000 56.745000  8.020000 ;
        RECT 56.545000  8.250000 56.745000  8.450000 ;
        RECT 56.545000  8.680000 56.745000  8.880000 ;
        RECT 56.545000  9.110000 56.745000  9.310000 ;
        RECT 56.545000  9.540000 56.745000  9.740000 ;
        RECT 56.545000  9.970000 56.745000 10.170000 ;
        RECT 56.545000 10.400000 56.745000 10.600000 ;
        RECT 56.545000 10.830000 56.745000 11.030000 ;
        RECT 56.545000 11.260000 56.745000 11.460000 ;
        RECT 56.950000  6.960000 57.150000  7.160000 ;
        RECT 56.950000  7.390000 57.150000  7.590000 ;
        RECT 56.950000  7.820000 57.150000  8.020000 ;
        RECT 56.950000  8.250000 57.150000  8.450000 ;
        RECT 56.950000  8.680000 57.150000  8.880000 ;
        RECT 56.950000  9.110000 57.150000  9.310000 ;
        RECT 56.950000  9.540000 57.150000  9.740000 ;
        RECT 56.950000  9.970000 57.150000 10.170000 ;
        RECT 56.950000 10.400000 57.150000 10.600000 ;
        RECT 56.950000 10.830000 57.150000 11.030000 ;
        RECT 56.950000 11.260000 57.150000 11.460000 ;
        RECT 57.355000  6.960000 57.555000  7.160000 ;
        RECT 57.355000  7.390000 57.555000  7.590000 ;
        RECT 57.355000  7.820000 57.555000  8.020000 ;
        RECT 57.355000  8.250000 57.555000  8.450000 ;
        RECT 57.355000  8.680000 57.555000  8.880000 ;
        RECT 57.355000  9.110000 57.555000  9.310000 ;
        RECT 57.355000  9.540000 57.555000  9.740000 ;
        RECT 57.355000  9.970000 57.555000 10.170000 ;
        RECT 57.355000 10.400000 57.555000 10.600000 ;
        RECT 57.355000 10.830000 57.555000 11.030000 ;
        RECT 57.355000 11.260000 57.555000 11.460000 ;
        RECT 57.760000  6.960000 57.960000  7.160000 ;
        RECT 57.760000  7.390000 57.960000  7.590000 ;
        RECT 57.760000  7.820000 57.960000  8.020000 ;
        RECT 57.760000  8.250000 57.960000  8.450000 ;
        RECT 57.760000  8.680000 57.960000  8.880000 ;
        RECT 57.760000  9.110000 57.960000  9.310000 ;
        RECT 57.760000  9.540000 57.960000  9.740000 ;
        RECT 57.760000  9.970000 57.960000 10.170000 ;
        RECT 57.760000 10.400000 57.960000 10.600000 ;
        RECT 57.760000 10.830000 57.960000 11.030000 ;
        RECT 57.760000 11.260000 57.960000 11.460000 ;
        RECT 58.165000  6.960000 58.365000  7.160000 ;
        RECT 58.165000  7.390000 58.365000  7.590000 ;
        RECT 58.165000  7.820000 58.365000  8.020000 ;
        RECT 58.165000  8.250000 58.365000  8.450000 ;
        RECT 58.165000  8.680000 58.365000  8.880000 ;
        RECT 58.165000  9.110000 58.365000  9.310000 ;
        RECT 58.165000  9.540000 58.365000  9.740000 ;
        RECT 58.165000  9.970000 58.365000 10.170000 ;
        RECT 58.165000 10.400000 58.365000 10.600000 ;
        RECT 58.165000 10.830000 58.365000 11.030000 ;
        RECT 58.165000 11.260000 58.365000 11.460000 ;
        RECT 58.570000  6.960000 58.770000  7.160000 ;
        RECT 58.570000  7.390000 58.770000  7.590000 ;
        RECT 58.570000  7.820000 58.770000  8.020000 ;
        RECT 58.570000  8.250000 58.770000  8.450000 ;
        RECT 58.570000  8.680000 58.770000  8.880000 ;
        RECT 58.570000  9.110000 58.770000  9.310000 ;
        RECT 58.570000  9.540000 58.770000  9.740000 ;
        RECT 58.570000  9.970000 58.770000 10.170000 ;
        RECT 58.570000 10.400000 58.770000 10.600000 ;
        RECT 58.570000 10.830000 58.770000 11.030000 ;
        RECT 58.570000 11.260000 58.770000 11.460000 ;
        RECT 58.975000  6.960000 59.175000  7.160000 ;
        RECT 58.975000  7.390000 59.175000  7.590000 ;
        RECT 58.975000  7.820000 59.175000  8.020000 ;
        RECT 58.975000  8.250000 59.175000  8.450000 ;
        RECT 58.975000  8.680000 59.175000  8.880000 ;
        RECT 58.975000  9.110000 59.175000  9.310000 ;
        RECT 58.975000  9.540000 59.175000  9.740000 ;
        RECT 58.975000  9.970000 59.175000 10.170000 ;
        RECT 58.975000 10.400000 59.175000 10.600000 ;
        RECT 58.975000 10.830000 59.175000 11.030000 ;
        RECT 58.975000 11.260000 59.175000 11.460000 ;
        RECT 59.380000  6.960000 59.580000  7.160000 ;
        RECT 59.380000  7.390000 59.580000  7.590000 ;
        RECT 59.380000  7.820000 59.580000  8.020000 ;
        RECT 59.380000  8.250000 59.580000  8.450000 ;
        RECT 59.380000  8.680000 59.580000  8.880000 ;
        RECT 59.380000  9.110000 59.580000  9.310000 ;
        RECT 59.380000  9.540000 59.580000  9.740000 ;
        RECT 59.380000  9.970000 59.580000 10.170000 ;
        RECT 59.380000 10.400000 59.580000 10.600000 ;
        RECT 59.380000 10.830000 59.580000 11.030000 ;
        RECT 59.380000 11.260000 59.580000 11.460000 ;
        RECT 59.785000  6.960000 59.985000  7.160000 ;
        RECT 59.785000  7.390000 59.985000  7.590000 ;
        RECT 59.785000  7.820000 59.985000  8.020000 ;
        RECT 59.785000  8.250000 59.985000  8.450000 ;
        RECT 59.785000  8.680000 59.985000  8.880000 ;
        RECT 59.785000  9.110000 59.985000  9.310000 ;
        RECT 59.785000  9.540000 59.985000  9.740000 ;
        RECT 59.785000  9.970000 59.985000 10.170000 ;
        RECT 59.785000 10.400000 59.985000 10.600000 ;
        RECT 59.785000 10.830000 59.985000 11.030000 ;
        RECT 59.785000 11.260000 59.985000 11.460000 ;
        RECT 60.190000  6.960000 60.390000  7.160000 ;
        RECT 60.190000  7.390000 60.390000  7.590000 ;
        RECT 60.190000  7.820000 60.390000  8.020000 ;
        RECT 60.190000  8.250000 60.390000  8.450000 ;
        RECT 60.190000  8.680000 60.390000  8.880000 ;
        RECT 60.190000  9.110000 60.390000  9.310000 ;
        RECT 60.190000  9.540000 60.390000  9.740000 ;
        RECT 60.190000  9.970000 60.390000 10.170000 ;
        RECT 60.190000 10.400000 60.390000 10.600000 ;
        RECT 60.190000 10.830000 60.390000 11.030000 ;
        RECT 60.190000 11.260000 60.390000 11.460000 ;
        RECT 60.595000  6.960000 60.795000  7.160000 ;
        RECT 60.595000  7.390000 60.795000  7.590000 ;
        RECT 60.595000  7.820000 60.795000  8.020000 ;
        RECT 60.595000  8.250000 60.795000  8.450000 ;
        RECT 60.595000  8.680000 60.795000  8.880000 ;
        RECT 60.595000  9.110000 60.795000  9.310000 ;
        RECT 60.595000  9.540000 60.795000  9.740000 ;
        RECT 60.595000  9.970000 60.795000 10.170000 ;
        RECT 60.595000 10.400000 60.795000 10.600000 ;
        RECT 60.595000 10.830000 60.795000 11.030000 ;
        RECT 60.595000 11.260000 60.795000 11.460000 ;
        RECT 61.000000  6.960000 61.200000  7.160000 ;
        RECT 61.000000  7.390000 61.200000  7.590000 ;
        RECT 61.000000  7.820000 61.200000  8.020000 ;
        RECT 61.000000  8.250000 61.200000  8.450000 ;
        RECT 61.000000  8.680000 61.200000  8.880000 ;
        RECT 61.000000  9.110000 61.200000  9.310000 ;
        RECT 61.000000  9.540000 61.200000  9.740000 ;
        RECT 61.000000  9.970000 61.200000 10.170000 ;
        RECT 61.000000 10.400000 61.200000 10.600000 ;
        RECT 61.000000 10.830000 61.200000 11.030000 ;
        RECT 61.000000 11.260000 61.200000 11.460000 ;
        RECT 61.405000  6.960000 61.605000  7.160000 ;
        RECT 61.405000  7.390000 61.605000  7.590000 ;
        RECT 61.405000  7.820000 61.605000  8.020000 ;
        RECT 61.405000  8.250000 61.605000  8.450000 ;
        RECT 61.405000  8.680000 61.605000  8.880000 ;
        RECT 61.405000  9.110000 61.605000  9.310000 ;
        RECT 61.405000  9.540000 61.605000  9.740000 ;
        RECT 61.405000  9.970000 61.605000 10.170000 ;
        RECT 61.405000 10.400000 61.605000 10.600000 ;
        RECT 61.405000 10.830000 61.605000 11.030000 ;
        RECT 61.405000 11.260000 61.605000 11.460000 ;
        RECT 61.810000  6.960000 62.010000  7.160000 ;
        RECT 61.810000  7.390000 62.010000  7.590000 ;
        RECT 61.810000  7.820000 62.010000  8.020000 ;
        RECT 61.810000  8.250000 62.010000  8.450000 ;
        RECT 61.810000  8.680000 62.010000  8.880000 ;
        RECT 61.810000  9.110000 62.010000  9.310000 ;
        RECT 61.810000  9.540000 62.010000  9.740000 ;
        RECT 61.810000  9.970000 62.010000 10.170000 ;
        RECT 61.810000 10.400000 62.010000 10.600000 ;
        RECT 61.810000 10.830000 62.010000 11.030000 ;
        RECT 61.810000 11.260000 62.010000 11.460000 ;
        RECT 62.215000  6.960000 62.415000  7.160000 ;
        RECT 62.215000  7.390000 62.415000  7.590000 ;
        RECT 62.215000  7.820000 62.415000  8.020000 ;
        RECT 62.215000  8.250000 62.415000  8.450000 ;
        RECT 62.215000  8.680000 62.415000  8.880000 ;
        RECT 62.215000  9.110000 62.415000  9.310000 ;
        RECT 62.215000  9.540000 62.415000  9.740000 ;
        RECT 62.215000  9.970000 62.415000 10.170000 ;
        RECT 62.215000 10.400000 62.415000 10.600000 ;
        RECT 62.215000 10.830000 62.415000 11.030000 ;
        RECT 62.215000 11.260000 62.415000 11.460000 ;
        RECT 62.620000  6.960000 62.820000  7.160000 ;
        RECT 62.620000  7.390000 62.820000  7.590000 ;
        RECT 62.620000  7.820000 62.820000  8.020000 ;
        RECT 62.620000  8.250000 62.820000  8.450000 ;
        RECT 62.620000  8.680000 62.820000  8.880000 ;
        RECT 62.620000  9.110000 62.820000  9.310000 ;
        RECT 62.620000  9.540000 62.820000  9.740000 ;
        RECT 62.620000  9.970000 62.820000 10.170000 ;
        RECT 62.620000 10.400000 62.820000 10.600000 ;
        RECT 62.620000 10.830000 62.820000 11.030000 ;
        RECT 62.620000 11.260000 62.820000 11.460000 ;
        RECT 63.025000  6.960000 63.225000  7.160000 ;
        RECT 63.025000  7.390000 63.225000  7.590000 ;
        RECT 63.025000  7.820000 63.225000  8.020000 ;
        RECT 63.025000  8.250000 63.225000  8.450000 ;
        RECT 63.025000  8.680000 63.225000  8.880000 ;
        RECT 63.025000  9.110000 63.225000  9.310000 ;
        RECT 63.025000  9.540000 63.225000  9.740000 ;
        RECT 63.025000  9.970000 63.225000 10.170000 ;
        RECT 63.025000 10.400000 63.225000 10.600000 ;
        RECT 63.025000 10.830000 63.225000 11.030000 ;
        RECT 63.025000 11.260000 63.225000 11.460000 ;
        RECT 63.430000  6.960000 63.630000  7.160000 ;
        RECT 63.430000  7.390000 63.630000  7.590000 ;
        RECT 63.430000  7.820000 63.630000  8.020000 ;
        RECT 63.430000  8.250000 63.630000  8.450000 ;
        RECT 63.430000  8.680000 63.630000  8.880000 ;
        RECT 63.430000  9.110000 63.630000  9.310000 ;
        RECT 63.430000  9.540000 63.630000  9.740000 ;
        RECT 63.430000  9.970000 63.630000 10.170000 ;
        RECT 63.430000 10.400000 63.630000 10.600000 ;
        RECT 63.430000 10.830000 63.630000 11.030000 ;
        RECT 63.430000 11.260000 63.630000 11.460000 ;
        RECT 63.835000  6.960000 64.035000  7.160000 ;
        RECT 63.835000  7.390000 64.035000  7.590000 ;
        RECT 63.835000  7.820000 64.035000  8.020000 ;
        RECT 63.835000  8.250000 64.035000  8.450000 ;
        RECT 63.835000  8.680000 64.035000  8.880000 ;
        RECT 63.835000  9.110000 64.035000  9.310000 ;
        RECT 63.835000  9.540000 64.035000  9.740000 ;
        RECT 63.835000  9.970000 64.035000 10.170000 ;
        RECT 63.835000 10.400000 64.035000 10.600000 ;
        RECT 63.835000 10.830000 64.035000 11.030000 ;
        RECT 63.835000 11.260000 64.035000 11.460000 ;
        RECT 64.240000  6.960000 64.440000  7.160000 ;
        RECT 64.240000  7.390000 64.440000  7.590000 ;
        RECT 64.240000  7.820000 64.440000  8.020000 ;
        RECT 64.240000  8.250000 64.440000  8.450000 ;
        RECT 64.240000  8.680000 64.440000  8.880000 ;
        RECT 64.240000  9.110000 64.440000  9.310000 ;
        RECT 64.240000  9.540000 64.440000  9.740000 ;
        RECT 64.240000  9.970000 64.440000 10.170000 ;
        RECT 64.240000 10.400000 64.440000 10.600000 ;
        RECT 64.240000 10.830000 64.440000 11.030000 ;
        RECT 64.240000 11.260000 64.440000 11.460000 ;
        RECT 64.645000  6.960000 64.845000  7.160000 ;
        RECT 64.645000  7.390000 64.845000  7.590000 ;
        RECT 64.645000  7.820000 64.845000  8.020000 ;
        RECT 64.645000  8.250000 64.845000  8.450000 ;
        RECT 64.645000  8.680000 64.845000  8.880000 ;
        RECT 64.645000  9.110000 64.845000  9.310000 ;
        RECT 64.645000  9.540000 64.845000  9.740000 ;
        RECT 64.645000  9.970000 64.845000 10.170000 ;
        RECT 64.645000 10.400000 64.845000 10.600000 ;
        RECT 64.645000 10.830000 64.845000 11.030000 ;
        RECT 64.645000 11.260000 64.845000 11.460000 ;
        RECT 65.050000  6.960000 65.250000  7.160000 ;
        RECT 65.050000  7.390000 65.250000  7.590000 ;
        RECT 65.050000  7.820000 65.250000  8.020000 ;
        RECT 65.050000  8.250000 65.250000  8.450000 ;
        RECT 65.050000  8.680000 65.250000  8.880000 ;
        RECT 65.050000  9.110000 65.250000  9.310000 ;
        RECT 65.050000  9.540000 65.250000  9.740000 ;
        RECT 65.050000  9.970000 65.250000 10.170000 ;
        RECT 65.050000 10.400000 65.250000 10.600000 ;
        RECT 65.050000 10.830000 65.250000 11.030000 ;
        RECT 65.050000 11.260000 65.250000 11.460000 ;
        RECT 65.455000  6.960000 65.655000  7.160000 ;
        RECT 65.455000  7.390000 65.655000  7.590000 ;
        RECT 65.455000  7.820000 65.655000  8.020000 ;
        RECT 65.455000  8.250000 65.655000  8.450000 ;
        RECT 65.455000  8.680000 65.655000  8.880000 ;
        RECT 65.455000  9.110000 65.655000  9.310000 ;
        RECT 65.455000  9.540000 65.655000  9.740000 ;
        RECT 65.455000  9.970000 65.655000 10.170000 ;
        RECT 65.455000 10.400000 65.655000 10.600000 ;
        RECT 65.455000 10.830000 65.655000 11.030000 ;
        RECT 65.455000 11.260000 65.655000 11.460000 ;
        RECT 65.860000  6.960000 66.060000  7.160000 ;
        RECT 65.860000  7.390000 66.060000  7.590000 ;
        RECT 65.860000  7.820000 66.060000  8.020000 ;
        RECT 65.860000  8.250000 66.060000  8.450000 ;
        RECT 65.860000  8.680000 66.060000  8.880000 ;
        RECT 65.860000  9.110000 66.060000  9.310000 ;
        RECT 65.860000  9.540000 66.060000  9.740000 ;
        RECT 65.860000  9.970000 66.060000 10.170000 ;
        RECT 65.860000 10.400000 66.060000 10.600000 ;
        RECT 65.860000 10.830000 66.060000 11.030000 ;
        RECT 65.860000 11.260000 66.060000 11.460000 ;
        RECT 66.265000  6.960000 66.465000  7.160000 ;
        RECT 66.265000  7.390000 66.465000  7.590000 ;
        RECT 66.265000  7.820000 66.465000  8.020000 ;
        RECT 66.265000  8.250000 66.465000  8.450000 ;
        RECT 66.265000  8.680000 66.465000  8.880000 ;
        RECT 66.265000  9.110000 66.465000  9.310000 ;
        RECT 66.265000  9.540000 66.465000  9.740000 ;
        RECT 66.265000  9.970000 66.465000 10.170000 ;
        RECT 66.265000 10.400000 66.465000 10.600000 ;
        RECT 66.265000 10.830000 66.465000 11.030000 ;
        RECT 66.265000 11.260000 66.465000 11.460000 ;
        RECT 66.670000  6.960000 66.870000  7.160000 ;
        RECT 66.670000  7.390000 66.870000  7.590000 ;
        RECT 66.670000  7.820000 66.870000  8.020000 ;
        RECT 66.670000  8.250000 66.870000  8.450000 ;
        RECT 66.670000  8.680000 66.870000  8.880000 ;
        RECT 66.670000  9.110000 66.870000  9.310000 ;
        RECT 66.670000  9.540000 66.870000  9.740000 ;
        RECT 66.670000  9.970000 66.870000 10.170000 ;
        RECT 66.670000 10.400000 66.870000 10.600000 ;
        RECT 66.670000 10.830000 66.870000 11.030000 ;
        RECT 66.670000 11.260000 66.870000 11.460000 ;
        RECT 67.075000  6.960000 67.275000  7.160000 ;
        RECT 67.075000  7.390000 67.275000  7.590000 ;
        RECT 67.075000  7.820000 67.275000  8.020000 ;
        RECT 67.075000  8.250000 67.275000  8.450000 ;
        RECT 67.075000  8.680000 67.275000  8.880000 ;
        RECT 67.075000  9.110000 67.275000  9.310000 ;
        RECT 67.075000  9.540000 67.275000  9.740000 ;
        RECT 67.075000  9.970000 67.275000 10.170000 ;
        RECT 67.075000 10.400000 67.275000 10.600000 ;
        RECT 67.075000 10.830000 67.275000 11.030000 ;
        RECT 67.075000 11.260000 67.275000 11.460000 ;
        RECT 67.480000  6.960000 67.680000  7.160000 ;
        RECT 67.480000  7.390000 67.680000  7.590000 ;
        RECT 67.480000  7.820000 67.680000  8.020000 ;
        RECT 67.480000  8.250000 67.680000  8.450000 ;
        RECT 67.480000  8.680000 67.680000  8.880000 ;
        RECT 67.480000  9.110000 67.680000  9.310000 ;
        RECT 67.480000  9.540000 67.680000  9.740000 ;
        RECT 67.480000  9.970000 67.680000 10.170000 ;
        RECT 67.480000 10.400000 67.680000 10.600000 ;
        RECT 67.480000 10.830000 67.680000 11.030000 ;
        RECT 67.480000 11.260000 67.680000 11.460000 ;
        RECT 67.885000  6.960000 68.085000  7.160000 ;
        RECT 67.885000  7.390000 68.085000  7.590000 ;
        RECT 67.885000  7.820000 68.085000  8.020000 ;
        RECT 67.885000  8.250000 68.085000  8.450000 ;
        RECT 67.885000  8.680000 68.085000  8.880000 ;
        RECT 67.885000  9.110000 68.085000  9.310000 ;
        RECT 67.885000  9.540000 68.085000  9.740000 ;
        RECT 67.885000  9.970000 68.085000 10.170000 ;
        RECT 67.885000 10.400000 68.085000 10.600000 ;
        RECT 67.885000 10.830000 68.085000 11.030000 ;
        RECT 67.885000 11.260000 68.085000 11.460000 ;
        RECT 68.290000  6.960000 68.490000  7.160000 ;
        RECT 68.290000  7.390000 68.490000  7.590000 ;
        RECT 68.290000  7.820000 68.490000  8.020000 ;
        RECT 68.290000  8.250000 68.490000  8.450000 ;
        RECT 68.290000  8.680000 68.490000  8.880000 ;
        RECT 68.290000  9.110000 68.490000  9.310000 ;
        RECT 68.290000  9.540000 68.490000  9.740000 ;
        RECT 68.290000  9.970000 68.490000 10.170000 ;
        RECT 68.290000 10.400000 68.490000 10.600000 ;
        RECT 68.290000 10.830000 68.490000 11.030000 ;
        RECT 68.290000 11.260000 68.490000 11.460000 ;
        RECT 68.695000  6.960000 68.895000  7.160000 ;
        RECT 68.695000  7.390000 68.895000  7.590000 ;
        RECT 68.695000  7.820000 68.895000  8.020000 ;
        RECT 68.695000  8.250000 68.895000  8.450000 ;
        RECT 68.695000  8.680000 68.895000  8.880000 ;
        RECT 68.695000  9.110000 68.895000  9.310000 ;
        RECT 68.695000  9.540000 68.895000  9.740000 ;
        RECT 68.695000  9.970000 68.895000 10.170000 ;
        RECT 68.695000 10.400000 68.895000 10.600000 ;
        RECT 68.695000 10.830000 68.895000 11.030000 ;
        RECT 68.695000 11.260000 68.895000 11.460000 ;
        RECT 69.100000  6.960000 69.300000  7.160000 ;
        RECT 69.100000  7.390000 69.300000  7.590000 ;
        RECT 69.100000  7.820000 69.300000  8.020000 ;
        RECT 69.100000  8.250000 69.300000  8.450000 ;
        RECT 69.100000  8.680000 69.300000  8.880000 ;
        RECT 69.100000  9.110000 69.300000  9.310000 ;
        RECT 69.100000  9.540000 69.300000  9.740000 ;
        RECT 69.100000  9.970000 69.300000 10.170000 ;
        RECT 69.100000 10.400000 69.300000 10.600000 ;
        RECT 69.100000 10.830000 69.300000 11.030000 ;
        RECT 69.100000 11.260000 69.300000 11.460000 ;
        RECT 69.505000  6.960000 69.705000  7.160000 ;
        RECT 69.505000  7.390000 69.705000  7.590000 ;
        RECT 69.505000  7.820000 69.705000  8.020000 ;
        RECT 69.505000  8.250000 69.705000  8.450000 ;
        RECT 69.505000  8.680000 69.705000  8.880000 ;
        RECT 69.505000  9.110000 69.705000  9.310000 ;
        RECT 69.505000  9.540000 69.705000  9.740000 ;
        RECT 69.505000  9.970000 69.705000 10.170000 ;
        RECT 69.505000 10.400000 69.705000 10.600000 ;
        RECT 69.505000 10.830000 69.705000 11.030000 ;
        RECT 69.505000 11.260000 69.705000 11.460000 ;
        RECT 69.910000  6.960000 70.110000  7.160000 ;
        RECT 69.910000  7.390000 70.110000  7.590000 ;
        RECT 69.910000  7.820000 70.110000  8.020000 ;
        RECT 69.910000  8.250000 70.110000  8.450000 ;
        RECT 69.910000  8.680000 70.110000  8.880000 ;
        RECT 69.910000  9.110000 70.110000  9.310000 ;
        RECT 69.910000  9.540000 70.110000  9.740000 ;
        RECT 69.910000  9.970000 70.110000 10.170000 ;
        RECT 69.910000 10.400000 70.110000 10.600000 ;
        RECT 69.910000 10.830000 70.110000 11.030000 ;
        RECT 69.910000 11.260000 70.110000 11.460000 ;
        RECT 70.315000  6.960000 70.515000  7.160000 ;
        RECT 70.315000  7.390000 70.515000  7.590000 ;
        RECT 70.315000  7.820000 70.515000  8.020000 ;
        RECT 70.315000  8.250000 70.515000  8.450000 ;
        RECT 70.315000  8.680000 70.515000  8.880000 ;
        RECT 70.315000  9.110000 70.515000  9.310000 ;
        RECT 70.315000  9.540000 70.515000  9.740000 ;
        RECT 70.315000  9.970000 70.515000 10.170000 ;
        RECT 70.315000 10.400000 70.515000 10.600000 ;
        RECT 70.315000 10.830000 70.515000 11.030000 ;
        RECT 70.315000 11.260000 70.515000 11.460000 ;
        RECT 70.720000  6.960000 70.920000  7.160000 ;
        RECT 70.720000  7.390000 70.920000  7.590000 ;
        RECT 70.720000  7.820000 70.920000  8.020000 ;
        RECT 70.720000  8.250000 70.920000  8.450000 ;
        RECT 70.720000  8.680000 70.920000  8.880000 ;
        RECT 70.720000  9.110000 70.920000  9.310000 ;
        RECT 70.720000  9.540000 70.920000  9.740000 ;
        RECT 70.720000  9.970000 70.920000 10.170000 ;
        RECT 70.720000 10.400000 70.920000 10.600000 ;
        RECT 70.720000 10.830000 70.920000 11.030000 ;
        RECT 70.720000 11.260000 70.920000 11.460000 ;
        RECT 71.125000  6.960000 71.325000  7.160000 ;
        RECT 71.125000  7.390000 71.325000  7.590000 ;
        RECT 71.125000  7.820000 71.325000  8.020000 ;
        RECT 71.125000  8.250000 71.325000  8.450000 ;
        RECT 71.125000  8.680000 71.325000  8.880000 ;
        RECT 71.125000  9.110000 71.325000  9.310000 ;
        RECT 71.125000  9.540000 71.325000  9.740000 ;
        RECT 71.125000  9.970000 71.325000 10.170000 ;
        RECT 71.125000 10.400000 71.325000 10.600000 ;
        RECT 71.125000 10.830000 71.325000 11.030000 ;
        RECT 71.125000 11.260000 71.325000 11.460000 ;
        RECT 71.530000  6.960000 71.730000  7.160000 ;
        RECT 71.530000  7.390000 71.730000  7.590000 ;
        RECT 71.530000  7.820000 71.730000  8.020000 ;
        RECT 71.530000  8.250000 71.730000  8.450000 ;
        RECT 71.530000  8.680000 71.730000  8.880000 ;
        RECT 71.530000  9.110000 71.730000  9.310000 ;
        RECT 71.530000  9.540000 71.730000  9.740000 ;
        RECT 71.530000  9.970000 71.730000 10.170000 ;
        RECT 71.530000 10.400000 71.730000 10.600000 ;
        RECT 71.530000 10.830000 71.730000 11.030000 ;
        RECT 71.530000 11.260000 71.730000 11.460000 ;
        RECT 71.935000  6.960000 72.135000  7.160000 ;
        RECT 71.935000  7.390000 72.135000  7.590000 ;
        RECT 71.935000  7.820000 72.135000  8.020000 ;
        RECT 71.935000  8.250000 72.135000  8.450000 ;
        RECT 71.935000  8.680000 72.135000  8.880000 ;
        RECT 71.935000  9.110000 72.135000  9.310000 ;
        RECT 71.935000  9.540000 72.135000  9.740000 ;
        RECT 71.935000  9.970000 72.135000 10.170000 ;
        RECT 71.935000 10.400000 72.135000 10.600000 ;
        RECT 71.935000 10.830000 72.135000 11.030000 ;
        RECT 71.935000 11.260000 72.135000 11.460000 ;
        RECT 72.340000  6.960000 72.540000  7.160000 ;
        RECT 72.340000  7.390000 72.540000  7.590000 ;
        RECT 72.340000  7.820000 72.540000  8.020000 ;
        RECT 72.340000  8.250000 72.540000  8.450000 ;
        RECT 72.340000  8.680000 72.540000  8.880000 ;
        RECT 72.340000  9.110000 72.540000  9.310000 ;
        RECT 72.340000  9.540000 72.540000  9.740000 ;
        RECT 72.340000  9.970000 72.540000 10.170000 ;
        RECT 72.340000 10.400000 72.540000 10.600000 ;
        RECT 72.340000 10.830000 72.540000 11.030000 ;
        RECT 72.340000 11.260000 72.540000 11.460000 ;
        RECT 72.745000  6.960000 72.945000  7.160000 ;
        RECT 72.745000  7.390000 72.945000  7.590000 ;
        RECT 72.745000  7.820000 72.945000  8.020000 ;
        RECT 72.745000  8.250000 72.945000  8.450000 ;
        RECT 72.745000  8.680000 72.945000  8.880000 ;
        RECT 72.745000  9.110000 72.945000  9.310000 ;
        RECT 72.745000  9.540000 72.945000  9.740000 ;
        RECT 72.745000  9.970000 72.945000 10.170000 ;
        RECT 72.745000 10.400000 72.945000 10.600000 ;
        RECT 72.745000 10.830000 72.945000 11.030000 ;
        RECT 72.745000 11.260000 72.945000 11.460000 ;
        RECT 73.150000  6.960000 73.350000  7.160000 ;
        RECT 73.150000  7.390000 73.350000  7.590000 ;
        RECT 73.150000  7.820000 73.350000  8.020000 ;
        RECT 73.150000  8.250000 73.350000  8.450000 ;
        RECT 73.150000  8.680000 73.350000  8.880000 ;
        RECT 73.150000  9.110000 73.350000  9.310000 ;
        RECT 73.150000  9.540000 73.350000  9.740000 ;
        RECT 73.150000  9.970000 73.350000 10.170000 ;
        RECT 73.150000 10.400000 73.350000 10.600000 ;
        RECT 73.150000 10.830000 73.350000 11.030000 ;
        RECT 73.150000 11.260000 73.350000 11.460000 ;
        RECT 73.555000  6.960000 73.755000  7.160000 ;
        RECT 73.555000  7.390000 73.755000  7.590000 ;
        RECT 73.555000  7.820000 73.755000  8.020000 ;
        RECT 73.555000  8.250000 73.755000  8.450000 ;
        RECT 73.555000  8.680000 73.755000  8.880000 ;
        RECT 73.555000  9.110000 73.755000  9.310000 ;
        RECT 73.555000  9.540000 73.755000  9.740000 ;
        RECT 73.555000  9.970000 73.755000 10.170000 ;
        RECT 73.555000 10.400000 73.755000 10.600000 ;
        RECT 73.555000 10.830000 73.755000 11.030000 ;
        RECT 73.555000 11.260000 73.755000 11.460000 ;
        RECT 73.960000  6.960000 74.160000  7.160000 ;
        RECT 73.960000  7.390000 74.160000  7.590000 ;
        RECT 73.960000  7.820000 74.160000  8.020000 ;
        RECT 73.960000  8.250000 74.160000  8.450000 ;
        RECT 73.960000  8.680000 74.160000  8.880000 ;
        RECT 73.960000  9.110000 74.160000  9.310000 ;
        RECT 73.960000  9.540000 74.160000  9.740000 ;
        RECT 73.960000  9.970000 74.160000 10.170000 ;
        RECT 73.960000 10.400000 74.160000 10.600000 ;
        RECT 73.960000 10.830000 74.160000 11.030000 ;
        RECT 73.960000 11.260000 74.160000 11.460000 ;
        RECT 74.365000  6.960000 74.565000  7.160000 ;
        RECT 74.365000  7.390000 74.565000  7.590000 ;
        RECT 74.365000  7.820000 74.565000  8.020000 ;
        RECT 74.365000  8.250000 74.565000  8.450000 ;
        RECT 74.365000  8.680000 74.565000  8.880000 ;
        RECT 74.365000  9.110000 74.565000  9.310000 ;
        RECT 74.365000  9.540000 74.565000  9.740000 ;
        RECT 74.365000  9.970000 74.565000 10.170000 ;
        RECT 74.365000 10.400000 74.565000 10.600000 ;
        RECT 74.365000 10.830000 74.565000 11.030000 ;
        RECT 74.365000 11.260000 74.565000 11.460000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
  END
END sky130_fd_io__overlay_vccd_lvc


MACRO sky130_fd_io__overlay_vssio_hvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT  0.495000 173.155000 13.500000 195.340000 ;
        RECT  0.495000 195.340000 13.500000 195.490000 ;
        RECT  0.495000 195.490000 13.650000 195.640000 ;
        RECT  0.495000 195.640000 13.800000 195.790000 ;
        RECT  0.495000 195.790000 13.950000 195.940000 ;
        RECT  0.495000 195.940000 14.100000 196.090000 ;
        RECT  0.495000 196.090000 14.250000 196.240000 ;
        RECT  0.495000 196.240000 14.400000 196.390000 ;
        RECT  0.495000 196.390000 14.550000 196.540000 ;
        RECT  0.495000 196.540000 14.700000 196.690000 ;
        RECT  0.495000 196.690000 14.850000 196.840000 ;
        RECT  0.495000 196.840000 15.000000 196.990000 ;
        RECT  0.495000 196.990000 15.150000 197.140000 ;
        RECT  0.495000 197.140000 15.300000 197.175000 ;
        RECT  0.495000 197.175000 74.290000 200.000000 ;
        RECT 59.700000 197.110000 74.290000 197.175000 ;
        RECT 59.850000 196.960000 74.290000 197.110000 ;
        RECT 60.000000 196.810000 74.290000 196.960000 ;
        RECT 60.150000 196.660000 74.290000 196.810000 ;
        RECT 60.300000 196.510000 74.290000 196.660000 ;
        RECT 60.450000 196.360000 74.290000 196.510000 ;
        RECT 60.600000 196.210000 74.290000 196.360000 ;
        RECT 60.750000 196.060000 74.290000 196.210000 ;
        RECT 60.900000 195.910000 74.290000 196.060000 ;
        RECT 61.050000 195.760000 74.290000 195.910000 ;
        RECT 61.200000 195.610000 74.290000 195.760000 ;
        RECT 61.350000 195.460000 74.290000 195.610000 ;
        RECT 61.500000 173.320000 74.290000 195.310000 ;
        RECT 61.500000 195.310000 74.290000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495000 25.840000 24.395000 30.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 25.840000 74.290000 30.480000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000  1.270000 175.930000 ;
        RECT 0.000000 175.930000 13.475000 199.920000 ;
        RECT 0.000000 199.920000  1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 24.370000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.595000 196.230000 14.255000 196.970000 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.630000 197.170000 61.325000 199.930000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.680000 196.230000 61.340000 196.970000 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.505000 175.930000 75.000000 199.920000 ;
        RECT 73.730000 175.785000 75.000000 175.930000 ;
        RECT 73.730000 199.920000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.585000  25.910000  0.785000  26.110000 ;
        RECT  0.585000  26.340000  0.785000  26.540000 ;
        RECT  0.585000  26.770000  0.785000  26.970000 ;
        RECT  0.585000  27.200000  0.785000  27.400000 ;
        RECT  0.585000  27.630000  0.785000  27.830000 ;
        RECT  0.585000  28.060000  0.785000  28.260000 ;
        RECT  0.585000  28.490000  0.785000  28.690000 ;
        RECT  0.585000  28.920000  0.785000  29.120000 ;
        RECT  0.585000  29.350000  0.785000  29.550000 ;
        RECT  0.585000  29.780000  0.785000  29.980000 ;
        RECT  0.585000  30.210000  0.785000  30.410000 ;
        RECT  0.685000 175.995000  0.885000 176.195000 ;
        RECT  0.685000 176.395000  0.885000 176.595000 ;
        RECT  0.685000 176.795000  0.885000 176.995000 ;
        RECT  0.685000 177.195000  0.885000 177.395000 ;
        RECT  0.685000 177.595000  0.885000 177.795000 ;
        RECT  0.685000 177.995000  0.885000 178.195000 ;
        RECT  0.685000 178.395000  0.885000 178.595000 ;
        RECT  0.685000 178.795000  0.885000 178.995000 ;
        RECT  0.685000 179.195000  0.885000 179.395000 ;
        RECT  0.685000 179.595000  0.885000 179.795000 ;
        RECT  0.685000 179.995000  0.885000 180.195000 ;
        RECT  0.685000 180.395000  0.885000 180.595000 ;
        RECT  0.685000 180.795000  0.885000 180.995000 ;
        RECT  0.685000 181.195000  0.885000 181.395000 ;
        RECT  0.685000 181.595000  0.885000 181.795000 ;
        RECT  0.685000 181.995000  0.885000 182.195000 ;
        RECT  0.685000 182.395000  0.885000 182.595000 ;
        RECT  0.685000 182.795000  0.885000 182.995000 ;
        RECT  0.685000 183.195000  0.885000 183.395000 ;
        RECT  0.685000 183.595000  0.885000 183.795000 ;
        RECT  0.685000 183.995000  0.885000 184.195000 ;
        RECT  0.685000 184.395000  0.885000 184.595000 ;
        RECT  0.685000 184.795000  0.885000 184.995000 ;
        RECT  0.685000 185.195000  0.885000 185.395000 ;
        RECT  0.685000 185.595000  0.885000 185.795000 ;
        RECT  0.685000 185.995000  0.885000 186.195000 ;
        RECT  0.685000 186.395000  0.885000 186.595000 ;
        RECT  0.685000 186.795000  0.885000 186.995000 ;
        RECT  0.685000 187.195000  0.885000 187.395000 ;
        RECT  0.685000 187.595000  0.885000 187.795000 ;
        RECT  0.685000 187.995000  0.885000 188.195000 ;
        RECT  0.685000 188.395000  0.885000 188.595000 ;
        RECT  0.685000 188.795000  0.885000 188.995000 ;
        RECT  0.685000 189.195000  0.885000 189.395000 ;
        RECT  0.685000 189.595000  0.885000 189.795000 ;
        RECT  0.685000 189.995000  0.885000 190.195000 ;
        RECT  0.685000 190.395000  0.885000 190.595000 ;
        RECT  0.685000 190.795000  0.885000 190.995000 ;
        RECT  0.685000 191.195000  0.885000 191.395000 ;
        RECT  0.685000 191.595000  0.885000 191.795000 ;
        RECT  0.685000 191.995000  0.885000 192.195000 ;
        RECT  0.685000 192.395000  0.885000 192.595000 ;
        RECT  0.685000 192.795000  0.885000 192.995000 ;
        RECT  0.685000 193.195000  0.885000 193.395000 ;
        RECT  0.685000 193.595000  0.885000 193.795000 ;
        RECT  0.685000 193.995000  0.885000 194.195000 ;
        RECT  0.685000 194.395000  0.885000 194.595000 ;
        RECT  0.685000 194.795000  0.885000 194.995000 ;
        RECT  0.685000 195.200000  0.885000 195.400000 ;
        RECT  0.685000 195.605000  0.885000 195.805000 ;
        RECT  0.685000 196.010000  0.885000 196.210000 ;
        RECT  0.685000 196.415000  0.885000 196.615000 ;
        RECT  0.685000 196.820000  0.885000 197.020000 ;
        RECT  0.685000 197.225000  0.885000 197.425000 ;
        RECT  0.685000 197.630000  0.885000 197.830000 ;
        RECT  0.685000 198.035000  0.885000 198.235000 ;
        RECT  0.685000 198.440000  0.885000 198.640000 ;
        RECT  0.685000 198.845000  0.885000 199.045000 ;
        RECT  0.685000 199.250000  0.885000 199.450000 ;
        RECT  0.685000 199.655000  0.885000 199.855000 ;
        RECT  0.995000  25.910000  1.195000  26.110000 ;
        RECT  0.995000  26.340000  1.195000  26.540000 ;
        RECT  0.995000  26.770000  1.195000  26.970000 ;
        RECT  0.995000  27.200000  1.195000  27.400000 ;
        RECT  0.995000  27.630000  1.195000  27.830000 ;
        RECT  0.995000  28.060000  1.195000  28.260000 ;
        RECT  0.995000  28.490000  1.195000  28.690000 ;
        RECT  0.995000  28.920000  1.195000  29.120000 ;
        RECT  0.995000  29.350000  1.195000  29.550000 ;
        RECT  0.995000  29.780000  1.195000  29.980000 ;
        RECT  0.995000  30.210000  1.195000  30.410000 ;
        RECT  1.085000 175.995000  1.285000 176.195000 ;
        RECT  1.085000 176.395000  1.285000 176.595000 ;
        RECT  1.085000 176.795000  1.285000 176.995000 ;
        RECT  1.085000 177.195000  1.285000 177.395000 ;
        RECT  1.085000 177.595000  1.285000 177.795000 ;
        RECT  1.085000 177.995000  1.285000 178.195000 ;
        RECT  1.085000 178.395000  1.285000 178.595000 ;
        RECT  1.085000 178.795000  1.285000 178.995000 ;
        RECT  1.085000 179.195000  1.285000 179.395000 ;
        RECT  1.085000 179.595000  1.285000 179.795000 ;
        RECT  1.085000 179.995000  1.285000 180.195000 ;
        RECT  1.085000 180.395000  1.285000 180.595000 ;
        RECT  1.085000 180.795000  1.285000 180.995000 ;
        RECT  1.085000 181.195000  1.285000 181.395000 ;
        RECT  1.085000 181.595000  1.285000 181.795000 ;
        RECT  1.085000 181.995000  1.285000 182.195000 ;
        RECT  1.085000 182.395000  1.285000 182.595000 ;
        RECT  1.085000 182.795000  1.285000 182.995000 ;
        RECT  1.085000 183.195000  1.285000 183.395000 ;
        RECT  1.085000 183.595000  1.285000 183.795000 ;
        RECT  1.085000 183.995000  1.285000 184.195000 ;
        RECT  1.085000 184.395000  1.285000 184.595000 ;
        RECT  1.085000 184.795000  1.285000 184.995000 ;
        RECT  1.085000 185.195000  1.285000 185.395000 ;
        RECT  1.085000 185.595000  1.285000 185.795000 ;
        RECT  1.085000 185.995000  1.285000 186.195000 ;
        RECT  1.085000 186.395000  1.285000 186.595000 ;
        RECT  1.085000 186.795000  1.285000 186.995000 ;
        RECT  1.085000 187.195000  1.285000 187.395000 ;
        RECT  1.085000 187.595000  1.285000 187.795000 ;
        RECT  1.085000 187.995000  1.285000 188.195000 ;
        RECT  1.085000 188.395000  1.285000 188.595000 ;
        RECT  1.085000 188.795000  1.285000 188.995000 ;
        RECT  1.085000 189.195000  1.285000 189.395000 ;
        RECT  1.085000 189.595000  1.285000 189.795000 ;
        RECT  1.085000 189.995000  1.285000 190.195000 ;
        RECT  1.085000 190.395000  1.285000 190.595000 ;
        RECT  1.085000 190.795000  1.285000 190.995000 ;
        RECT  1.085000 191.195000  1.285000 191.395000 ;
        RECT  1.085000 191.595000  1.285000 191.795000 ;
        RECT  1.085000 191.995000  1.285000 192.195000 ;
        RECT  1.085000 192.395000  1.285000 192.595000 ;
        RECT  1.085000 192.795000  1.285000 192.995000 ;
        RECT  1.085000 193.195000  1.285000 193.395000 ;
        RECT  1.085000 193.595000  1.285000 193.795000 ;
        RECT  1.085000 193.995000  1.285000 194.195000 ;
        RECT  1.085000 194.395000  1.285000 194.595000 ;
        RECT  1.085000 194.795000  1.285000 194.995000 ;
        RECT  1.085000 195.200000  1.285000 195.400000 ;
        RECT  1.085000 195.605000  1.285000 195.805000 ;
        RECT  1.085000 196.010000  1.285000 196.210000 ;
        RECT  1.085000 196.415000  1.285000 196.615000 ;
        RECT  1.085000 196.820000  1.285000 197.020000 ;
        RECT  1.085000 197.225000  1.285000 197.425000 ;
        RECT  1.085000 197.630000  1.285000 197.830000 ;
        RECT  1.085000 198.035000  1.285000 198.235000 ;
        RECT  1.085000 198.440000  1.285000 198.640000 ;
        RECT  1.085000 198.845000  1.285000 199.045000 ;
        RECT  1.085000 199.250000  1.285000 199.450000 ;
        RECT  1.085000 199.655000  1.285000 199.855000 ;
        RECT  1.405000  25.910000  1.605000  26.110000 ;
        RECT  1.405000  26.340000  1.605000  26.540000 ;
        RECT  1.405000  26.770000  1.605000  26.970000 ;
        RECT  1.405000  27.200000  1.605000  27.400000 ;
        RECT  1.405000  27.630000  1.605000  27.830000 ;
        RECT  1.405000  28.060000  1.605000  28.260000 ;
        RECT  1.405000  28.490000  1.605000  28.690000 ;
        RECT  1.405000  28.920000  1.605000  29.120000 ;
        RECT  1.405000  29.350000  1.605000  29.550000 ;
        RECT  1.405000  29.780000  1.605000  29.980000 ;
        RECT  1.405000  30.210000  1.605000  30.410000 ;
        RECT  1.485000 175.995000  1.685000 176.195000 ;
        RECT  1.485000 176.395000  1.685000 176.595000 ;
        RECT  1.485000 176.795000  1.685000 176.995000 ;
        RECT  1.485000 177.195000  1.685000 177.395000 ;
        RECT  1.485000 177.595000  1.685000 177.795000 ;
        RECT  1.485000 177.995000  1.685000 178.195000 ;
        RECT  1.485000 178.395000  1.685000 178.595000 ;
        RECT  1.485000 178.795000  1.685000 178.995000 ;
        RECT  1.485000 179.195000  1.685000 179.395000 ;
        RECT  1.485000 179.595000  1.685000 179.795000 ;
        RECT  1.485000 179.995000  1.685000 180.195000 ;
        RECT  1.485000 180.395000  1.685000 180.595000 ;
        RECT  1.485000 180.795000  1.685000 180.995000 ;
        RECT  1.485000 181.195000  1.685000 181.395000 ;
        RECT  1.485000 181.595000  1.685000 181.795000 ;
        RECT  1.485000 181.995000  1.685000 182.195000 ;
        RECT  1.485000 182.395000  1.685000 182.595000 ;
        RECT  1.485000 182.795000  1.685000 182.995000 ;
        RECT  1.485000 183.195000  1.685000 183.395000 ;
        RECT  1.485000 183.595000  1.685000 183.795000 ;
        RECT  1.485000 183.995000  1.685000 184.195000 ;
        RECT  1.485000 184.395000  1.685000 184.595000 ;
        RECT  1.485000 184.795000  1.685000 184.995000 ;
        RECT  1.485000 185.195000  1.685000 185.395000 ;
        RECT  1.485000 185.595000  1.685000 185.795000 ;
        RECT  1.485000 185.995000  1.685000 186.195000 ;
        RECT  1.485000 186.395000  1.685000 186.595000 ;
        RECT  1.485000 186.795000  1.685000 186.995000 ;
        RECT  1.485000 187.195000  1.685000 187.395000 ;
        RECT  1.485000 187.595000  1.685000 187.795000 ;
        RECT  1.485000 187.995000  1.685000 188.195000 ;
        RECT  1.485000 188.395000  1.685000 188.595000 ;
        RECT  1.485000 188.795000  1.685000 188.995000 ;
        RECT  1.485000 189.195000  1.685000 189.395000 ;
        RECT  1.485000 189.595000  1.685000 189.795000 ;
        RECT  1.485000 189.995000  1.685000 190.195000 ;
        RECT  1.485000 190.395000  1.685000 190.595000 ;
        RECT  1.485000 190.795000  1.685000 190.995000 ;
        RECT  1.485000 191.195000  1.685000 191.395000 ;
        RECT  1.485000 191.595000  1.685000 191.795000 ;
        RECT  1.485000 191.995000  1.685000 192.195000 ;
        RECT  1.485000 192.395000  1.685000 192.595000 ;
        RECT  1.485000 192.795000  1.685000 192.995000 ;
        RECT  1.485000 193.195000  1.685000 193.395000 ;
        RECT  1.485000 193.595000  1.685000 193.795000 ;
        RECT  1.485000 193.995000  1.685000 194.195000 ;
        RECT  1.485000 194.395000  1.685000 194.595000 ;
        RECT  1.485000 194.795000  1.685000 194.995000 ;
        RECT  1.485000 195.200000  1.685000 195.400000 ;
        RECT  1.485000 195.605000  1.685000 195.805000 ;
        RECT  1.485000 196.010000  1.685000 196.210000 ;
        RECT  1.485000 196.415000  1.685000 196.615000 ;
        RECT  1.485000 196.820000  1.685000 197.020000 ;
        RECT  1.485000 197.225000  1.685000 197.425000 ;
        RECT  1.485000 197.630000  1.685000 197.830000 ;
        RECT  1.485000 198.035000  1.685000 198.235000 ;
        RECT  1.485000 198.440000  1.685000 198.640000 ;
        RECT  1.485000 198.845000  1.685000 199.045000 ;
        RECT  1.485000 199.250000  1.685000 199.450000 ;
        RECT  1.485000 199.655000  1.685000 199.855000 ;
        RECT  1.815000  25.910000  2.015000  26.110000 ;
        RECT  1.815000  26.340000  2.015000  26.540000 ;
        RECT  1.815000  26.770000  2.015000  26.970000 ;
        RECT  1.815000  27.200000  2.015000  27.400000 ;
        RECT  1.815000  27.630000  2.015000  27.830000 ;
        RECT  1.815000  28.060000  2.015000  28.260000 ;
        RECT  1.815000  28.490000  2.015000  28.690000 ;
        RECT  1.815000  28.920000  2.015000  29.120000 ;
        RECT  1.815000  29.350000  2.015000  29.550000 ;
        RECT  1.815000  29.780000  2.015000  29.980000 ;
        RECT  1.815000  30.210000  2.015000  30.410000 ;
        RECT  1.885000 175.995000  2.085000 176.195000 ;
        RECT  1.885000 176.395000  2.085000 176.595000 ;
        RECT  1.885000 176.795000  2.085000 176.995000 ;
        RECT  1.885000 177.195000  2.085000 177.395000 ;
        RECT  1.885000 177.595000  2.085000 177.795000 ;
        RECT  1.885000 177.995000  2.085000 178.195000 ;
        RECT  1.885000 178.395000  2.085000 178.595000 ;
        RECT  1.885000 178.795000  2.085000 178.995000 ;
        RECT  1.885000 179.195000  2.085000 179.395000 ;
        RECT  1.885000 179.595000  2.085000 179.795000 ;
        RECT  1.885000 179.995000  2.085000 180.195000 ;
        RECT  1.885000 180.395000  2.085000 180.595000 ;
        RECT  1.885000 180.795000  2.085000 180.995000 ;
        RECT  1.885000 181.195000  2.085000 181.395000 ;
        RECT  1.885000 181.595000  2.085000 181.795000 ;
        RECT  1.885000 181.995000  2.085000 182.195000 ;
        RECT  1.885000 182.395000  2.085000 182.595000 ;
        RECT  1.885000 182.795000  2.085000 182.995000 ;
        RECT  1.885000 183.195000  2.085000 183.395000 ;
        RECT  1.885000 183.595000  2.085000 183.795000 ;
        RECT  1.885000 183.995000  2.085000 184.195000 ;
        RECT  1.885000 184.395000  2.085000 184.595000 ;
        RECT  1.885000 184.795000  2.085000 184.995000 ;
        RECT  1.885000 185.195000  2.085000 185.395000 ;
        RECT  1.885000 185.595000  2.085000 185.795000 ;
        RECT  1.885000 185.995000  2.085000 186.195000 ;
        RECT  1.885000 186.395000  2.085000 186.595000 ;
        RECT  1.885000 186.795000  2.085000 186.995000 ;
        RECT  1.885000 187.195000  2.085000 187.395000 ;
        RECT  1.885000 187.595000  2.085000 187.795000 ;
        RECT  1.885000 187.995000  2.085000 188.195000 ;
        RECT  1.885000 188.395000  2.085000 188.595000 ;
        RECT  1.885000 188.795000  2.085000 188.995000 ;
        RECT  1.885000 189.195000  2.085000 189.395000 ;
        RECT  1.885000 189.595000  2.085000 189.795000 ;
        RECT  1.885000 189.995000  2.085000 190.195000 ;
        RECT  1.885000 190.395000  2.085000 190.595000 ;
        RECT  1.885000 190.795000  2.085000 190.995000 ;
        RECT  1.885000 191.195000  2.085000 191.395000 ;
        RECT  1.885000 191.595000  2.085000 191.795000 ;
        RECT  1.885000 191.995000  2.085000 192.195000 ;
        RECT  1.885000 192.395000  2.085000 192.595000 ;
        RECT  1.885000 192.795000  2.085000 192.995000 ;
        RECT  1.885000 193.195000  2.085000 193.395000 ;
        RECT  1.885000 193.595000  2.085000 193.795000 ;
        RECT  1.885000 193.995000  2.085000 194.195000 ;
        RECT  1.885000 194.395000  2.085000 194.595000 ;
        RECT  1.885000 194.795000  2.085000 194.995000 ;
        RECT  1.885000 195.200000  2.085000 195.400000 ;
        RECT  1.885000 195.605000  2.085000 195.805000 ;
        RECT  1.885000 196.010000  2.085000 196.210000 ;
        RECT  1.885000 196.415000  2.085000 196.615000 ;
        RECT  1.885000 196.820000  2.085000 197.020000 ;
        RECT  1.885000 197.225000  2.085000 197.425000 ;
        RECT  1.885000 197.630000  2.085000 197.830000 ;
        RECT  1.885000 198.035000  2.085000 198.235000 ;
        RECT  1.885000 198.440000  2.085000 198.640000 ;
        RECT  1.885000 198.845000  2.085000 199.045000 ;
        RECT  1.885000 199.250000  2.085000 199.450000 ;
        RECT  1.885000 199.655000  2.085000 199.855000 ;
        RECT  2.225000  25.910000  2.425000  26.110000 ;
        RECT  2.225000  26.340000  2.425000  26.540000 ;
        RECT  2.225000  26.770000  2.425000  26.970000 ;
        RECT  2.225000  27.200000  2.425000  27.400000 ;
        RECT  2.225000  27.630000  2.425000  27.830000 ;
        RECT  2.225000  28.060000  2.425000  28.260000 ;
        RECT  2.225000  28.490000  2.425000  28.690000 ;
        RECT  2.225000  28.920000  2.425000  29.120000 ;
        RECT  2.225000  29.350000  2.425000  29.550000 ;
        RECT  2.225000  29.780000  2.425000  29.980000 ;
        RECT  2.225000  30.210000  2.425000  30.410000 ;
        RECT  2.285000 175.995000  2.485000 176.195000 ;
        RECT  2.285000 176.395000  2.485000 176.595000 ;
        RECT  2.285000 176.795000  2.485000 176.995000 ;
        RECT  2.285000 177.195000  2.485000 177.395000 ;
        RECT  2.285000 177.595000  2.485000 177.795000 ;
        RECT  2.285000 177.995000  2.485000 178.195000 ;
        RECT  2.285000 178.395000  2.485000 178.595000 ;
        RECT  2.285000 178.795000  2.485000 178.995000 ;
        RECT  2.285000 179.195000  2.485000 179.395000 ;
        RECT  2.285000 179.595000  2.485000 179.795000 ;
        RECT  2.285000 179.995000  2.485000 180.195000 ;
        RECT  2.285000 180.395000  2.485000 180.595000 ;
        RECT  2.285000 180.795000  2.485000 180.995000 ;
        RECT  2.285000 181.195000  2.485000 181.395000 ;
        RECT  2.285000 181.595000  2.485000 181.795000 ;
        RECT  2.285000 181.995000  2.485000 182.195000 ;
        RECT  2.285000 182.395000  2.485000 182.595000 ;
        RECT  2.285000 182.795000  2.485000 182.995000 ;
        RECT  2.285000 183.195000  2.485000 183.395000 ;
        RECT  2.285000 183.595000  2.485000 183.795000 ;
        RECT  2.285000 183.995000  2.485000 184.195000 ;
        RECT  2.285000 184.395000  2.485000 184.595000 ;
        RECT  2.285000 184.795000  2.485000 184.995000 ;
        RECT  2.285000 185.195000  2.485000 185.395000 ;
        RECT  2.285000 185.595000  2.485000 185.795000 ;
        RECT  2.285000 185.995000  2.485000 186.195000 ;
        RECT  2.285000 186.395000  2.485000 186.595000 ;
        RECT  2.285000 186.795000  2.485000 186.995000 ;
        RECT  2.285000 187.195000  2.485000 187.395000 ;
        RECT  2.285000 187.595000  2.485000 187.795000 ;
        RECT  2.285000 187.995000  2.485000 188.195000 ;
        RECT  2.285000 188.395000  2.485000 188.595000 ;
        RECT  2.285000 188.795000  2.485000 188.995000 ;
        RECT  2.285000 189.195000  2.485000 189.395000 ;
        RECT  2.285000 189.595000  2.485000 189.795000 ;
        RECT  2.285000 189.995000  2.485000 190.195000 ;
        RECT  2.285000 190.395000  2.485000 190.595000 ;
        RECT  2.285000 190.795000  2.485000 190.995000 ;
        RECT  2.285000 191.195000  2.485000 191.395000 ;
        RECT  2.285000 191.595000  2.485000 191.795000 ;
        RECT  2.285000 191.995000  2.485000 192.195000 ;
        RECT  2.285000 192.395000  2.485000 192.595000 ;
        RECT  2.285000 192.795000  2.485000 192.995000 ;
        RECT  2.285000 193.195000  2.485000 193.395000 ;
        RECT  2.285000 193.595000  2.485000 193.795000 ;
        RECT  2.285000 193.995000  2.485000 194.195000 ;
        RECT  2.285000 194.395000  2.485000 194.595000 ;
        RECT  2.285000 194.795000  2.485000 194.995000 ;
        RECT  2.285000 195.200000  2.485000 195.400000 ;
        RECT  2.285000 195.605000  2.485000 195.805000 ;
        RECT  2.285000 196.010000  2.485000 196.210000 ;
        RECT  2.285000 196.415000  2.485000 196.615000 ;
        RECT  2.285000 196.820000  2.485000 197.020000 ;
        RECT  2.285000 197.225000  2.485000 197.425000 ;
        RECT  2.285000 197.630000  2.485000 197.830000 ;
        RECT  2.285000 198.035000  2.485000 198.235000 ;
        RECT  2.285000 198.440000  2.485000 198.640000 ;
        RECT  2.285000 198.845000  2.485000 199.045000 ;
        RECT  2.285000 199.250000  2.485000 199.450000 ;
        RECT  2.285000 199.655000  2.485000 199.855000 ;
        RECT  2.635000  25.910000  2.835000  26.110000 ;
        RECT  2.635000  26.340000  2.835000  26.540000 ;
        RECT  2.635000  26.770000  2.835000  26.970000 ;
        RECT  2.635000  27.200000  2.835000  27.400000 ;
        RECT  2.635000  27.630000  2.835000  27.830000 ;
        RECT  2.635000  28.060000  2.835000  28.260000 ;
        RECT  2.635000  28.490000  2.835000  28.690000 ;
        RECT  2.635000  28.920000  2.835000  29.120000 ;
        RECT  2.635000  29.350000  2.835000  29.550000 ;
        RECT  2.635000  29.780000  2.835000  29.980000 ;
        RECT  2.635000  30.210000  2.835000  30.410000 ;
        RECT  2.685000 175.995000  2.885000 176.195000 ;
        RECT  2.685000 176.395000  2.885000 176.595000 ;
        RECT  2.685000 176.795000  2.885000 176.995000 ;
        RECT  2.685000 177.195000  2.885000 177.395000 ;
        RECT  2.685000 177.595000  2.885000 177.795000 ;
        RECT  2.685000 177.995000  2.885000 178.195000 ;
        RECT  2.685000 178.395000  2.885000 178.595000 ;
        RECT  2.685000 178.795000  2.885000 178.995000 ;
        RECT  2.685000 179.195000  2.885000 179.395000 ;
        RECT  2.685000 179.595000  2.885000 179.795000 ;
        RECT  2.685000 179.995000  2.885000 180.195000 ;
        RECT  2.685000 180.395000  2.885000 180.595000 ;
        RECT  2.685000 180.795000  2.885000 180.995000 ;
        RECT  2.685000 181.195000  2.885000 181.395000 ;
        RECT  2.685000 181.595000  2.885000 181.795000 ;
        RECT  2.685000 181.995000  2.885000 182.195000 ;
        RECT  2.685000 182.395000  2.885000 182.595000 ;
        RECT  2.685000 182.795000  2.885000 182.995000 ;
        RECT  2.685000 183.195000  2.885000 183.395000 ;
        RECT  2.685000 183.595000  2.885000 183.795000 ;
        RECT  2.685000 183.995000  2.885000 184.195000 ;
        RECT  2.685000 184.395000  2.885000 184.595000 ;
        RECT  2.685000 184.795000  2.885000 184.995000 ;
        RECT  2.685000 185.195000  2.885000 185.395000 ;
        RECT  2.685000 185.595000  2.885000 185.795000 ;
        RECT  2.685000 185.995000  2.885000 186.195000 ;
        RECT  2.685000 186.395000  2.885000 186.595000 ;
        RECT  2.685000 186.795000  2.885000 186.995000 ;
        RECT  2.685000 187.195000  2.885000 187.395000 ;
        RECT  2.685000 187.595000  2.885000 187.795000 ;
        RECT  2.685000 187.995000  2.885000 188.195000 ;
        RECT  2.685000 188.395000  2.885000 188.595000 ;
        RECT  2.685000 188.795000  2.885000 188.995000 ;
        RECT  2.685000 189.195000  2.885000 189.395000 ;
        RECT  2.685000 189.595000  2.885000 189.795000 ;
        RECT  2.685000 189.995000  2.885000 190.195000 ;
        RECT  2.685000 190.395000  2.885000 190.595000 ;
        RECT  2.685000 190.795000  2.885000 190.995000 ;
        RECT  2.685000 191.195000  2.885000 191.395000 ;
        RECT  2.685000 191.595000  2.885000 191.795000 ;
        RECT  2.685000 191.995000  2.885000 192.195000 ;
        RECT  2.685000 192.395000  2.885000 192.595000 ;
        RECT  2.685000 192.795000  2.885000 192.995000 ;
        RECT  2.685000 193.195000  2.885000 193.395000 ;
        RECT  2.685000 193.595000  2.885000 193.795000 ;
        RECT  2.685000 193.995000  2.885000 194.195000 ;
        RECT  2.685000 194.395000  2.885000 194.595000 ;
        RECT  2.685000 194.795000  2.885000 194.995000 ;
        RECT  2.685000 195.200000  2.885000 195.400000 ;
        RECT  2.685000 195.605000  2.885000 195.805000 ;
        RECT  2.685000 196.010000  2.885000 196.210000 ;
        RECT  2.685000 196.415000  2.885000 196.615000 ;
        RECT  2.685000 196.820000  2.885000 197.020000 ;
        RECT  2.685000 197.225000  2.885000 197.425000 ;
        RECT  2.685000 197.630000  2.885000 197.830000 ;
        RECT  2.685000 198.035000  2.885000 198.235000 ;
        RECT  2.685000 198.440000  2.885000 198.640000 ;
        RECT  2.685000 198.845000  2.885000 199.045000 ;
        RECT  2.685000 199.250000  2.885000 199.450000 ;
        RECT  2.685000 199.655000  2.885000 199.855000 ;
        RECT  3.045000  25.910000  3.245000  26.110000 ;
        RECT  3.045000  26.340000  3.245000  26.540000 ;
        RECT  3.045000  26.770000  3.245000  26.970000 ;
        RECT  3.045000  27.200000  3.245000  27.400000 ;
        RECT  3.045000  27.630000  3.245000  27.830000 ;
        RECT  3.045000  28.060000  3.245000  28.260000 ;
        RECT  3.045000  28.490000  3.245000  28.690000 ;
        RECT  3.045000  28.920000  3.245000  29.120000 ;
        RECT  3.045000  29.350000  3.245000  29.550000 ;
        RECT  3.045000  29.780000  3.245000  29.980000 ;
        RECT  3.045000  30.210000  3.245000  30.410000 ;
        RECT  3.085000 175.995000  3.285000 176.195000 ;
        RECT  3.085000 176.395000  3.285000 176.595000 ;
        RECT  3.085000 176.795000  3.285000 176.995000 ;
        RECT  3.085000 177.195000  3.285000 177.395000 ;
        RECT  3.085000 177.595000  3.285000 177.795000 ;
        RECT  3.085000 177.995000  3.285000 178.195000 ;
        RECT  3.085000 178.395000  3.285000 178.595000 ;
        RECT  3.085000 178.795000  3.285000 178.995000 ;
        RECT  3.085000 179.195000  3.285000 179.395000 ;
        RECT  3.085000 179.595000  3.285000 179.795000 ;
        RECT  3.085000 179.995000  3.285000 180.195000 ;
        RECT  3.085000 180.395000  3.285000 180.595000 ;
        RECT  3.085000 180.795000  3.285000 180.995000 ;
        RECT  3.085000 181.195000  3.285000 181.395000 ;
        RECT  3.085000 181.595000  3.285000 181.795000 ;
        RECT  3.085000 181.995000  3.285000 182.195000 ;
        RECT  3.085000 182.395000  3.285000 182.595000 ;
        RECT  3.085000 182.795000  3.285000 182.995000 ;
        RECT  3.085000 183.195000  3.285000 183.395000 ;
        RECT  3.085000 183.595000  3.285000 183.795000 ;
        RECT  3.085000 183.995000  3.285000 184.195000 ;
        RECT  3.085000 184.395000  3.285000 184.595000 ;
        RECT  3.085000 184.795000  3.285000 184.995000 ;
        RECT  3.085000 185.195000  3.285000 185.395000 ;
        RECT  3.085000 185.595000  3.285000 185.795000 ;
        RECT  3.085000 185.995000  3.285000 186.195000 ;
        RECT  3.085000 186.395000  3.285000 186.595000 ;
        RECT  3.085000 186.795000  3.285000 186.995000 ;
        RECT  3.085000 187.195000  3.285000 187.395000 ;
        RECT  3.085000 187.595000  3.285000 187.795000 ;
        RECT  3.085000 187.995000  3.285000 188.195000 ;
        RECT  3.085000 188.395000  3.285000 188.595000 ;
        RECT  3.085000 188.795000  3.285000 188.995000 ;
        RECT  3.085000 189.195000  3.285000 189.395000 ;
        RECT  3.085000 189.595000  3.285000 189.795000 ;
        RECT  3.085000 189.995000  3.285000 190.195000 ;
        RECT  3.085000 190.395000  3.285000 190.595000 ;
        RECT  3.085000 190.795000  3.285000 190.995000 ;
        RECT  3.085000 191.195000  3.285000 191.395000 ;
        RECT  3.085000 191.595000  3.285000 191.795000 ;
        RECT  3.085000 191.995000  3.285000 192.195000 ;
        RECT  3.085000 192.395000  3.285000 192.595000 ;
        RECT  3.085000 192.795000  3.285000 192.995000 ;
        RECT  3.085000 193.195000  3.285000 193.395000 ;
        RECT  3.085000 193.595000  3.285000 193.795000 ;
        RECT  3.085000 193.995000  3.285000 194.195000 ;
        RECT  3.085000 194.395000  3.285000 194.595000 ;
        RECT  3.085000 194.795000  3.285000 194.995000 ;
        RECT  3.085000 195.200000  3.285000 195.400000 ;
        RECT  3.085000 195.605000  3.285000 195.805000 ;
        RECT  3.085000 196.010000  3.285000 196.210000 ;
        RECT  3.085000 196.415000  3.285000 196.615000 ;
        RECT  3.085000 196.820000  3.285000 197.020000 ;
        RECT  3.085000 197.225000  3.285000 197.425000 ;
        RECT  3.085000 197.630000  3.285000 197.830000 ;
        RECT  3.085000 198.035000  3.285000 198.235000 ;
        RECT  3.085000 198.440000  3.285000 198.640000 ;
        RECT  3.085000 198.845000  3.285000 199.045000 ;
        RECT  3.085000 199.250000  3.285000 199.450000 ;
        RECT  3.085000 199.655000  3.285000 199.855000 ;
        RECT  3.450000  25.910000  3.650000  26.110000 ;
        RECT  3.450000  26.340000  3.650000  26.540000 ;
        RECT  3.450000  26.770000  3.650000  26.970000 ;
        RECT  3.450000  27.200000  3.650000  27.400000 ;
        RECT  3.450000  27.630000  3.650000  27.830000 ;
        RECT  3.450000  28.060000  3.650000  28.260000 ;
        RECT  3.450000  28.490000  3.650000  28.690000 ;
        RECT  3.450000  28.920000  3.650000  29.120000 ;
        RECT  3.450000  29.350000  3.650000  29.550000 ;
        RECT  3.450000  29.780000  3.650000  29.980000 ;
        RECT  3.450000  30.210000  3.650000  30.410000 ;
        RECT  3.485000 175.995000  3.685000 176.195000 ;
        RECT  3.485000 176.395000  3.685000 176.595000 ;
        RECT  3.485000 176.795000  3.685000 176.995000 ;
        RECT  3.485000 177.195000  3.685000 177.395000 ;
        RECT  3.485000 177.595000  3.685000 177.795000 ;
        RECT  3.485000 177.995000  3.685000 178.195000 ;
        RECT  3.485000 178.395000  3.685000 178.595000 ;
        RECT  3.485000 178.795000  3.685000 178.995000 ;
        RECT  3.485000 179.195000  3.685000 179.395000 ;
        RECT  3.485000 179.595000  3.685000 179.795000 ;
        RECT  3.485000 179.995000  3.685000 180.195000 ;
        RECT  3.485000 180.395000  3.685000 180.595000 ;
        RECT  3.485000 180.795000  3.685000 180.995000 ;
        RECT  3.485000 181.195000  3.685000 181.395000 ;
        RECT  3.485000 181.595000  3.685000 181.795000 ;
        RECT  3.485000 181.995000  3.685000 182.195000 ;
        RECT  3.485000 182.395000  3.685000 182.595000 ;
        RECT  3.485000 182.795000  3.685000 182.995000 ;
        RECT  3.485000 183.195000  3.685000 183.395000 ;
        RECT  3.485000 183.595000  3.685000 183.795000 ;
        RECT  3.485000 183.995000  3.685000 184.195000 ;
        RECT  3.485000 184.395000  3.685000 184.595000 ;
        RECT  3.485000 184.795000  3.685000 184.995000 ;
        RECT  3.485000 185.195000  3.685000 185.395000 ;
        RECT  3.485000 185.595000  3.685000 185.795000 ;
        RECT  3.485000 185.995000  3.685000 186.195000 ;
        RECT  3.485000 186.395000  3.685000 186.595000 ;
        RECT  3.485000 186.795000  3.685000 186.995000 ;
        RECT  3.485000 187.195000  3.685000 187.395000 ;
        RECT  3.485000 187.595000  3.685000 187.795000 ;
        RECT  3.485000 187.995000  3.685000 188.195000 ;
        RECT  3.485000 188.395000  3.685000 188.595000 ;
        RECT  3.485000 188.795000  3.685000 188.995000 ;
        RECT  3.485000 189.195000  3.685000 189.395000 ;
        RECT  3.485000 189.595000  3.685000 189.795000 ;
        RECT  3.485000 189.995000  3.685000 190.195000 ;
        RECT  3.485000 190.395000  3.685000 190.595000 ;
        RECT  3.485000 190.795000  3.685000 190.995000 ;
        RECT  3.485000 191.195000  3.685000 191.395000 ;
        RECT  3.485000 191.595000  3.685000 191.795000 ;
        RECT  3.485000 191.995000  3.685000 192.195000 ;
        RECT  3.485000 192.395000  3.685000 192.595000 ;
        RECT  3.485000 192.795000  3.685000 192.995000 ;
        RECT  3.485000 193.195000  3.685000 193.395000 ;
        RECT  3.485000 193.595000  3.685000 193.795000 ;
        RECT  3.485000 193.995000  3.685000 194.195000 ;
        RECT  3.485000 194.395000  3.685000 194.595000 ;
        RECT  3.485000 194.795000  3.685000 194.995000 ;
        RECT  3.485000 195.200000  3.685000 195.400000 ;
        RECT  3.485000 195.605000  3.685000 195.805000 ;
        RECT  3.485000 196.010000  3.685000 196.210000 ;
        RECT  3.485000 196.415000  3.685000 196.615000 ;
        RECT  3.485000 196.820000  3.685000 197.020000 ;
        RECT  3.485000 197.225000  3.685000 197.425000 ;
        RECT  3.485000 197.630000  3.685000 197.830000 ;
        RECT  3.485000 198.035000  3.685000 198.235000 ;
        RECT  3.485000 198.440000  3.685000 198.640000 ;
        RECT  3.485000 198.845000  3.685000 199.045000 ;
        RECT  3.485000 199.250000  3.685000 199.450000 ;
        RECT  3.485000 199.655000  3.685000 199.855000 ;
        RECT  3.855000  25.910000  4.055000  26.110000 ;
        RECT  3.855000  26.340000  4.055000  26.540000 ;
        RECT  3.855000  26.770000  4.055000  26.970000 ;
        RECT  3.855000  27.200000  4.055000  27.400000 ;
        RECT  3.855000  27.630000  4.055000  27.830000 ;
        RECT  3.855000  28.060000  4.055000  28.260000 ;
        RECT  3.855000  28.490000  4.055000  28.690000 ;
        RECT  3.855000  28.920000  4.055000  29.120000 ;
        RECT  3.855000  29.350000  4.055000  29.550000 ;
        RECT  3.855000  29.780000  4.055000  29.980000 ;
        RECT  3.855000  30.210000  4.055000  30.410000 ;
        RECT  3.885000 175.995000  4.085000 176.195000 ;
        RECT  3.885000 176.395000  4.085000 176.595000 ;
        RECT  3.885000 176.795000  4.085000 176.995000 ;
        RECT  3.885000 177.195000  4.085000 177.395000 ;
        RECT  3.885000 177.595000  4.085000 177.795000 ;
        RECT  3.885000 177.995000  4.085000 178.195000 ;
        RECT  3.885000 178.395000  4.085000 178.595000 ;
        RECT  3.885000 178.795000  4.085000 178.995000 ;
        RECT  3.885000 179.195000  4.085000 179.395000 ;
        RECT  3.885000 179.595000  4.085000 179.795000 ;
        RECT  3.885000 179.995000  4.085000 180.195000 ;
        RECT  3.885000 180.395000  4.085000 180.595000 ;
        RECT  3.885000 180.795000  4.085000 180.995000 ;
        RECT  3.885000 181.195000  4.085000 181.395000 ;
        RECT  3.885000 181.595000  4.085000 181.795000 ;
        RECT  3.885000 181.995000  4.085000 182.195000 ;
        RECT  3.885000 182.395000  4.085000 182.595000 ;
        RECT  3.885000 182.795000  4.085000 182.995000 ;
        RECT  3.885000 183.195000  4.085000 183.395000 ;
        RECT  3.885000 183.595000  4.085000 183.795000 ;
        RECT  3.885000 183.995000  4.085000 184.195000 ;
        RECT  3.885000 184.395000  4.085000 184.595000 ;
        RECT  3.885000 184.795000  4.085000 184.995000 ;
        RECT  3.885000 185.195000  4.085000 185.395000 ;
        RECT  3.885000 185.595000  4.085000 185.795000 ;
        RECT  3.885000 185.995000  4.085000 186.195000 ;
        RECT  3.885000 186.395000  4.085000 186.595000 ;
        RECT  3.885000 186.795000  4.085000 186.995000 ;
        RECT  3.885000 187.195000  4.085000 187.395000 ;
        RECT  3.885000 187.595000  4.085000 187.795000 ;
        RECT  3.885000 187.995000  4.085000 188.195000 ;
        RECT  3.885000 188.395000  4.085000 188.595000 ;
        RECT  3.885000 188.795000  4.085000 188.995000 ;
        RECT  3.885000 189.195000  4.085000 189.395000 ;
        RECT  3.885000 189.595000  4.085000 189.795000 ;
        RECT  3.885000 189.995000  4.085000 190.195000 ;
        RECT  3.885000 190.395000  4.085000 190.595000 ;
        RECT  3.885000 190.795000  4.085000 190.995000 ;
        RECT  3.885000 191.195000  4.085000 191.395000 ;
        RECT  3.885000 191.595000  4.085000 191.795000 ;
        RECT  3.885000 191.995000  4.085000 192.195000 ;
        RECT  3.885000 192.395000  4.085000 192.595000 ;
        RECT  3.885000 192.795000  4.085000 192.995000 ;
        RECT  3.885000 193.195000  4.085000 193.395000 ;
        RECT  3.885000 193.595000  4.085000 193.795000 ;
        RECT  3.885000 193.995000  4.085000 194.195000 ;
        RECT  3.885000 194.395000  4.085000 194.595000 ;
        RECT  3.885000 194.795000  4.085000 194.995000 ;
        RECT  3.885000 195.200000  4.085000 195.400000 ;
        RECT  3.885000 195.605000  4.085000 195.805000 ;
        RECT  3.885000 196.010000  4.085000 196.210000 ;
        RECT  3.885000 196.415000  4.085000 196.615000 ;
        RECT  3.885000 196.820000  4.085000 197.020000 ;
        RECT  3.885000 197.225000  4.085000 197.425000 ;
        RECT  3.885000 197.630000  4.085000 197.830000 ;
        RECT  3.885000 198.035000  4.085000 198.235000 ;
        RECT  3.885000 198.440000  4.085000 198.640000 ;
        RECT  3.885000 198.845000  4.085000 199.045000 ;
        RECT  3.885000 199.250000  4.085000 199.450000 ;
        RECT  3.885000 199.655000  4.085000 199.855000 ;
        RECT  4.260000  25.910000  4.460000  26.110000 ;
        RECT  4.260000  26.340000  4.460000  26.540000 ;
        RECT  4.260000  26.770000  4.460000  26.970000 ;
        RECT  4.260000  27.200000  4.460000  27.400000 ;
        RECT  4.260000  27.630000  4.460000  27.830000 ;
        RECT  4.260000  28.060000  4.460000  28.260000 ;
        RECT  4.260000  28.490000  4.460000  28.690000 ;
        RECT  4.260000  28.920000  4.460000  29.120000 ;
        RECT  4.260000  29.350000  4.460000  29.550000 ;
        RECT  4.260000  29.780000  4.460000  29.980000 ;
        RECT  4.260000  30.210000  4.460000  30.410000 ;
        RECT  4.285000 175.995000  4.485000 176.195000 ;
        RECT  4.285000 176.395000  4.485000 176.595000 ;
        RECT  4.285000 176.795000  4.485000 176.995000 ;
        RECT  4.285000 177.195000  4.485000 177.395000 ;
        RECT  4.285000 177.595000  4.485000 177.795000 ;
        RECT  4.285000 177.995000  4.485000 178.195000 ;
        RECT  4.285000 178.395000  4.485000 178.595000 ;
        RECT  4.285000 178.795000  4.485000 178.995000 ;
        RECT  4.285000 179.195000  4.485000 179.395000 ;
        RECT  4.285000 179.595000  4.485000 179.795000 ;
        RECT  4.285000 179.995000  4.485000 180.195000 ;
        RECT  4.285000 180.395000  4.485000 180.595000 ;
        RECT  4.285000 180.795000  4.485000 180.995000 ;
        RECT  4.285000 181.195000  4.485000 181.395000 ;
        RECT  4.285000 181.595000  4.485000 181.795000 ;
        RECT  4.285000 181.995000  4.485000 182.195000 ;
        RECT  4.285000 182.395000  4.485000 182.595000 ;
        RECT  4.285000 182.795000  4.485000 182.995000 ;
        RECT  4.285000 183.195000  4.485000 183.395000 ;
        RECT  4.285000 183.595000  4.485000 183.795000 ;
        RECT  4.285000 183.995000  4.485000 184.195000 ;
        RECT  4.285000 184.395000  4.485000 184.595000 ;
        RECT  4.285000 184.795000  4.485000 184.995000 ;
        RECT  4.285000 185.195000  4.485000 185.395000 ;
        RECT  4.285000 185.595000  4.485000 185.795000 ;
        RECT  4.285000 185.995000  4.485000 186.195000 ;
        RECT  4.285000 186.395000  4.485000 186.595000 ;
        RECT  4.285000 186.795000  4.485000 186.995000 ;
        RECT  4.285000 187.195000  4.485000 187.395000 ;
        RECT  4.285000 187.595000  4.485000 187.795000 ;
        RECT  4.285000 187.995000  4.485000 188.195000 ;
        RECT  4.285000 188.395000  4.485000 188.595000 ;
        RECT  4.285000 188.795000  4.485000 188.995000 ;
        RECT  4.285000 189.195000  4.485000 189.395000 ;
        RECT  4.285000 189.595000  4.485000 189.795000 ;
        RECT  4.285000 189.995000  4.485000 190.195000 ;
        RECT  4.285000 190.395000  4.485000 190.595000 ;
        RECT  4.285000 190.795000  4.485000 190.995000 ;
        RECT  4.285000 191.195000  4.485000 191.395000 ;
        RECT  4.285000 191.595000  4.485000 191.795000 ;
        RECT  4.285000 191.995000  4.485000 192.195000 ;
        RECT  4.285000 192.395000  4.485000 192.595000 ;
        RECT  4.285000 192.795000  4.485000 192.995000 ;
        RECT  4.285000 193.195000  4.485000 193.395000 ;
        RECT  4.285000 193.595000  4.485000 193.795000 ;
        RECT  4.285000 193.995000  4.485000 194.195000 ;
        RECT  4.285000 194.395000  4.485000 194.595000 ;
        RECT  4.285000 194.795000  4.485000 194.995000 ;
        RECT  4.285000 195.200000  4.485000 195.400000 ;
        RECT  4.285000 195.605000  4.485000 195.805000 ;
        RECT  4.285000 196.010000  4.485000 196.210000 ;
        RECT  4.285000 196.415000  4.485000 196.615000 ;
        RECT  4.285000 196.820000  4.485000 197.020000 ;
        RECT  4.285000 197.225000  4.485000 197.425000 ;
        RECT  4.285000 197.630000  4.485000 197.830000 ;
        RECT  4.285000 198.035000  4.485000 198.235000 ;
        RECT  4.285000 198.440000  4.485000 198.640000 ;
        RECT  4.285000 198.845000  4.485000 199.045000 ;
        RECT  4.285000 199.250000  4.485000 199.450000 ;
        RECT  4.285000 199.655000  4.485000 199.855000 ;
        RECT  4.665000  25.910000  4.865000  26.110000 ;
        RECT  4.665000  26.340000  4.865000  26.540000 ;
        RECT  4.665000  26.770000  4.865000  26.970000 ;
        RECT  4.665000  27.200000  4.865000  27.400000 ;
        RECT  4.665000  27.630000  4.865000  27.830000 ;
        RECT  4.665000  28.060000  4.865000  28.260000 ;
        RECT  4.665000  28.490000  4.865000  28.690000 ;
        RECT  4.665000  28.920000  4.865000  29.120000 ;
        RECT  4.665000  29.350000  4.865000  29.550000 ;
        RECT  4.665000  29.780000  4.865000  29.980000 ;
        RECT  4.665000  30.210000  4.865000  30.410000 ;
        RECT  4.685000 175.995000  4.885000 176.195000 ;
        RECT  4.685000 176.395000  4.885000 176.595000 ;
        RECT  4.685000 176.795000  4.885000 176.995000 ;
        RECT  4.685000 177.195000  4.885000 177.395000 ;
        RECT  4.685000 177.595000  4.885000 177.795000 ;
        RECT  4.685000 177.995000  4.885000 178.195000 ;
        RECT  4.685000 178.395000  4.885000 178.595000 ;
        RECT  4.685000 178.795000  4.885000 178.995000 ;
        RECT  4.685000 179.195000  4.885000 179.395000 ;
        RECT  4.685000 179.595000  4.885000 179.795000 ;
        RECT  4.685000 179.995000  4.885000 180.195000 ;
        RECT  4.685000 180.395000  4.885000 180.595000 ;
        RECT  4.685000 180.795000  4.885000 180.995000 ;
        RECT  4.685000 181.195000  4.885000 181.395000 ;
        RECT  4.685000 181.595000  4.885000 181.795000 ;
        RECT  4.685000 181.995000  4.885000 182.195000 ;
        RECT  4.685000 182.395000  4.885000 182.595000 ;
        RECT  4.685000 182.795000  4.885000 182.995000 ;
        RECT  4.685000 183.195000  4.885000 183.395000 ;
        RECT  4.685000 183.595000  4.885000 183.795000 ;
        RECT  4.685000 183.995000  4.885000 184.195000 ;
        RECT  4.685000 184.395000  4.885000 184.595000 ;
        RECT  4.685000 184.795000  4.885000 184.995000 ;
        RECT  4.685000 185.195000  4.885000 185.395000 ;
        RECT  4.685000 185.595000  4.885000 185.795000 ;
        RECT  4.685000 185.995000  4.885000 186.195000 ;
        RECT  4.685000 186.395000  4.885000 186.595000 ;
        RECT  4.685000 186.795000  4.885000 186.995000 ;
        RECT  4.685000 187.195000  4.885000 187.395000 ;
        RECT  4.685000 187.595000  4.885000 187.795000 ;
        RECT  4.685000 187.995000  4.885000 188.195000 ;
        RECT  4.685000 188.395000  4.885000 188.595000 ;
        RECT  4.685000 188.795000  4.885000 188.995000 ;
        RECT  4.685000 189.195000  4.885000 189.395000 ;
        RECT  4.685000 189.595000  4.885000 189.795000 ;
        RECT  4.685000 189.995000  4.885000 190.195000 ;
        RECT  4.685000 190.395000  4.885000 190.595000 ;
        RECT  4.685000 190.795000  4.885000 190.995000 ;
        RECT  4.685000 191.195000  4.885000 191.395000 ;
        RECT  4.685000 191.595000  4.885000 191.795000 ;
        RECT  4.685000 191.995000  4.885000 192.195000 ;
        RECT  4.685000 192.395000  4.885000 192.595000 ;
        RECT  4.685000 192.795000  4.885000 192.995000 ;
        RECT  4.685000 193.195000  4.885000 193.395000 ;
        RECT  4.685000 193.595000  4.885000 193.795000 ;
        RECT  4.685000 193.995000  4.885000 194.195000 ;
        RECT  4.685000 194.395000  4.885000 194.595000 ;
        RECT  4.685000 194.795000  4.885000 194.995000 ;
        RECT  4.685000 195.200000  4.885000 195.400000 ;
        RECT  4.685000 195.605000  4.885000 195.805000 ;
        RECT  4.685000 196.010000  4.885000 196.210000 ;
        RECT  4.685000 196.415000  4.885000 196.615000 ;
        RECT  4.685000 196.820000  4.885000 197.020000 ;
        RECT  4.685000 197.225000  4.885000 197.425000 ;
        RECT  4.685000 197.630000  4.885000 197.830000 ;
        RECT  4.685000 198.035000  4.885000 198.235000 ;
        RECT  4.685000 198.440000  4.885000 198.640000 ;
        RECT  4.685000 198.845000  4.885000 199.045000 ;
        RECT  4.685000 199.250000  4.885000 199.450000 ;
        RECT  4.685000 199.655000  4.885000 199.855000 ;
        RECT  5.070000  25.910000  5.270000  26.110000 ;
        RECT  5.070000  26.340000  5.270000  26.540000 ;
        RECT  5.070000  26.770000  5.270000  26.970000 ;
        RECT  5.070000  27.200000  5.270000  27.400000 ;
        RECT  5.070000  27.630000  5.270000  27.830000 ;
        RECT  5.070000  28.060000  5.270000  28.260000 ;
        RECT  5.070000  28.490000  5.270000  28.690000 ;
        RECT  5.070000  28.920000  5.270000  29.120000 ;
        RECT  5.070000  29.350000  5.270000  29.550000 ;
        RECT  5.070000  29.780000  5.270000  29.980000 ;
        RECT  5.070000  30.210000  5.270000  30.410000 ;
        RECT  5.085000 175.995000  5.285000 176.195000 ;
        RECT  5.085000 176.395000  5.285000 176.595000 ;
        RECT  5.085000 176.795000  5.285000 176.995000 ;
        RECT  5.085000 177.195000  5.285000 177.395000 ;
        RECT  5.085000 177.595000  5.285000 177.795000 ;
        RECT  5.085000 177.995000  5.285000 178.195000 ;
        RECT  5.085000 178.395000  5.285000 178.595000 ;
        RECT  5.085000 178.795000  5.285000 178.995000 ;
        RECT  5.085000 179.195000  5.285000 179.395000 ;
        RECT  5.085000 179.595000  5.285000 179.795000 ;
        RECT  5.085000 179.995000  5.285000 180.195000 ;
        RECT  5.085000 180.395000  5.285000 180.595000 ;
        RECT  5.085000 180.795000  5.285000 180.995000 ;
        RECT  5.085000 181.195000  5.285000 181.395000 ;
        RECT  5.085000 181.595000  5.285000 181.795000 ;
        RECT  5.085000 181.995000  5.285000 182.195000 ;
        RECT  5.085000 182.395000  5.285000 182.595000 ;
        RECT  5.085000 182.795000  5.285000 182.995000 ;
        RECT  5.085000 183.195000  5.285000 183.395000 ;
        RECT  5.085000 183.595000  5.285000 183.795000 ;
        RECT  5.085000 183.995000  5.285000 184.195000 ;
        RECT  5.085000 184.395000  5.285000 184.595000 ;
        RECT  5.085000 184.795000  5.285000 184.995000 ;
        RECT  5.085000 185.195000  5.285000 185.395000 ;
        RECT  5.085000 185.595000  5.285000 185.795000 ;
        RECT  5.085000 185.995000  5.285000 186.195000 ;
        RECT  5.085000 186.395000  5.285000 186.595000 ;
        RECT  5.085000 186.795000  5.285000 186.995000 ;
        RECT  5.085000 187.195000  5.285000 187.395000 ;
        RECT  5.085000 187.595000  5.285000 187.795000 ;
        RECT  5.085000 187.995000  5.285000 188.195000 ;
        RECT  5.085000 188.395000  5.285000 188.595000 ;
        RECT  5.085000 188.795000  5.285000 188.995000 ;
        RECT  5.085000 189.195000  5.285000 189.395000 ;
        RECT  5.085000 189.595000  5.285000 189.795000 ;
        RECT  5.085000 189.995000  5.285000 190.195000 ;
        RECT  5.085000 190.395000  5.285000 190.595000 ;
        RECT  5.085000 190.795000  5.285000 190.995000 ;
        RECT  5.085000 191.195000  5.285000 191.395000 ;
        RECT  5.085000 191.595000  5.285000 191.795000 ;
        RECT  5.085000 191.995000  5.285000 192.195000 ;
        RECT  5.085000 192.395000  5.285000 192.595000 ;
        RECT  5.085000 192.795000  5.285000 192.995000 ;
        RECT  5.085000 193.195000  5.285000 193.395000 ;
        RECT  5.085000 193.595000  5.285000 193.795000 ;
        RECT  5.085000 193.995000  5.285000 194.195000 ;
        RECT  5.085000 194.395000  5.285000 194.595000 ;
        RECT  5.085000 194.795000  5.285000 194.995000 ;
        RECT  5.085000 195.200000  5.285000 195.400000 ;
        RECT  5.085000 195.605000  5.285000 195.805000 ;
        RECT  5.085000 196.010000  5.285000 196.210000 ;
        RECT  5.085000 196.415000  5.285000 196.615000 ;
        RECT  5.085000 196.820000  5.285000 197.020000 ;
        RECT  5.085000 197.225000  5.285000 197.425000 ;
        RECT  5.085000 197.630000  5.285000 197.830000 ;
        RECT  5.085000 198.035000  5.285000 198.235000 ;
        RECT  5.085000 198.440000  5.285000 198.640000 ;
        RECT  5.085000 198.845000  5.285000 199.045000 ;
        RECT  5.085000 199.250000  5.285000 199.450000 ;
        RECT  5.085000 199.655000  5.285000 199.855000 ;
        RECT  5.475000  25.910000  5.675000  26.110000 ;
        RECT  5.475000  26.340000  5.675000  26.540000 ;
        RECT  5.475000  26.770000  5.675000  26.970000 ;
        RECT  5.475000  27.200000  5.675000  27.400000 ;
        RECT  5.475000  27.630000  5.675000  27.830000 ;
        RECT  5.475000  28.060000  5.675000  28.260000 ;
        RECT  5.475000  28.490000  5.675000  28.690000 ;
        RECT  5.475000  28.920000  5.675000  29.120000 ;
        RECT  5.475000  29.350000  5.675000  29.550000 ;
        RECT  5.475000  29.780000  5.675000  29.980000 ;
        RECT  5.475000  30.210000  5.675000  30.410000 ;
        RECT  5.485000 175.995000  5.685000 176.195000 ;
        RECT  5.485000 176.395000  5.685000 176.595000 ;
        RECT  5.485000 176.795000  5.685000 176.995000 ;
        RECT  5.485000 177.195000  5.685000 177.395000 ;
        RECT  5.485000 177.595000  5.685000 177.795000 ;
        RECT  5.485000 177.995000  5.685000 178.195000 ;
        RECT  5.485000 178.395000  5.685000 178.595000 ;
        RECT  5.485000 178.795000  5.685000 178.995000 ;
        RECT  5.485000 179.195000  5.685000 179.395000 ;
        RECT  5.485000 179.595000  5.685000 179.795000 ;
        RECT  5.485000 179.995000  5.685000 180.195000 ;
        RECT  5.485000 180.395000  5.685000 180.595000 ;
        RECT  5.485000 180.795000  5.685000 180.995000 ;
        RECT  5.485000 181.195000  5.685000 181.395000 ;
        RECT  5.485000 181.595000  5.685000 181.795000 ;
        RECT  5.485000 181.995000  5.685000 182.195000 ;
        RECT  5.485000 182.395000  5.685000 182.595000 ;
        RECT  5.485000 182.795000  5.685000 182.995000 ;
        RECT  5.485000 183.195000  5.685000 183.395000 ;
        RECT  5.485000 183.595000  5.685000 183.795000 ;
        RECT  5.485000 183.995000  5.685000 184.195000 ;
        RECT  5.485000 184.395000  5.685000 184.595000 ;
        RECT  5.485000 184.795000  5.685000 184.995000 ;
        RECT  5.485000 185.195000  5.685000 185.395000 ;
        RECT  5.485000 185.595000  5.685000 185.795000 ;
        RECT  5.485000 185.995000  5.685000 186.195000 ;
        RECT  5.485000 186.395000  5.685000 186.595000 ;
        RECT  5.485000 186.795000  5.685000 186.995000 ;
        RECT  5.485000 187.195000  5.685000 187.395000 ;
        RECT  5.485000 187.595000  5.685000 187.795000 ;
        RECT  5.485000 187.995000  5.685000 188.195000 ;
        RECT  5.485000 188.395000  5.685000 188.595000 ;
        RECT  5.485000 188.795000  5.685000 188.995000 ;
        RECT  5.485000 189.195000  5.685000 189.395000 ;
        RECT  5.485000 189.595000  5.685000 189.795000 ;
        RECT  5.485000 189.995000  5.685000 190.195000 ;
        RECT  5.485000 190.395000  5.685000 190.595000 ;
        RECT  5.485000 190.795000  5.685000 190.995000 ;
        RECT  5.485000 191.195000  5.685000 191.395000 ;
        RECT  5.485000 191.595000  5.685000 191.795000 ;
        RECT  5.485000 191.995000  5.685000 192.195000 ;
        RECT  5.485000 192.395000  5.685000 192.595000 ;
        RECT  5.485000 192.795000  5.685000 192.995000 ;
        RECT  5.485000 193.195000  5.685000 193.395000 ;
        RECT  5.485000 193.595000  5.685000 193.795000 ;
        RECT  5.485000 193.995000  5.685000 194.195000 ;
        RECT  5.485000 194.395000  5.685000 194.595000 ;
        RECT  5.485000 194.795000  5.685000 194.995000 ;
        RECT  5.485000 195.200000  5.685000 195.400000 ;
        RECT  5.485000 195.605000  5.685000 195.805000 ;
        RECT  5.485000 196.010000  5.685000 196.210000 ;
        RECT  5.485000 196.415000  5.685000 196.615000 ;
        RECT  5.485000 196.820000  5.685000 197.020000 ;
        RECT  5.485000 197.225000  5.685000 197.425000 ;
        RECT  5.485000 197.630000  5.685000 197.830000 ;
        RECT  5.485000 198.035000  5.685000 198.235000 ;
        RECT  5.485000 198.440000  5.685000 198.640000 ;
        RECT  5.485000 198.845000  5.685000 199.045000 ;
        RECT  5.485000 199.250000  5.685000 199.450000 ;
        RECT  5.485000 199.655000  5.685000 199.855000 ;
        RECT  5.880000  25.910000  6.080000  26.110000 ;
        RECT  5.880000  26.340000  6.080000  26.540000 ;
        RECT  5.880000  26.770000  6.080000  26.970000 ;
        RECT  5.880000  27.200000  6.080000  27.400000 ;
        RECT  5.880000  27.630000  6.080000  27.830000 ;
        RECT  5.880000  28.060000  6.080000  28.260000 ;
        RECT  5.880000  28.490000  6.080000  28.690000 ;
        RECT  5.880000  28.920000  6.080000  29.120000 ;
        RECT  5.880000  29.350000  6.080000  29.550000 ;
        RECT  5.880000  29.780000  6.080000  29.980000 ;
        RECT  5.880000  30.210000  6.080000  30.410000 ;
        RECT  5.885000 175.995000  6.085000 176.195000 ;
        RECT  5.885000 176.395000  6.085000 176.595000 ;
        RECT  5.885000 176.795000  6.085000 176.995000 ;
        RECT  5.885000 177.195000  6.085000 177.395000 ;
        RECT  5.885000 177.595000  6.085000 177.795000 ;
        RECT  5.885000 177.995000  6.085000 178.195000 ;
        RECT  5.885000 178.395000  6.085000 178.595000 ;
        RECT  5.885000 178.795000  6.085000 178.995000 ;
        RECT  5.885000 179.195000  6.085000 179.395000 ;
        RECT  5.885000 179.595000  6.085000 179.795000 ;
        RECT  5.885000 179.995000  6.085000 180.195000 ;
        RECT  5.885000 180.395000  6.085000 180.595000 ;
        RECT  5.885000 180.795000  6.085000 180.995000 ;
        RECT  5.885000 181.195000  6.085000 181.395000 ;
        RECT  5.885000 181.595000  6.085000 181.795000 ;
        RECT  5.885000 181.995000  6.085000 182.195000 ;
        RECT  5.885000 182.395000  6.085000 182.595000 ;
        RECT  5.885000 182.795000  6.085000 182.995000 ;
        RECT  5.885000 183.195000  6.085000 183.395000 ;
        RECT  5.885000 183.595000  6.085000 183.795000 ;
        RECT  5.885000 183.995000  6.085000 184.195000 ;
        RECT  5.885000 184.395000  6.085000 184.595000 ;
        RECT  5.885000 184.795000  6.085000 184.995000 ;
        RECT  5.885000 185.195000  6.085000 185.395000 ;
        RECT  5.885000 185.595000  6.085000 185.795000 ;
        RECT  5.885000 185.995000  6.085000 186.195000 ;
        RECT  5.885000 186.395000  6.085000 186.595000 ;
        RECT  5.885000 186.795000  6.085000 186.995000 ;
        RECT  5.885000 187.195000  6.085000 187.395000 ;
        RECT  5.885000 187.595000  6.085000 187.795000 ;
        RECT  5.885000 187.995000  6.085000 188.195000 ;
        RECT  5.885000 188.395000  6.085000 188.595000 ;
        RECT  5.885000 188.795000  6.085000 188.995000 ;
        RECT  5.885000 189.195000  6.085000 189.395000 ;
        RECT  5.885000 189.595000  6.085000 189.795000 ;
        RECT  5.885000 189.995000  6.085000 190.195000 ;
        RECT  5.885000 190.395000  6.085000 190.595000 ;
        RECT  5.885000 190.795000  6.085000 190.995000 ;
        RECT  5.885000 191.195000  6.085000 191.395000 ;
        RECT  5.885000 191.595000  6.085000 191.795000 ;
        RECT  5.885000 191.995000  6.085000 192.195000 ;
        RECT  5.885000 192.395000  6.085000 192.595000 ;
        RECT  5.885000 192.795000  6.085000 192.995000 ;
        RECT  5.885000 193.195000  6.085000 193.395000 ;
        RECT  5.885000 193.595000  6.085000 193.795000 ;
        RECT  5.885000 193.995000  6.085000 194.195000 ;
        RECT  5.885000 194.395000  6.085000 194.595000 ;
        RECT  5.885000 194.795000  6.085000 194.995000 ;
        RECT  5.885000 195.200000  6.085000 195.400000 ;
        RECT  5.885000 195.605000  6.085000 195.805000 ;
        RECT  5.885000 196.010000  6.085000 196.210000 ;
        RECT  5.885000 196.415000  6.085000 196.615000 ;
        RECT  5.885000 196.820000  6.085000 197.020000 ;
        RECT  5.885000 197.225000  6.085000 197.425000 ;
        RECT  5.885000 197.630000  6.085000 197.830000 ;
        RECT  5.885000 198.035000  6.085000 198.235000 ;
        RECT  5.885000 198.440000  6.085000 198.640000 ;
        RECT  5.885000 198.845000  6.085000 199.045000 ;
        RECT  5.885000 199.250000  6.085000 199.450000 ;
        RECT  5.885000 199.655000  6.085000 199.855000 ;
        RECT  6.285000  25.910000  6.485000  26.110000 ;
        RECT  6.285000  26.340000  6.485000  26.540000 ;
        RECT  6.285000  26.770000  6.485000  26.970000 ;
        RECT  6.285000  27.200000  6.485000  27.400000 ;
        RECT  6.285000  27.630000  6.485000  27.830000 ;
        RECT  6.285000  28.060000  6.485000  28.260000 ;
        RECT  6.285000  28.490000  6.485000  28.690000 ;
        RECT  6.285000  28.920000  6.485000  29.120000 ;
        RECT  6.285000  29.350000  6.485000  29.550000 ;
        RECT  6.285000  29.780000  6.485000  29.980000 ;
        RECT  6.285000  30.210000  6.485000  30.410000 ;
        RECT  6.285000 175.995000  6.485000 176.195000 ;
        RECT  6.285000 176.395000  6.485000 176.595000 ;
        RECT  6.285000 176.795000  6.485000 176.995000 ;
        RECT  6.285000 177.195000  6.485000 177.395000 ;
        RECT  6.285000 177.595000  6.485000 177.795000 ;
        RECT  6.285000 177.995000  6.485000 178.195000 ;
        RECT  6.285000 178.395000  6.485000 178.595000 ;
        RECT  6.285000 178.795000  6.485000 178.995000 ;
        RECT  6.285000 179.195000  6.485000 179.395000 ;
        RECT  6.285000 179.595000  6.485000 179.795000 ;
        RECT  6.285000 179.995000  6.485000 180.195000 ;
        RECT  6.285000 180.395000  6.485000 180.595000 ;
        RECT  6.285000 180.795000  6.485000 180.995000 ;
        RECT  6.285000 181.195000  6.485000 181.395000 ;
        RECT  6.285000 181.595000  6.485000 181.795000 ;
        RECT  6.285000 181.995000  6.485000 182.195000 ;
        RECT  6.285000 182.395000  6.485000 182.595000 ;
        RECT  6.285000 182.795000  6.485000 182.995000 ;
        RECT  6.285000 183.195000  6.485000 183.395000 ;
        RECT  6.285000 183.595000  6.485000 183.795000 ;
        RECT  6.285000 183.995000  6.485000 184.195000 ;
        RECT  6.285000 184.395000  6.485000 184.595000 ;
        RECT  6.285000 184.795000  6.485000 184.995000 ;
        RECT  6.285000 185.195000  6.485000 185.395000 ;
        RECT  6.285000 185.595000  6.485000 185.795000 ;
        RECT  6.285000 185.995000  6.485000 186.195000 ;
        RECT  6.285000 186.395000  6.485000 186.595000 ;
        RECT  6.285000 186.795000  6.485000 186.995000 ;
        RECT  6.285000 187.195000  6.485000 187.395000 ;
        RECT  6.285000 187.595000  6.485000 187.795000 ;
        RECT  6.285000 187.995000  6.485000 188.195000 ;
        RECT  6.285000 188.395000  6.485000 188.595000 ;
        RECT  6.285000 188.795000  6.485000 188.995000 ;
        RECT  6.285000 189.195000  6.485000 189.395000 ;
        RECT  6.285000 189.595000  6.485000 189.795000 ;
        RECT  6.285000 189.995000  6.485000 190.195000 ;
        RECT  6.285000 190.395000  6.485000 190.595000 ;
        RECT  6.285000 190.795000  6.485000 190.995000 ;
        RECT  6.285000 191.195000  6.485000 191.395000 ;
        RECT  6.285000 191.595000  6.485000 191.795000 ;
        RECT  6.285000 191.995000  6.485000 192.195000 ;
        RECT  6.285000 192.395000  6.485000 192.595000 ;
        RECT  6.285000 192.795000  6.485000 192.995000 ;
        RECT  6.285000 193.195000  6.485000 193.395000 ;
        RECT  6.285000 193.595000  6.485000 193.795000 ;
        RECT  6.285000 193.995000  6.485000 194.195000 ;
        RECT  6.285000 194.395000  6.485000 194.595000 ;
        RECT  6.285000 194.795000  6.485000 194.995000 ;
        RECT  6.285000 195.200000  6.485000 195.400000 ;
        RECT  6.285000 195.605000  6.485000 195.805000 ;
        RECT  6.285000 196.010000  6.485000 196.210000 ;
        RECT  6.285000 196.415000  6.485000 196.615000 ;
        RECT  6.285000 196.820000  6.485000 197.020000 ;
        RECT  6.285000 197.225000  6.485000 197.425000 ;
        RECT  6.285000 197.630000  6.485000 197.830000 ;
        RECT  6.285000 198.035000  6.485000 198.235000 ;
        RECT  6.285000 198.440000  6.485000 198.640000 ;
        RECT  6.285000 198.845000  6.485000 199.045000 ;
        RECT  6.285000 199.250000  6.485000 199.450000 ;
        RECT  6.285000 199.655000  6.485000 199.855000 ;
        RECT  6.685000 175.995000  6.885000 176.195000 ;
        RECT  6.685000 176.395000  6.885000 176.595000 ;
        RECT  6.685000 176.795000  6.885000 176.995000 ;
        RECT  6.685000 177.195000  6.885000 177.395000 ;
        RECT  6.685000 177.595000  6.885000 177.795000 ;
        RECT  6.685000 177.995000  6.885000 178.195000 ;
        RECT  6.685000 178.395000  6.885000 178.595000 ;
        RECT  6.685000 178.795000  6.885000 178.995000 ;
        RECT  6.685000 179.195000  6.885000 179.395000 ;
        RECT  6.685000 179.595000  6.885000 179.795000 ;
        RECT  6.685000 179.995000  6.885000 180.195000 ;
        RECT  6.685000 180.395000  6.885000 180.595000 ;
        RECT  6.685000 180.795000  6.885000 180.995000 ;
        RECT  6.685000 181.195000  6.885000 181.395000 ;
        RECT  6.685000 181.595000  6.885000 181.795000 ;
        RECT  6.685000 181.995000  6.885000 182.195000 ;
        RECT  6.685000 182.395000  6.885000 182.595000 ;
        RECT  6.685000 182.795000  6.885000 182.995000 ;
        RECT  6.685000 183.195000  6.885000 183.395000 ;
        RECT  6.685000 183.595000  6.885000 183.795000 ;
        RECT  6.685000 183.995000  6.885000 184.195000 ;
        RECT  6.685000 184.395000  6.885000 184.595000 ;
        RECT  6.685000 184.795000  6.885000 184.995000 ;
        RECT  6.685000 185.195000  6.885000 185.395000 ;
        RECT  6.685000 185.595000  6.885000 185.795000 ;
        RECT  6.685000 185.995000  6.885000 186.195000 ;
        RECT  6.685000 186.395000  6.885000 186.595000 ;
        RECT  6.685000 186.795000  6.885000 186.995000 ;
        RECT  6.685000 187.195000  6.885000 187.395000 ;
        RECT  6.685000 187.595000  6.885000 187.795000 ;
        RECT  6.685000 187.995000  6.885000 188.195000 ;
        RECT  6.685000 188.395000  6.885000 188.595000 ;
        RECT  6.685000 188.795000  6.885000 188.995000 ;
        RECT  6.685000 189.195000  6.885000 189.395000 ;
        RECT  6.685000 189.595000  6.885000 189.795000 ;
        RECT  6.685000 189.995000  6.885000 190.195000 ;
        RECT  6.685000 190.395000  6.885000 190.595000 ;
        RECT  6.685000 190.795000  6.885000 190.995000 ;
        RECT  6.685000 191.195000  6.885000 191.395000 ;
        RECT  6.685000 191.595000  6.885000 191.795000 ;
        RECT  6.685000 191.995000  6.885000 192.195000 ;
        RECT  6.685000 192.395000  6.885000 192.595000 ;
        RECT  6.685000 192.795000  6.885000 192.995000 ;
        RECT  6.685000 193.195000  6.885000 193.395000 ;
        RECT  6.685000 193.595000  6.885000 193.795000 ;
        RECT  6.685000 193.995000  6.885000 194.195000 ;
        RECT  6.685000 194.395000  6.885000 194.595000 ;
        RECT  6.685000 194.795000  6.885000 194.995000 ;
        RECT  6.685000 195.200000  6.885000 195.400000 ;
        RECT  6.685000 195.605000  6.885000 195.805000 ;
        RECT  6.685000 196.010000  6.885000 196.210000 ;
        RECT  6.685000 196.415000  6.885000 196.615000 ;
        RECT  6.685000 196.820000  6.885000 197.020000 ;
        RECT  6.685000 197.225000  6.885000 197.425000 ;
        RECT  6.685000 197.630000  6.885000 197.830000 ;
        RECT  6.685000 198.035000  6.885000 198.235000 ;
        RECT  6.685000 198.440000  6.885000 198.640000 ;
        RECT  6.685000 198.845000  6.885000 199.045000 ;
        RECT  6.685000 199.250000  6.885000 199.450000 ;
        RECT  6.685000 199.655000  6.885000 199.855000 ;
        RECT  6.690000  25.910000  6.890000  26.110000 ;
        RECT  6.690000  26.340000  6.890000  26.540000 ;
        RECT  6.690000  26.770000  6.890000  26.970000 ;
        RECT  6.690000  27.200000  6.890000  27.400000 ;
        RECT  6.690000  27.630000  6.890000  27.830000 ;
        RECT  6.690000  28.060000  6.890000  28.260000 ;
        RECT  6.690000  28.490000  6.890000  28.690000 ;
        RECT  6.690000  28.920000  6.890000  29.120000 ;
        RECT  6.690000  29.350000  6.890000  29.550000 ;
        RECT  6.690000  29.780000  6.890000  29.980000 ;
        RECT  6.690000  30.210000  6.890000  30.410000 ;
        RECT  7.085000 175.995000  7.285000 176.195000 ;
        RECT  7.085000 176.395000  7.285000 176.595000 ;
        RECT  7.085000 176.795000  7.285000 176.995000 ;
        RECT  7.085000 177.195000  7.285000 177.395000 ;
        RECT  7.085000 177.595000  7.285000 177.795000 ;
        RECT  7.085000 177.995000  7.285000 178.195000 ;
        RECT  7.085000 178.395000  7.285000 178.595000 ;
        RECT  7.085000 178.795000  7.285000 178.995000 ;
        RECT  7.085000 179.195000  7.285000 179.395000 ;
        RECT  7.085000 179.595000  7.285000 179.795000 ;
        RECT  7.085000 179.995000  7.285000 180.195000 ;
        RECT  7.085000 180.395000  7.285000 180.595000 ;
        RECT  7.085000 180.795000  7.285000 180.995000 ;
        RECT  7.085000 181.195000  7.285000 181.395000 ;
        RECT  7.085000 181.595000  7.285000 181.795000 ;
        RECT  7.085000 181.995000  7.285000 182.195000 ;
        RECT  7.085000 182.395000  7.285000 182.595000 ;
        RECT  7.085000 182.795000  7.285000 182.995000 ;
        RECT  7.085000 183.195000  7.285000 183.395000 ;
        RECT  7.085000 183.595000  7.285000 183.795000 ;
        RECT  7.085000 183.995000  7.285000 184.195000 ;
        RECT  7.085000 184.395000  7.285000 184.595000 ;
        RECT  7.085000 184.795000  7.285000 184.995000 ;
        RECT  7.085000 185.195000  7.285000 185.395000 ;
        RECT  7.085000 185.595000  7.285000 185.795000 ;
        RECT  7.085000 185.995000  7.285000 186.195000 ;
        RECT  7.085000 186.395000  7.285000 186.595000 ;
        RECT  7.085000 186.795000  7.285000 186.995000 ;
        RECT  7.085000 187.195000  7.285000 187.395000 ;
        RECT  7.085000 187.595000  7.285000 187.795000 ;
        RECT  7.085000 187.995000  7.285000 188.195000 ;
        RECT  7.085000 188.395000  7.285000 188.595000 ;
        RECT  7.085000 188.795000  7.285000 188.995000 ;
        RECT  7.085000 189.195000  7.285000 189.395000 ;
        RECT  7.085000 189.595000  7.285000 189.795000 ;
        RECT  7.085000 189.995000  7.285000 190.195000 ;
        RECT  7.085000 190.395000  7.285000 190.595000 ;
        RECT  7.085000 190.795000  7.285000 190.995000 ;
        RECT  7.085000 191.195000  7.285000 191.395000 ;
        RECT  7.085000 191.595000  7.285000 191.795000 ;
        RECT  7.085000 191.995000  7.285000 192.195000 ;
        RECT  7.085000 192.395000  7.285000 192.595000 ;
        RECT  7.085000 192.795000  7.285000 192.995000 ;
        RECT  7.085000 193.195000  7.285000 193.395000 ;
        RECT  7.085000 193.595000  7.285000 193.795000 ;
        RECT  7.085000 193.995000  7.285000 194.195000 ;
        RECT  7.085000 194.395000  7.285000 194.595000 ;
        RECT  7.085000 194.795000  7.285000 194.995000 ;
        RECT  7.085000 195.200000  7.285000 195.400000 ;
        RECT  7.085000 195.605000  7.285000 195.805000 ;
        RECT  7.085000 196.010000  7.285000 196.210000 ;
        RECT  7.085000 196.415000  7.285000 196.615000 ;
        RECT  7.085000 196.820000  7.285000 197.020000 ;
        RECT  7.085000 197.225000  7.285000 197.425000 ;
        RECT  7.085000 197.630000  7.285000 197.830000 ;
        RECT  7.085000 198.035000  7.285000 198.235000 ;
        RECT  7.085000 198.440000  7.285000 198.640000 ;
        RECT  7.085000 198.845000  7.285000 199.045000 ;
        RECT  7.085000 199.250000  7.285000 199.450000 ;
        RECT  7.085000 199.655000  7.285000 199.855000 ;
        RECT  7.095000  25.910000  7.295000  26.110000 ;
        RECT  7.095000  26.340000  7.295000  26.540000 ;
        RECT  7.095000  26.770000  7.295000  26.970000 ;
        RECT  7.095000  27.200000  7.295000  27.400000 ;
        RECT  7.095000  27.630000  7.295000  27.830000 ;
        RECT  7.095000  28.060000  7.295000  28.260000 ;
        RECT  7.095000  28.490000  7.295000  28.690000 ;
        RECT  7.095000  28.920000  7.295000  29.120000 ;
        RECT  7.095000  29.350000  7.295000  29.550000 ;
        RECT  7.095000  29.780000  7.295000  29.980000 ;
        RECT  7.095000  30.210000  7.295000  30.410000 ;
        RECT  7.485000 175.995000  7.685000 176.195000 ;
        RECT  7.485000 176.395000  7.685000 176.595000 ;
        RECT  7.485000 176.795000  7.685000 176.995000 ;
        RECT  7.485000 177.195000  7.685000 177.395000 ;
        RECT  7.485000 177.595000  7.685000 177.795000 ;
        RECT  7.485000 177.995000  7.685000 178.195000 ;
        RECT  7.485000 178.395000  7.685000 178.595000 ;
        RECT  7.485000 178.795000  7.685000 178.995000 ;
        RECT  7.485000 179.195000  7.685000 179.395000 ;
        RECT  7.485000 179.595000  7.685000 179.795000 ;
        RECT  7.485000 179.995000  7.685000 180.195000 ;
        RECT  7.485000 180.395000  7.685000 180.595000 ;
        RECT  7.485000 180.795000  7.685000 180.995000 ;
        RECT  7.485000 181.195000  7.685000 181.395000 ;
        RECT  7.485000 181.595000  7.685000 181.795000 ;
        RECT  7.485000 181.995000  7.685000 182.195000 ;
        RECT  7.485000 182.395000  7.685000 182.595000 ;
        RECT  7.485000 182.795000  7.685000 182.995000 ;
        RECT  7.485000 183.195000  7.685000 183.395000 ;
        RECT  7.485000 183.595000  7.685000 183.795000 ;
        RECT  7.485000 183.995000  7.685000 184.195000 ;
        RECT  7.485000 184.395000  7.685000 184.595000 ;
        RECT  7.485000 184.795000  7.685000 184.995000 ;
        RECT  7.485000 185.195000  7.685000 185.395000 ;
        RECT  7.485000 185.595000  7.685000 185.795000 ;
        RECT  7.485000 185.995000  7.685000 186.195000 ;
        RECT  7.485000 186.395000  7.685000 186.595000 ;
        RECT  7.485000 186.795000  7.685000 186.995000 ;
        RECT  7.485000 187.195000  7.685000 187.395000 ;
        RECT  7.485000 187.595000  7.685000 187.795000 ;
        RECT  7.485000 187.995000  7.685000 188.195000 ;
        RECT  7.485000 188.395000  7.685000 188.595000 ;
        RECT  7.485000 188.795000  7.685000 188.995000 ;
        RECT  7.485000 189.195000  7.685000 189.395000 ;
        RECT  7.485000 189.595000  7.685000 189.795000 ;
        RECT  7.485000 189.995000  7.685000 190.195000 ;
        RECT  7.485000 190.395000  7.685000 190.595000 ;
        RECT  7.485000 190.795000  7.685000 190.995000 ;
        RECT  7.485000 191.195000  7.685000 191.395000 ;
        RECT  7.485000 191.595000  7.685000 191.795000 ;
        RECT  7.485000 191.995000  7.685000 192.195000 ;
        RECT  7.485000 192.395000  7.685000 192.595000 ;
        RECT  7.485000 192.795000  7.685000 192.995000 ;
        RECT  7.485000 193.195000  7.685000 193.395000 ;
        RECT  7.485000 193.595000  7.685000 193.795000 ;
        RECT  7.485000 193.995000  7.685000 194.195000 ;
        RECT  7.485000 194.395000  7.685000 194.595000 ;
        RECT  7.485000 194.795000  7.685000 194.995000 ;
        RECT  7.485000 195.200000  7.685000 195.400000 ;
        RECT  7.485000 195.605000  7.685000 195.805000 ;
        RECT  7.485000 196.010000  7.685000 196.210000 ;
        RECT  7.485000 196.415000  7.685000 196.615000 ;
        RECT  7.485000 196.820000  7.685000 197.020000 ;
        RECT  7.485000 197.225000  7.685000 197.425000 ;
        RECT  7.485000 197.630000  7.685000 197.830000 ;
        RECT  7.485000 198.035000  7.685000 198.235000 ;
        RECT  7.485000 198.440000  7.685000 198.640000 ;
        RECT  7.485000 198.845000  7.685000 199.045000 ;
        RECT  7.485000 199.250000  7.685000 199.450000 ;
        RECT  7.485000 199.655000  7.685000 199.855000 ;
        RECT  7.500000  25.910000  7.700000  26.110000 ;
        RECT  7.500000  26.340000  7.700000  26.540000 ;
        RECT  7.500000  26.770000  7.700000  26.970000 ;
        RECT  7.500000  27.200000  7.700000  27.400000 ;
        RECT  7.500000  27.630000  7.700000  27.830000 ;
        RECT  7.500000  28.060000  7.700000  28.260000 ;
        RECT  7.500000  28.490000  7.700000  28.690000 ;
        RECT  7.500000  28.920000  7.700000  29.120000 ;
        RECT  7.500000  29.350000  7.700000  29.550000 ;
        RECT  7.500000  29.780000  7.700000  29.980000 ;
        RECT  7.500000  30.210000  7.700000  30.410000 ;
        RECT  7.885000 175.995000  8.085000 176.195000 ;
        RECT  7.885000 176.395000  8.085000 176.595000 ;
        RECT  7.885000 176.795000  8.085000 176.995000 ;
        RECT  7.885000 177.195000  8.085000 177.395000 ;
        RECT  7.885000 177.595000  8.085000 177.795000 ;
        RECT  7.885000 177.995000  8.085000 178.195000 ;
        RECT  7.885000 178.395000  8.085000 178.595000 ;
        RECT  7.885000 178.795000  8.085000 178.995000 ;
        RECT  7.885000 179.195000  8.085000 179.395000 ;
        RECT  7.885000 179.595000  8.085000 179.795000 ;
        RECT  7.885000 179.995000  8.085000 180.195000 ;
        RECT  7.885000 180.395000  8.085000 180.595000 ;
        RECT  7.885000 180.795000  8.085000 180.995000 ;
        RECT  7.885000 181.195000  8.085000 181.395000 ;
        RECT  7.885000 181.595000  8.085000 181.795000 ;
        RECT  7.885000 181.995000  8.085000 182.195000 ;
        RECT  7.885000 182.395000  8.085000 182.595000 ;
        RECT  7.885000 182.795000  8.085000 182.995000 ;
        RECT  7.885000 183.195000  8.085000 183.395000 ;
        RECT  7.885000 183.595000  8.085000 183.795000 ;
        RECT  7.885000 183.995000  8.085000 184.195000 ;
        RECT  7.885000 184.395000  8.085000 184.595000 ;
        RECT  7.885000 184.795000  8.085000 184.995000 ;
        RECT  7.885000 185.195000  8.085000 185.395000 ;
        RECT  7.885000 185.595000  8.085000 185.795000 ;
        RECT  7.885000 185.995000  8.085000 186.195000 ;
        RECT  7.885000 186.395000  8.085000 186.595000 ;
        RECT  7.885000 186.795000  8.085000 186.995000 ;
        RECT  7.885000 187.195000  8.085000 187.395000 ;
        RECT  7.885000 187.595000  8.085000 187.795000 ;
        RECT  7.885000 187.995000  8.085000 188.195000 ;
        RECT  7.885000 188.395000  8.085000 188.595000 ;
        RECT  7.885000 188.795000  8.085000 188.995000 ;
        RECT  7.885000 189.195000  8.085000 189.395000 ;
        RECT  7.885000 189.595000  8.085000 189.795000 ;
        RECT  7.885000 189.995000  8.085000 190.195000 ;
        RECT  7.885000 190.395000  8.085000 190.595000 ;
        RECT  7.885000 190.795000  8.085000 190.995000 ;
        RECT  7.885000 191.195000  8.085000 191.395000 ;
        RECT  7.885000 191.595000  8.085000 191.795000 ;
        RECT  7.885000 191.995000  8.085000 192.195000 ;
        RECT  7.885000 192.395000  8.085000 192.595000 ;
        RECT  7.885000 192.795000  8.085000 192.995000 ;
        RECT  7.885000 193.195000  8.085000 193.395000 ;
        RECT  7.885000 193.595000  8.085000 193.795000 ;
        RECT  7.885000 193.995000  8.085000 194.195000 ;
        RECT  7.885000 194.395000  8.085000 194.595000 ;
        RECT  7.885000 194.795000  8.085000 194.995000 ;
        RECT  7.885000 195.200000  8.085000 195.400000 ;
        RECT  7.885000 195.605000  8.085000 195.805000 ;
        RECT  7.885000 196.010000  8.085000 196.210000 ;
        RECT  7.885000 196.415000  8.085000 196.615000 ;
        RECT  7.885000 196.820000  8.085000 197.020000 ;
        RECT  7.885000 197.225000  8.085000 197.425000 ;
        RECT  7.885000 197.630000  8.085000 197.830000 ;
        RECT  7.885000 198.035000  8.085000 198.235000 ;
        RECT  7.885000 198.440000  8.085000 198.640000 ;
        RECT  7.885000 198.845000  8.085000 199.045000 ;
        RECT  7.885000 199.250000  8.085000 199.450000 ;
        RECT  7.885000 199.655000  8.085000 199.855000 ;
        RECT  7.905000  25.910000  8.105000  26.110000 ;
        RECT  7.905000  26.340000  8.105000  26.540000 ;
        RECT  7.905000  26.770000  8.105000  26.970000 ;
        RECT  7.905000  27.200000  8.105000  27.400000 ;
        RECT  7.905000  27.630000  8.105000  27.830000 ;
        RECT  7.905000  28.060000  8.105000  28.260000 ;
        RECT  7.905000  28.490000  8.105000  28.690000 ;
        RECT  7.905000  28.920000  8.105000  29.120000 ;
        RECT  7.905000  29.350000  8.105000  29.550000 ;
        RECT  7.905000  29.780000  8.105000  29.980000 ;
        RECT  7.905000  30.210000  8.105000  30.410000 ;
        RECT  8.285000 175.995000  8.485000 176.195000 ;
        RECT  8.285000 176.395000  8.485000 176.595000 ;
        RECT  8.285000 176.795000  8.485000 176.995000 ;
        RECT  8.285000 177.195000  8.485000 177.395000 ;
        RECT  8.285000 177.595000  8.485000 177.795000 ;
        RECT  8.285000 177.995000  8.485000 178.195000 ;
        RECT  8.285000 178.395000  8.485000 178.595000 ;
        RECT  8.285000 178.795000  8.485000 178.995000 ;
        RECT  8.285000 179.195000  8.485000 179.395000 ;
        RECT  8.285000 179.595000  8.485000 179.795000 ;
        RECT  8.285000 179.995000  8.485000 180.195000 ;
        RECT  8.285000 180.395000  8.485000 180.595000 ;
        RECT  8.285000 180.795000  8.485000 180.995000 ;
        RECT  8.285000 181.195000  8.485000 181.395000 ;
        RECT  8.285000 181.595000  8.485000 181.795000 ;
        RECT  8.285000 181.995000  8.485000 182.195000 ;
        RECT  8.285000 182.395000  8.485000 182.595000 ;
        RECT  8.285000 182.795000  8.485000 182.995000 ;
        RECT  8.285000 183.195000  8.485000 183.395000 ;
        RECT  8.285000 183.595000  8.485000 183.795000 ;
        RECT  8.285000 183.995000  8.485000 184.195000 ;
        RECT  8.285000 184.395000  8.485000 184.595000 ;
        RECT  8.285000 184.795000  8.485000 184.995000 ;
        RECT  8.285000 185.195000  8.485000 185.395000 ;
        RECT  8.285000 185.595000  8.485000 185.795000 ;
        RECT  8.285000 185.995000  8.485000 186.195000 ;
        RECT  8.285000 186.395000  8.485000 186.595000 ;
        RECT  8.285000 186.795000  8.485000 186.995000 ;
        RECT  8.285000 187.195000  8.485000 187.395000 ;
        RECT  8.285000 187.595000  8.485000 187.795000 ;
        RECT  8.285000 187.995000  8.485000 188.195000 ;
        RECT  8.285000 188.395000  8.485000 188.595000 ;
        RECT  8.285000 188.795000  8.485000 188.995000 ;
        RECT  8.285000 189.195000  8.485000 189.395000 ;
        RECT  8.285000 189.595000  8.485000 189.795000 ;
        RECT  8.285000 189.995000  8.485000 190.195000 ;
        RECT  8.285000 190.395000  8.485000 190.595000 ;
        RECT  8.285000 190.795000  8.485000 190.995000 ;
        RECT  8.285000 191.195000  8.485000 191.395000 ;
        RECT  8.285000 191.595000  8.485000 191.795000 ;
        RECT  8.285000 191.995000  8.485000 192.195000 ;
        RECT  8.285000 192.395000  8.485000 192.595000 ;
        RECT  8.285000 192.795000  8.485000 192.995000 ;
        RECT  8.285000 193.195000  8.485000 193.395000 ;
        RECT  8.285000 193.595000  8.485000 193.795000 ;
        RECT  8.285000 193.995000  8.485000 194.195000 ;
        RECT  8.285000 194.395000  8.485000 194.595000 ;
        RECT  8.285000 194.795000  8.485000 194.995000 ;
        RECT  8.285000 195.200000  8.485000 195.400000 ;
        RECT  8.285000 195.605000  8.485000 195.805000 ;
        RECT  8.285000 196.010000  8.485000 196.210000 ;
        RECT  8.285000 196.415000  8.485000 196.615000 ;
        RECT  8.285000 196.820000  8.485000 197.020000 ;
        RECT  8.285000 197.225000  8.485000 197.425000 ;
        RECT  8.285000 197.630000  8.485000 197.830000 ;
        RECT  8.285000 198.035000  8.485000 198.235000 ;
        RECT  8.285000 198.440000  8.485000 198.640000 ;
        RECT  8.285000 198.845000  8.485000 199.045000 ;
        RECT  8.285000 199.250000  8.485000 199.450000 ;
        RECT  8.285000 199.655000  8.485000 199.855000 ;
        RECT  8.310000  25.910000  8.510000  26.110000 ;
        RECT  8.310000  26.340000  8.510000  26.540000 ;
        RECT  8.310000  26.770000  8.510000  26.970000 ;
        RECT  8.310000  27.200000  8.510000  27.400000 ;
        RECT  8.310000  27.630000  8.510000  27.830000 ;
        RECT  8.310000  28.060000  8.510000  28.260000 ;
        RECT  8.310000  28.490000  8.510000  28.690000 ;
        RECT  8.310000  28.920000  8.510000  29.120000 ;
        RECT  8.310000  29.350000  8.510000  29.550000 ;
        RECT  8.310000  29.780000  8.510000  29.980000 ;
        RECT  8.310000  30.210000  8.510000  30.410000 ;
        RECT  8.685000 175.995000  8.885000 176.195000 ;
        RECT  8.685000 176.395000  8.885000 176.595000 ;
        RECT  8.685000 176.795000  8.885000 176.995000 ;
        RECT  8.685000 177.195000  8.885000 177.395000 ;
        RECT  8.685000 177.595000  8.885000 177.795000 ;
        RECT  8.685000 177.995000  8.885000 178.195000 ;
        RECT  8.685000 178.395000  8.885000 178.595000 ;
        RECT  8.685000 178.795000  8.885000 178.995000 ;
        RECT  8.685000 179.195000  8.885000 179.395000 ;
        RECT  8.685000 179.595000  8.885000 179.795000 ;
        RECT  8.685000 179.995000  8.885000 180.195000 ;
        RECT  8.685000 180.395000  8.885000 180.595000 ;
        RECT  8.685000 180.795000  8.885000 180.995000 ;
        RECT  8.685000 181.195000  8.885000 181.395000 ;
        RECT  8.685000 181.595000  8.885000 181.795000 ;
        RECT  8.685000 181.995000  8.885000 182.195000 ;
        RECT  8.685000 182.395000  8.885000 182.595000 ;
        RECT  8.685000 182.795000  8.885000 182.995000 ;
        RECT  8.685000 183.195000  8.885000 183.395000 ;
        RECT  8.685000 183.595000  8.885000 183.795000 ;
        RECT  8.685000 183.995000  8.885000 184.195000 ;
        RECT  8.685000 184.395000  8.885000 184.595000 ;
        RECT  8.685000 184.795000  8.885000 184.995000 ;
        RECT  8.685000 185.195000  8.885000 185.395000 ;
        RECT  8.685000 185.595000  8.885000 185.795000 ;
        RECT  8.685000 185.995000  8.885000 186.195000 ;
        RECT  8.685000 186.395000  8.885000 186.595000 ;
        RECT  8.685000 186.795000  8.885000 186.995000 ;
        RECT  8.685000 187.195000  8.885000 187.395000 ;
        RECT  8.685000 187.595000  8.885000 187.795000 ;
        RECT  8.685000 187.995000  8.885000 188.195000 ;
        RECT  8.685000 188.395000  8.885000 188.595000 ;
        RECT  8.685000 188.795000  8.885000 188.995000 ;
        RECT  8.685000 189.195000  8.885000 189.395000 ;
        RECT  8.685000 189.595000  8.885000 189.795000 ;
        RECT  8.685000 189.995000  8.885000 190.195000 ;
        RECT  8.685000 190.395000  8.885000 190.595000 ;
        RECT  8.685000 190.795000  8.885000 190.995000 ;
        RECT  8.685000 191.195000  8.885000 191.395000 ;
        RECT  8.685000 191.595000  8.885000 191.795000 ;
        RECT  8.685000 191.995000  8.885000 192.195000 ;
        RECT  8.685000 192.395000  8.885000 192.595000 ;
        RECT  8.685000 192.795000  8.885000 192.995000 ;
        RECT  8.685000 193.195000  8.885000 193.395000 ;
        RECT  8.685000 193.595000  8.885000 193.795000 ;
        RECT  8.685000 193.995000  8.885000 194.195000 ;
        RECT  8.685000 194.395000  8.885000 194.595000 ;
        RECT  8.685000 194.795000  8.885000 194.995000 ;
        RECT  8.685000 195.200000  8.885000 195.400000 ;
        RECT  8.685000 195.605000  8.885000 195.805000 ;
        RECT  8.685000 196.010000  8.885000 196.210000 ;
        RECT  8.685000 196.415000  8.885000 196.615000 ;
        RECT  8.685000 196.820000  8.885000 197.020000 ;
        RECT  8.685000 197.225000  8.885000 197.425000 ;
        RECT  8.685000 197.630000  8.885000 197.830000 ;
        RECT  8.685000 198.035000  8.885000 198.235000 ;
        RECT  8.685000 198.440000  8.885000 198.640000 ;
        RECT  8.685000 198.845000  8.885000 199.045000 ;
        RECT  8.685000 199.250000  8.885000 199.450000 ;
        RECT  8.685000 199.655000  8.885000 199.855000 ;
        RECT  8.715000  25.910000  8.915000  26.110000 ;
        RECT  8.715000  26.340000  8.915000  26.540000 ;
        RECT  8.715000  26.770000  8.915000  26.970000 ;
        RECT  8.715000  27.200000  8.915000  27.400000 ;
        RECT  8.715000  27.630000  8.915000  27.830000 ;
        RECT  8.715000  28.060000  8.915000  28.260000 ;
        RECT  8.715000  28.490000  8.915000  28.690000 ;
        RECT  8.715000  28.920000  8.915000  29.120000 ;
        RECT  8.715000  29.350000  8.915000  29.550000 ;
        RECT  8.715000  29.780000  8.915000  29.980000 ;
        RECT  8.715000  30.210000  8.915000  30.410000 ;
        RECT  9.085000 175.995000  9.285000 176.195000 ;
        RECT  9.085000 176.395000  9.285000 176.595000 ;
        RECT  9.085000 176.795000  9.285000 176.995000 ;
        RECT  9.085000 177.195000  9.285000 177.395000 ;
        RECT  9.085000 177.595000  9.285000 177.795000 ;
        RECT  9.085000 177.995000  9.285000 178.195000 ;
        RECT  9.085000 178.395000  9.285000 178.595000 ;
        RECT  9.085000 178.795000  9.285000 178.995000 ;
        RECT  9.085000 179.195000  9.285000 179.395000 ;
        RECT  9.085000 179.595000  9.285000 179.795000 ;
        RECT  9.085000 179.995000  9.285000 180.195000 ;
        RECT  9.085000 180.395000  9.285000 180.595000 ;
        RECT  9.085000 180.795000  9.285000 180.995000 ;
        RECT  9.085000 181.195000  9.285000 181.395000 ;
        RECT  9.085000 181.595000  9.285000 181.795000 ;
        RECT  9.085000 181.995000  9.285000 182.195000 ;
        RECT  9.085000 182.395000  9.285000 182.595000 ;
        RECT  9.085000 182.795000  9.285000 182.995000 ;
        RECT  9.085000 183.195000  9.285000 183.395000 ;
        RECT  9.085000 183.595000  9.285000 183.795000 ;
        RECT  9.085000 183.995000  9.285000 184.195000 ;
        RECT  9.085000 184.395000  9.285000 184.595000 ;
        RECT  9.085000 184.795000  9.285000 184.995000 ;
        RECT  9.085000 185.195000  9.285000 185.395000 ;
        RECT  9.085000 185.595000  9.285000 185.795000 ;
        RECT  9.085000 185.995000  9.285000 186.195000 ;
        RECT  9.085000 186.395000  9.285000 186.595000 ;
        RECT  9.085000 186.795000  9.285000 186.995000 ;
        RECT  9.085000 187.195000  9.285000 187.395000 ;
        RECT  9.085000 187.595000  9.285000 187.795000 ;
        RECT  9.085000 187.995000  9.285000 188.195000 ;
        RECT  9.085000 188.395000  9.285000 188.595000 ;
        RECT  9.085000 188.795000  9.285000 188.995000 ;
        RECT  9.085000 189.195000  9.285000 189.395000 ;
        RECT  9.085000 189.595000  9.285000 189.795000 ;
        RECT  9.085000 189.995000  9.285000 190.195000 ;
        RECT  9.085000 190.395000  9.285000 190.595000 ;
        RECT  9.085000 190.795000  9.285000 190.995000 ;
        RECT  9.085000 191.195000  9.285000 191.395000 ;
        RECT  9.085000 191.595000  9.285000 191.795000 ;
        RECT  9.085000 191.995000  9.285000 192.195000 ;
        RECT  9.085000 192.395000  9.285000 192.595000 ;
        RECT  9.085000 192.795000  9.285000 192.995000 ;
        RECT  9.085000 193.195000  9.285000 193.395000 ;
        RECT  9.085000 193.595000  9.285000 193.795000 ;
        RECT  9.085000 193.995000  9.285000 194.195000 ;
        RECT  9.085000 194.395000  9.285000 194.595000 ;
        RECT  9.085000 194.795000  9.285000 194.995000 ;
        RECT  9.085000 195.200000  9.285000 195.400000 ;
        RECT  9.085000 195.605000  9.285000 195.805000 ;
        RECT  9.085000 196.010000  9.285000 196.210000 ;
        RECT  9.085000 196.415000  9.285000 196.615000 ;
        RECT  9.085000 196.820000  9.285000 197.020000 ;
        RECT  9.085000 197.225000  9.285000 197.425000 ;
        RECT  9.085000 197.630000  9.285000 197.830000 ;
        RECT  9.085000 198.035000  9.285000 198.235000 ;
        RECT  9.085000 198.440000  9.285000 198.640000 ;
        RECT  9.085000 198.845000  9.285000 199.045000 ;
        RECT  9.085000 199.250000  9.285000 199.450000 ;
        RECT  9.085000 199.655000  9.285000 199.855000 ;
        RECT  9.120000  25.910000  9.320000  26.110000 ;
        RECT  9.120000  26.340000  9.320000  26.540000 ;
        RECT  9.120000  26.770000  9.320000  26.970000 ;
        RECT  9.120000  27.200000  9.320000  27.400000 ;
        RECT  9.120000  27.630000  9.320000  27.830000 ;
        RECT  9.120000  28.060000  9.320000  28.260000 ;
        RECT  9.120000  28.490000  9.320000  28.690000 ;
        RECT  9.120000  28.920000  9.320000  29.120000 ;
        RECT  9.120000  29.350000  9.320000  29.550000 ;
        RECT  9.120000  29.780000  9.320000  29.980000 ;
        RECT  9.120000  30.210000  9.320000  30.410000 ;
        RECT  9.485000 175.995000  9.685000 176.195000 ;
        RECT  9.485000 176.395000  9.685000 176.595000 ;
        RECT  9.485000 176.795000  9.685000 176.995000 ;
        RECT  9.485000 177.195000  9.685000 177.395000 ;
        RECT  9.485000 177.595000  9.685000 177.795000 ;
        RECT  9.485000 177.995000  9.685000 178.195000 ;
        RECT  9.485000 178.395000  9.685000 178.595000 ;
        RECT  9.485000 178.795000  9.685000 178.995000 ;
        RECT  9.485000 179.195000  9.685000 179.395000 ;
        RECT  9.485000 179.595000  9.685000 179.795000 ;
        RECT  9.485000 179.995000  9.685000 180.195000 ;
        RECT  9.485000 180.395000  9.685000 180.595000 ;
        RECT  9.485000 180.795000  9.685000 180.995000 ;
        RECT  9.485000 181.195000  9.685000 181.395000 ;
        RECT  9.485000 181.595000  9.685000 181.795000 ;
        RECT  9.485000 181.995000  9.685000 182.195000 ;
        RECT  9.485000 182.395000  9.685000 182.595000 ;
        RECT  9.485000 182.795000  9.685000 182.995000 ;
        RECT  9.485000 183.195000  9.685000 183.395000 ;
        RECT  9.485000 183.595000  9.685000 183.795000 ;
        RECT  9.485000 183.995000  9.685000 184.195000 ;
        RECT  9.485000 184.395000  9.685000 184.595000 ;
        RECT  9.485000 184.795000  9.685000 184.995000 ;
        RECT  9.485000 185.195000  9.685000 185.395000 ;
        RECT  9.485000 185.595000  9.685000 185.795000 ;
        RECT  9.485000 185.995000  9.685000 186.195000 ;
        RECT  9.485000 186.395000  9.685000 186.595000 ;
        RECT  9.485000 186.795000  9.685000 186.995000 ;
        RECT  9.485000 187.195000  9.685000 187.395000 ;
        RECT  9.485000 187.595000  9.685000 187.795000 ;
        RECT  9.485000 187.995000  9.685000 188.195000 ;
        RECT  9.485000 188.395000  9.685000 188.595000 ;
        RECT  9.485000 188.795000  9.685000 188.995000 ;
        RECT  9.485000 189.195000  9.685000 189.395000 ;
        RECT  9.485000 189.595000  9.685000 189.795000 ;
        RECT  9.485000 189.995000  9.685000 190.195000 ;
        RECT  9.485000 190.395000  9.685000 190.595000 ;
        RECT  9.485000 190.795000  9.685000 190.995000 ;
        RECT  9.485000 191.195000  9.685000 191.395000 ;
        RECT  9.485000 191.595000  9.685000 191.795000 ;
        RECT  9.485000 191.995000  9.685000 192.195000 ;
        RECT  9.485000 192.395000  9.685000 192.595000 ;
        RECT  9.485000 192.795000  9.685000 192.995000 ;
        RECT  9.485000 193.195000  9.685000 193.395000 ;
        RECT  9.485000 193.595000  9.685000 193.795000 ;
        RECT  9.485000 193.995000  9.685000 194.195000 ;
        RECT  9.485000 194.395000  9.685000 194.595000 ;
        RECT  9.485000 194.795000  9.685000 194.995000 ;
        RECT  9.485000 195.200000  9.685000 195.400000 ;
        RECT  9.485000 195.605000  9.685000 195.805000 ;
        RECT  9.485000 196.010000  9.685000 196.210000 ;
        RECT  9.485000 196.415000  9.685000 196.615000 ;
        RECT  9.485000 196.820000  9.685000 197.020000 ;
        RECT  9.485000 197.225000  9.685000 197.425000 ;
        RECT  9.485000 197.630000  9.685000 197.830000 ;
        RECT  9.485000 198.035000  9.685000 198.235000 ;
        RECT  9.485000 198.440000  9.685000 198.640000 ;
        RECT  9.485000 198.845000  9.685000 199.045000 ;
        RECT  9.485000 199.250000  9.685000 199.450000 ;
        RECT  9.485000 199.655000  9.685000 199.855000 ;
        RECT  9.525000  25.910000  9.725000  26.110000 ;
        RECT  9.525000  26.340000  9.725000  26.540000 ;
        RECT  9.525000  26.770000  9.725000  26.970000 ;
        RECT  9.525000  27.200000  9.725000  27.400000 ;
        RECT  9.525000  27.630000  9.725000  27.830000 ;
        RECT  9.525000  28.060000  9.725000  28.260000 ;
        RECT  9.525000  28.490000  9.725000  28.690000 ;
        RECT  9.525000  28.920000  9.725000  29.120000 ;
        RECT  9.525000  29.350000  9.725000  29.550000 ;
        RECT  9.525000  29.780000  9.725000  29.980000 ;
        RECT  9.525000  30.210000  9.725000  30.410000 ;
        RECT  9.885000 175.995000 10.085000 176.195000 ;
        RECT  9.885000 176.395000 10.085000 176.595000 ;
        RECT  9.885000 176.795000 10.085000 176.995000 ;
        RECT  9.885000 177.195000 10.085000 177.395000 ;
        RECT  9.885000 177.595000 10.085000 177.795000 ;
        RECT  9.885000 177.995000 10.085000 178.195000 ;
        RECT  9.885000 178.395000 10.085000 178.595000 ;
        RECT  9.885000 178.795000 10.085000 178.995000 ;
        RECT  9.885000 179.195000 10.085000 179.395000 ;
        RECT  9.885000 179.595000 10.085000 179.795000 ;
        RECT  9.885000 179.995000 10.085000 180.195000 ;
        RECT  9.885000 180.395000 10.085000 180.595000 ;
        RECT  9.885000 180.795000 10.085000 180.995000 ;
        RECT  9.885000 181.195000 10.085000 181.395000 ;
        RECT  9.885000 181.595000 10.085000 181.795000 ;
        RECT  9.885000 181.995000 10.085000 182.195000 ;
        RECT  9.885000 182.395000 10.085000 182.595000 ;
        RECT  9.885000 182.795000 10.085000 182.995000 ;
        RECT  9.885000 183.195000 10.085000 183.395000 ;
        RECT  9.885000 183.595000 10.085000 183.795000 ;
        RECT  9.885000 183.995000 10.085000 184.195000 ;
        RECT  9.885000 184.395000 10.085000 184.595000 ;
        RECT  9.885000 184.795000 10.085000 184.995000 ;
        RECT  9.885000 185.195000 10.085000 185.395000 ;
        RECT  9.885000 185.595000 10.085000 185.795000 ;
        RECT  9.885000 185.995000 10.085000 186.195000 ;
        RECT  9.885000 186.395000 10.085000 186.595000 ;
        RECT  9.885000 186.795000 10.085000 186.995000 ;
        RECT  9.885000 187.195000 10.085000 187.395000 ;
        RECT  9.885000 187.595000 10.085000 187.795000 ;
        RECT  9.885000 187.995000 10.085000 188.195000 ;
        RECT  9.885000 188.395000 10.085000 188.595000 ;
        RECT  9.885000 188.795000 10.085000 188.995000 ;
        RECT  9.885000 189.195000 10.085000 189.395000 ;
        RECT  9.885000 189.595000 10.085000 189.795000 ;
        RECT  9.885000 189.995000 10.085000 190.195000 ;
        RECT  9.885000 190.395000 10.085000 190.595000 ;
        RECT  9.885000 190.795000 10.085000 190.995000 ;
        RECT  9.885000 191.195000 10.085000 191.395000 ;
        RECT  9.885000 191.595000 10.085000 191.795000 ;
        RECT  9.885000 191.995000 10.085000 192.195000 ;
        RECT  9.885000 192.395000 10.085000 192.595000 ;
        RECT  9.885000 192.795000 10.085000 192.995000 ;
        RECT  9.885000 193.195000 10.085000 193.395000 ;
        RECT  9.885000 193.595000 10.085000 193.795000 ;
        RECT  9.885000 193.995000 10.085000 194.195000 ;
        RECT  9.885000 194.395000 10.085000 194.595000 ;
        RECT  9.885000 194.795000 10.085000 194.995000 ;
        RECT  9.885000 195.200000 10.085000 195.400000 ;
        RECT  9.885000 195.605000 10.085000 195.805000 ;
        RECT  9.885000 196.010000 10.085000 196.210000 ;
        RECT  9.885000 196.415000 10.085000 196.615000 ;
        RECT  9.885000 196.820000 10.085000 197.020000 ;
        RECT  9.885000 197.225000 10.085000 197.425000 ;
        RECT  9.885000 197.630000 10.085000 197.830000 ;
        RECT  9.885000 198.035000 10.085000 198.235000 ;
        RECT  9.885000 198.440000 10.085000 198.640000 ;
        RECT  9.885000 198.845000 10.085000 199.045000 ;
        RECT  9.885000 199.250000 10.085000 199.450000 ;
        RECT  9.885000 199.655000 10.085000 199.855000 ;
        RECT  9.930000  25.910000 10.130000  26.110000 ;
        RECT  9.930000  26.340000 10.130000  26.540000 ;
        RECT  9.930000  26.770000 10.130000  26.970000 ;
        RECT  9.930000  27.200000 10.130000  27.400000 ;
        RECT  9.930000  27.630000 10.130000  27.830000 ;
        RECT  9.930000  28.060000 10.130000  28.260000 ;
        RECT  9.930000  28.490000 10.130000  28.690000 ;
        RECT  9.930000  28.920000 10.130000  29.120000 ;
        RECT  9.930000  29.350000 10.130000  29.550000 ;
        RECT  9.930000  29.780000 10.130000  29.980000 ;
        RECT  9.930000  30.210000 10.130000  30.410000 ;
        RECT 10.285000 175.995000 10.485000 176.195000 ;
        RECT 10.285000 176.395000 10.485000 176.595000 ;
        RECT 10.285000 176.795000 10.485000 176.995000 ;
        RECT 10.285000 177.195000 10.485000 177.395000 ;
        RECT 10.285000 177.595000 10.485000 177.795000 ;
        RECT 10.285000 177.995000 10.485000 178.195000 ;
        RECT 10.285000 178.395000 10.485000 178.595000 ;
        RECT 10.285000 178.795000 10.485000 178.995000 ;
        RECT 10.285000 179.195000 10.485000 179.395000 ;
        RECT 10.285000 179.595000 10.485000 179.795000 ;
        RECT 10.285000 179.995000 10.485000 180.195000 ;
        RECT 10.285000 180.395000 10.485000 180.595000 ;
        RECT 10.285000 180.795000 10.485000 180.995000 ;
        RECT 10.285000 181.195000 10.485000 181.395000 ;
        RECT 10.285000 181.595000 10.485000 181.795000 ;
        RECT 10.285000 181.995000 10.485000 182.195000 ;
        RECT 10.285000 182.395000 10.485000 182.595000 ;
        RECT 10.285000 182.795000 10.485000 182.995000 ;
        RECT 10.285000 183.195000 10.485000 183.395000 ;
        RECT 10.285000 183.595000 10.485000 183.795000 ;
        RECT 10.285000 183.995000 10.485000 184.195000 ;
        RECT 10.285000 184.395000 10.485000 184.595000 ;
        RECT 10.285000 184.795000 10.485000 184.995000 ;
        RECT 10.285000 185.195000 10.485000 185.395000 ;
        RECT 10.285000 185.595000 10.485000 185.795000 ;
        RECT 10.285000 185.995000 10.485000 186.195000 ;
        RECT 10.285000 186.395000 10.485000 186.595000 ;
        RECT 10.285000 186.795000 10.485000 186.995000 ;
        RECT 10.285000 187.195000 10.485000 187.395000 ;
        RECT 10.285000 187.595000 10.485000 187.795000 ;
        RECT 10.285000 187.995000 10.485000 188.195000 ;
        RECT 10.285000 188.395000 10.485000 188.595000 ;
        RECT 10.285000 188.795000 10.485000 188.995000 ;
        RECT 10.285000 189.195000 10.485000 189.395000 ;
        RECT 10.285000 189.595000 10.485000 189.795000 ;
        RECT 10.285000 189.995000 10.485000 190.195000 ;
        RECT 10.285000 190.395000 10.485000 190.595000 ;
        RECT 10.285000 190.795000 10.485000 190.995000 ;
        RECT 10.285000 191.195000 10.485000 191.395000 ;
        RECT 10.285000 191.595000 10.485000 191.795000 ;
        RECT 10.285000 191.995000 10.485000 192.195000 ;
        RECT 10.285000 192.395000 10.485000 192.595000 ;
        RECT 10.285000 192.795000 10.485000 192.995000 ;
        RECT 10.285000 193.195000 10.485000 193.395000 ;
        RECT 10.285000 193.595000 10.485000 193.795000 ;
        RECT 10.285000 193.995000 10.485000 194.195000 ;
        RECT 10.285000 194.395000 10.485000 194.595000 ;
        RECT 10.285000 194.795000 10.485000 194.995000 ;
        RECT 10.285000 195.200000 10.485000 195.400000 ;
        RECT 10.285000 195.605000 10.485000 195.805000 ;
        RECT 10.285000 196.010000 10.485000 196.210000 ;
        RECT 10.285000 196.415000 10.485000 196.615000 ;
        RECT 10.285000 196.820000 10.485000 197.020000 ;
        RECT 10.285000 197.225000 10.485000 197.425000 ;
        RECT 10.285000 197.630000 10.485000 197.830000 ;
        RECT 10.285000 198.035000 10.485000 198.235000 ;
        RECT 10.285000 198.440000 10.485000 198.640000 ;
        RECT 10.285000 198.845000 10.485000 199.045000 ;
        RECT 10.285000 199.250000 10.485000 199.450000 ;
        RECT 10.285000 199.655000 10.485000 199.855000 ;
        RECT 10.335000  25.910000 10.535000  26.110000 ;
        RECT 10.335000  26.340000 10.535000  26.540000 ;
        RECT 10.335000  26.770000 10.535000  26.970000 ;
        RECT 10.335000  27.200000 10.535000  27.400000 ;
        RECT 10.335000  27.630000 10.535000  27.830000 ;
        RECT 10.335000  28.060000 10.535000  28.260000 ;
        RECT 10.335000  28.490000 10.535000  28.690000 ;
        RECT 10.335000  28.920000 10.535000  29.120000 ;
        RECT 10.335000  29.350000 10.535000  29.550000 ;
        RECT 10.335000  29.780000 10.535000  29.980000 ;
        RECT 10.335000  30.210000 10.535000  30.410000 ;
        RECT 10.685000 175.995000 10.885000 176.195000 ;
        RECT 10.685000 176.395000 10.885000 176.595000 ;
        RECT 10.685000 176.795000 10.885000 176.995000 ;
        RECT 10.685000 177.195000 10.885000 177.395000 ;
        RECT 10.685000 177.595000 10.885000 177.795000 ;
        RECT 10.685000 177.995000 10.885000 178.195000 ;
        RECT 10.685000 178.395000 10.885000 178.595000 ;
        RECT 10.685000 178.795000 10.885000 178.995000 ;
        RECT 10.685000 179.195000 10.885000 179.395000 ;
        RECT 10.685000 179.595000 10.885000 179.795000 ;
        RECT 10.685000 179.995000 10.885000 180.195000 ;
        RECT 10.685000 180.395000 10.885000 180.595000 ;
        RECT 10.685000 180.795000 10.885000 180.995000 ;
        RECT 10.685000 181.195000 10.885000 181.395000 ;
        RECT 10.685000 181.595000 10.885000 181.795000 ;
        RECT 10.685000 181.995000 10.885000 182.195000 ;
        RECT 10.685000 182.395000 10.885000 182.595000 ;
        RECT 10.685000 182.795000 10.885000 182.995000 ;
        RECT 10.685000 183.195000 10.885000 183.395000 ;
        RECT 10.685000 183.595000 10.885000 183.795000 ;
        RECT 10.685000 183.995000 10.885000 184.195000 ;
        RECT 10.685000 184.395000 10.885000 184.595000 ;
        RECT 10.685000 184.795000 10.885000 184.995000 ;
        RECT 10.685000 185.195000 10.885000 185.395000 ;
        RECT 10.685000 185.595000 10.885000 185.795000 ;
        RECT 10.685000 185.995000 10.885000 186.195000 ;
        RECT 10.685000 186.395000 10.885000 186.595000 ;
        RECT 10.685000 186.795000 10.885000 186.995000 ;
        RECT 10.685000 187.195000 10.885000 187.395000 ;
        RECT 10.685000 187.595000 10.885000 187.795000 ;
        RECT 10.685000 187.995000 10.885000 188.195000 ;
        RECT 10.685000 188.395000 10.885000 188.595000 ;
        RECT 10.685000 188.795000 10.885000 188.995000 ;
        RECT 10.685000 189.195000 10.885000 189.395000 ;
        RECT 10.685000 189.595000 10.885000 189.795000 ;
        RECT 10.685000 189.995000 10.885000 190.195000 ;
        RECT 10.685000 190.395000 10.885000 190.595000 ;
        RECT 10.685000 190.795000 10.885000 190.995000 ;
        RECT 10.685000 191.195000 10.885000 191.395000 ;
        RECT 10.685000 191.595000 10.885000 191.795000 ;
        RECT 10.685000 191.995000 10.885000 192.195000 ;
        RECT 10.685000 192.395000 10.885000 192.595000 ;
        RECT 10.685000 192.795000 10.885000 192.995000 ;
        RECT 10.685000 193.195000 10.885000 193.395000 ;
        RECT 10.685000 193.595000 10.885000 193.795000 ;
        RECT 10.685000 193.995000 10.885000 194.195000 ;
        RECT 10.685000 194.395000 10.885000 194.595000 ;
        RECT 10.685000 194.795000 10.885000 194.995000 ;
        RECT 10.685000 195.200000 10.885000 195.400000 ;
        RECT 10.685000 195.605000 10.885000 195.805000 ;
        RECT 10.685000 196.010000 10.885000 196.210000 ;
        RECT 10.685000 196.415000 10.885000 196.615000 ;
        RECT 10.685000 196.820000 10.885000 197.020000 ;
        RECT 10.685000 197.225000 10.885000 197.425000 ;
        RECT 10.685000 197.630000 10.885000 197.830000 ;
        RECT 10.685000 198.035000 10.885000 198.235000 ;
        RECT 10.685000 198.440000 10.885000 198.640000 ;
        RECT 10.685000 198.845000 10.885000 199.045000 ;
        RECT 10.685000 199.250000 10.885000 199.450000 ;
        RECT 10.685000 199.655000 10.885000 199.855000 ;
        RECT 10.740000  25.910000 10.940000  26.110000 ;
        RECT 10.740000  26.340000 10.940000  26.540000 ;
        RECT 10.740000  26.770000 10.940000  26.970000 ;
        RECT 10.740000  27.200000 10.940000  27.400000 ;
        RECT 10.740000  27.630000 10.940000  27.830000 ;
        RECT 10.740000  28.060000 10.940000  28.260000 ;
        RECT 10.740000  28.490000 10.940000  28.690000 ;
        RECT 10.740000  28.920000 10.940000  29.120000 ;
        RECT 10.740000  29.350000 10.940000  29.550000 ;
        RECT 10.740000  29.780000 10.940000  29.980000 ;
        RECT 10.740000  30.210000 10.940000  30.410000 ;
        RECT 11.085000 175.995000 11.285000 176.195000 ;
        RECT 11.085000 176.395000 11.285000 176.595000 ;
        RECT 11.085000 176.795000 11.285000 176.995000 ;
        RECT 11.085000 177.195000 11.285000 177.395000 ;
        RECT 11.085000 177.595000 11.285000 177.795000 ;
        RECT 11.085000 177.995000 11.285000 178.195000 ;
        RECT 11.085000 178.395000 11.285000 178.595000 ;
        RECT 11.085000 178.795000 11.285000 178.995000 ;
        RECT 11.085000 179.195000 11.285000 179.395000 ;
        RECT 11.085000 179.595000 11.285000 179.795000 ;
        RECT 11.085000 179.995000 11.285000 180.195000 ;
        RECT 11.085000 180.395000 11.285000 180.595000 ;
        RECT 11.085000 180.795000 11.285000 180.995000 ;
        RECT 11.085000 181.195000 11.285000 181.395000 ;
        RECT 11.085000 181.595000 11.285000 181.795000 ;
        RECT 11.085000 181.995000 11.285000 182.195000 ;
        RECT 11.085000 182.395000 11.285000 182.595000 ;
        RECT 11.085000 182.795000 11.285000 182.995000 ;
        RECT 11.085000 183.195000 11.285000 183.395000 ;
        RECT 11.085000 183.595000 11.285000 183.795000 ;
        RECT 11.085000 183.995000 11.285000 184.195000 ;
        RECT 11.085000 184.395000 11.285000 184.595000 ;
        RECT 11.085000 184.795000 11.285000 184.995000 ;
        RECT 11.085000 185.195000 11.285000 185.395000 ;
        RECT 11.085000 185.595000 11.285000 185.795000 ;
        RECT 11.085000 185.995000 11.285000 186.195000 ;
        RECT 11.085000 186.395000 11.285000 186.595000 ;
        RECT 11.085000 186.795000 11.285000 186.995000 ;
        RECT 11.085000 187.195000 11.285000 187.395000 ;
        RECT 11.085000 187.595000 11.285000 187.795000 ;
        RECT 11.085000 187.995000 11.285000 188.195000 ;
        RECT 11.085000 188.395000 11.285000 188.595000 ;
        RECT 11.085000 188.795000 11.285000 188.995000 ;
        RECT 11.085000 189.195000 11.285000 189.395000 ;
        RECT 11.085000 189.595000 11.285000 189.795000 ;
        RECT 11.085000 189.995000 11.285000 190.195000 ;
        RECT 11.085000 190.395000 11.285000 190.595000 ;
        RECT 11.085000 190.795000 11.285000 190.995000 ;
        RECT 11.085000 191.195000 11.285000 191.395000 ;
        RECT 11.085000 191.595000 11.285000 191.795000 ;
        RECT 11.085000 191.995000 11.285000 192.195000 ;
        RECT 11.085000 192.395000 11.285000 192.595000 ;
        RECT 11.085000 192.795000 11.285000 192.995000 ;
        RECT 11.085000 193.195000 11.285000 193.395000 ;
        RECT 11.085000 193.595000 11.285000 193.795000 ;
        RECT 11.085000 193.995000 11.285000 194.195000 ;
        RECT 11.085000 194.395000 11.285000 194.595000 ;
        RECT 11.085000 194.795000 11.285000 194.995000 ;
        RECT 11.085000 195.200000 11.285000 195.400000 ;
        RECT 11.085000 195.605000 11.285000 195.805000 ;
        RECT 11.085000 196.010000 11.285000 196.210000 ;
        RECT 11.085000 196.415000 11.285000 196.615000 ;
        RECT 11.085000 196.820000 11.285000 197.020000 ;
        RECT 11.085000 197.225000 11.285000 197.425000 ;
        RECT 11.085000 197.630000 11.285000 197.830000 ;
        RECT 11.085000 198.035000 11.285000 198.235000 ;
        RECT 11.085000 198.440000 11.285000 198.640000 ;
        RECT 11.085000 198.845000 11.285000 199.045000 ;
        RECT 11.085000 199.250000 11.285000 199.450000 ;
        RECT 11.085000 199.655000 11.285000 199.855000 ;
        RECT 11.145000  25.910000 11.345000  26.110000 ;
        RECT 11.145000  26.340000 11.345000  26.540000 ;
        RECT 11.145000  26.770000 11.345000  26.970000 ;
        RECT 11.145000  27.200000 11.345000  27.400000 ;
        RECT 11.145000  27.630000 11.345000  27.830000 ;
        RECT 11.145000  28.060000 11.345000  28.260000 ;
        RECT 11.145000  28.490000 11.345000  28.690000 ;
        RECT 11.145000  28.920000 11.345000  29.120000 ;
        RECT 11.145000  29.350000 11.345000  29.550000 ;
        RECT 11.145000  29.780000 11.345000  29.980000 ;
        RECT 11.145000  30.210000 11.345000  30.410000 ;
        RECT 11.485000 175.995000 11.685000 176.195000 ;
        RECT 11.485000 176.395000 11.685000 176.595000 ;
        RECT 11.485000 176.795000 11.685000 176.995000 ;
        RECT 11.485000 177.195000 11.685000 177.395000 ;
        RECT 11.485000 177.595000 11.685000 177.795000 ;
        RECT 11.485000 177.995000 11.685000 178.195000 ;
        RECT 11.485000 178.395000 11.685000 178.595000 ;
        RECT 11.485000 178.795000 11.685000 178.995000 ;
        RECT 11.485000 179.195000 11.685000 179.395000 ;
        RECT 11.485000 179.595000 11.685000 179.795000 ;
        RECT 11.485000 179.995000 11.685000 180.195000 ;
        RECT 11.485000 180.395000 11.685000 180.595000 ;
        RECT 11.485000 180.795000 11.685000 180.995000 ;
        RECT 11.485000 181.195000 11.685000 181.395000 ;
        RECT 11.485000 181.595000 11.685000 181.795000 ;
        RECT 11.485000 181.995000 11.685000 182.195000 ;
        RECT 11.485000 182.395000 11.685000 182.595000 ;
        RECT 11.485000 182.795000 11.685000 182.995000 ;
        RECT 11.485000 183.195000 11.685000 183.395000 ;
        RECT 11.485000 183.595000 11.685000 183.795000 ;
        RECT 11.485000 183.995000 11.685000 184.195000 ;
        RECT 11.485000 184.395000 11.685000 184.595000 ;
        RECT 11.485000 184.795000 11.685000 184.995000 ;
        RECT 11.485000 185.195000 11.685000 185.395000 ;
        RECT 11.485000 185.595000 11.685000 185.795000 ;
        RECT 11.485000 185.995000 11.685000 186.195000 ;
        RECT 11.485000 186.395000 11.685000 186.595000 ;
        RECT 11.485000 186.795000 11.685000 186.995000 ;
        RECT 11.485000 187.195000 11.685000 187.395000 ;
        RECT 11.485000 187.595000 11.685000 187.795000 ;
        RECT 11.485000 187.995000 11.685000 188.195000 ;
        RECT 11.485000 188.395000 11.685000 188.595000 ;
        RECT 11.485000 188.795000 11.685000 188.995000 ;
        RECT 11.485000 189.195000 11.685000 189.395000 ;
        RECT 11.485000 189.595000 11.685000 189.795000 ;
        RECT 11.485000 189.995000 11.685000 190.195000 ;
        RECT 11.485000 190.395000 11.685000 190.595000 ;
        RECT 11.485000 190.795000 11.685000 190.995000 ;
        RECT 11.485000 191.195000 11.685000 191.395000 ;
        RECT 11.485000 191.595000 11.685000 191.795000 ;
        RECT 11.485000 191.995000 11.685000 192.195000 ;
        RECT 11.485000 192.395000 11.685000 192.595000 ;
        RECT 11.485000 192.795000 11.685000 192.995000 ;
        RECT 11.485000 193.195000 11.685000 193.395000 ;
        RECT 11.485000 193.595000 11.685000 193.795000 ;
        RECT 11.485000 193.995000 11.685000 194.195000 ;
        RECT 11.485000 194.395000 11.685000 194.595000 ;
        RECT 11.485000 194.795000 11.685000 194.995000 ;
        RECT 11.485000 195.200000 11.685000 195.400000 ;
        RECT 11.485000 195.605000 11.685000 195.805000 ;
        RECT 11.485000 196.010000 11.685000 196.210000 ;
        RECT 11.485000 196.415000 11.685000 196.615000 ;
        RECT 11.485000 196.820000 11.685000 197.020000 ;
        RECT 11.485000 197.225000 11.685000 197.425000 ;
        RECT 11.485000 197.630000 11.685000 197.830000 ;
        RECT 11.485000 198.035000 11.685000 198.235000 ;
        RECT 11.485000 198.440000 11.685000 198.640000 ;
        RECT 11.485000 198.845000 11.685000 199.045000 ;
        RECT 11.485000 199.250000 11.685000 199.450000 ;
        RECT 11.485000 199.655000 11.685000 199.855000 ;
        RECT 11.550000  25.910000 11.750000  26.110000 ;
        RECT 11.550000  26.340000 11.750000  26.540000 ;
        RECT 11.550000  26.770000 11.750000  26.970000 ;
        RECT 11.550000  27.200000 11.750000  27.400000 ;
        RECT 11.550000  27.630000 11.750000  27.830000 ;
        RECT 11.550000  28.060000 11.750000  28.260000 ;
        RECT 11.550000  28.490000 11.750000  28.690000 ;
        RECT 11.550000  28.920000 11.750000  29.120000 ;
        RECT 11.550000  29.350000 11.750000  29.550000 ;
        RECT 11.550000  29.780000 11.750000  29.980000 ;
        RECT 11.550000  30.210000 11.750000  30.410000 ;
        RECT 11.885000 175.995000 12.085000 176.195000 ;
        RECT 11.885000 176.395000 12.085000 176.595000 ;
        RECT 11.885000 176.795000 12.085000 176.995000 ;
        RECT 11.885000 177.195000 12.085000 177.395000 ;
        RECT 11.885000 177.595000 12.085000 177.795000 ;
        RECT 11.885000 177.995000 12.085000 178.195000 ;
        RECT 11.885000 178.395000 12.085000 178.595000 ;
        RECT 11.885000 178.795000 12.085000 178.995000 ;
        RECT 11.885000 179.195000 12.085000 179.395000 ;
        RECT 11.885000 179.595000 12.085000 179.795000 ;
        RECT 11.885000 179.995000 12.085000 180.195000 ;
        RECT 11.885000 180.395000 12.085000 180.595000 ;
        RECT 11.885000 180.795000 12.085000 180.995000 ;
        RECT 11.885000 181.195000 12.085000 181.395000 ;
        RECT 11.885000 181.595000 12.085000 181.795000 ;
        RECT 11.885000 181.995000 12.085000 182.195000 ;
        RECT 11.885000 182.395000 12.085000 182.595000 ;
        RECT 11.885000 182.795000 12.085000 182.995000 ;
        RECT 11.885000 183.195000 12.085000 183.395000 ;
        RECT 11.885000 183.595000 12.085000 183.795000 ;
        RECT 11.885000 183.995000 12.085000 184.195000 ;
        RECT 11.885000 184.395000 12.085000 184.595000 ;
        RECT 11.885000 184.795000 12.085000 184.995000 ;
        RECT 11.885000 185.195000 12.085000 185.395000 ;
        RECT 11.885000 185.595000 12.085000 185.795000 ;
        RECT 11.885000 185.995000 12.085000 186.195000 ;
        RECT 11.885000 186.395000 12.085000 186.595000 ;
        RECT 11.885000 186.795000 12.085000 186.995000 ;
        RECT 11.885000 187.195000 12.085000 187.395000 ;
        RECT 11.885000 187.595000 12.085000 187.795000 ;
        RECT 11.885000 187.995000 12.085000 188.195000 ;
        RECT 11.885000 188.395000 12.085000 188.595000 ;
        RECT 11.885000 188.795000 12.085000 188.995000 ;
        RECT 11.885000 189.195000 12.085000 189.395000 ;
        RECT 11.885000 189.595000 12.085000 189.795000 ;
        RECT 11.885000 189.995000 12.085000 190.195000 ;
        RECT 11.885000 190.395000 12.085000 190.595000 ;
        RECT 11.885000 190.795000 12.085000 190.995000 ;
        RECT 11.885000 191.195000 12.085000 191.395000 ;
        RECT 11.885000 191.595000 12.085000 191.795000 ;
        RECT 11.885000 191.995000 12.085000 192.195000 ;
        RECT 11.885000 192.395000 12.085000 192.595000 ;
        RECT 11.885000 192.795000 12.085000 192.995000 ;
        RECT 11.885000 193.195000 12.085000 193.395000 ;
        RECT 11.885000 193.595000 12.085000 193.795000 ;
        RECT 11.885000 193.995000 12.085000 194.195000 ;
        RECT 11.885000 194.395000 12.085000 194.595000 ;
        RECT 11.885000 194.795000 12.085000 194.995000 ;
        RECT 11.885000 195.200000 12.085000 195.400000 ;
        RECT 11.885000 195.605000 12.085000 195.805000 ;
        RECT 11.885000 196.010000 12.085000 196.210000 ;
        RECT 11.885000 196.415000 12.085000 196.615000 ;
        RECT 11.885000 196.820000 12.085000 197.020000 ;
        RECT 11.885000 197.225000 12.085000 197.425000 ;
        RECT 11.885000 197.630000 12.085000 197.830000 ;
        RECT 11.885000 198.035000 12.085000 198.235000 ;
        RECT 11.885000 198.440000 12.085000 198.640000 ;
        RECT 11.885000 198.845000 12.085000 199.045000 ;
        RECT 11.885000 199.250000 12.085000 199.450000 ;
        RECT 11.885000 199.655000 12.085000 199.855000 ;
        RECT 11.955000  25.910000 12.155000  26.110000 ;
        RECT 11.955000  26.340000 12.155000  26.540000 ;
        RECT 11.955000  26.770000 12.155000  26.970000 ;
        RECT 11.955000  27.200000 12.155000  27.400000 ;
        RECT 11.955000  27.630000 12.155000  27.830000 ;
        RECT 11.955000  28.060000 12.155000  28.260000 ;
        RECT 11.955000  28.490000 12.155000  28.690000 ;
        RECT 11.955000  28.920000 12.155000  29.120000 ;
        RECT 11.955000  29.350000 12.155000  29.550000 ;
        RECT 11.955000  29.780000 12.155000  29.980000 ;
        RECT 11.955000  30.210000 12.155000  30.410000 ;
        RECT 12.285000 175.995000 12.485000 176.195000 ;
        RECT 12.285000 176.395000 12.485000 176.595000 ;
        RECT 12.285000 176.795000 12.485000 176.995000 ;
        RECT 12.285000 177.195000 12.485000 177.395000 ;
        RECT 12.285000 177.595000 12.485000 177.795000 ;
        RECT 12.285000 177.995000 12.485000 178.195000 ;
        RECT 12.285000 178.395000 12.485000 178.595000 ;
        RECT 12.285000 178.795000 12.485000 178.995000 ;
        RECT 12.285000 179.195000 12.485000 179.395000 ;
        RECT 12.285000 179.595000 12.485000 179.795000 ;
        RECT 12.285000 179.995000 12.485000 180.195000 ;
        RECT 12.285000 180.395000 12.485000 180.595000 ;
        RECT 12.285000 180.795000 12.485000 180.995000 ;
        RECT 12.285000 181.195000 12.485000 181.395000 ;
        RECT 12.285000 181.595000 12.485000 181.795000 ;
        RECT 12.285000 181.995000 12.485000 182.195000 ;
        RECT 12.285000 182.395000 12.485000 182.595000 ;
        RECT 12.285000 182.795000 12.485000 182.995000 ;
        RECT 12.285000 183.195000 12.485000 183.395000 ;
        RECT 12.285000 183.595000 12.485000 183.795000 ;
        RECT 12.285000 183.995000 12.485000 184.195000 ;
        RECT 12.285000 184.395000 12.485000 184.595000 ;
        RECT 12.285000 184.795000 12.485000 184.995000 ;
        RECT 12.285000 185.195000 12.485000 185.395000 ;
        RECT 12.285000 185.595000 12.485000 185.795000 ;
        RECT 12.285000 185.995000 12.485000 186.195000 ;
        RECT 12.285000 186.395000 12.485000 186.595000 ;
        RECT 12.285000 186.795000 12.485000 186.995000 ;
        RECT 12.285000 187.195000 12.485000 187.395000 ;
        RECT 12.285000 187.595000 12.485000 187.795000 ;
        RECT 12.285000 187.995000 12.485000 188.195000 ;
        RECT 12.285000 188.395000 12.485000 188.595000 ;
        RECT 12.285000 188.795000 12.485000 188.995000 ;
        RECT 12.285000 189.195000 12.485000 189.395000 ;
        RECT 12.285000 189.595000 12.485000 189.795000 ;
        RECT 12.285000 189.995000 12.485000 190.195000 ;
        RECT 12.285000 190.395000 12.485000 190.595000 ;
        RECT 12.285000 190.795000 12.485000 190.995000 ;
        RECT 12.285000 191.195000 12.485000 191.395000 ;
        RECT 12.285000 191.595000 12.485000 191.795000 ;
        RECT 12.285000 191.995000 12.485000 192.195000 ;
        RECT 12.285000 192.395000 12.485000 192.595000 ;
        RECT 12.285000 192.795000 12.485000 192.995000 ;
        RECT 12.285000 193.195000 12.485000 193.395000 ;
        RECT 12.285000 193.595000 12.485000 193.795000 ;
        RECT 12.285000 193.995000 12.485000 194.195000 ;
        RECT 12.285000 194.395000 12.485000 194.595000 ;
        RECT 12.285000 194.795000 12.485000 194.995000 ;
        RECT 12.285000 195.200000 12.485000 195.400000 ;
        RECT 12.285000 195.605000 12.485000 195.805000 ;
        RECT 12.285000 196.010000 12.485000 196.210000 ;
        RECT 12.285000 196.415000 12.485000 196.615000 ;
        RECT 12.285000 196.820000 12.485000 197.020000 ;
        RECT 12.285000 197.225000 12.485000 197.425000 ;
        RECT 12.285000 197.630000 12.485000 197.830000 ;
        RECT 12.285000 198.035000 12.485000 198.235000 ;
        RECT 12.285000 198.440000 12.485000 198.640000 ;
        RECT 12.285000 198.845000 12.485000 199.045000 ;
        RECT 12.285000 199.250000 12.485000 199.450000 ;
        RECT 12.285000 199.655000 12.485000 199.855000 ;
        RECT 12.360000  25.910000 12.560000  26.110000 ;
        RECT 12.360000  26.340000 12.560000  26.540000 ;
        RECT 12.360000  26.770000 12.560000  26.970000 ;
        RECT 12.360000  27.200000 12.560000  27.400000 ;
        RECT 12.360000  27.630000 12.560000  27.830000 ;
        RECT 12.360000  28.060000 12.560000  28.260000 ;
        RECT 12.360000  28.490000 12.560000  28.690000 ;
        RECT 12.360000  28.920000 12.560000  29.120000 ;
        RECT 12.360000  29.350000 12.560000  29.550000 ;
        RECT 12.360000  29.780000 12.560000  29.980000 ;
        RECT 12.360000  30.210000 12.560000  30.410000 ;
        RECT 12.685000 175.995000 12.885000 176.195000 ;
        RECT 12.685000 176.395000 12.885000 176.595000 ;
        RECT 12.685000 176.795000 12.885000 176.995000 ;
        RECT 12.685000 177.195000 12.885000 177.395000 ;
        RECT 12.685000 177.595000 12.885000 177.795000 ;
        RECT 12.685000 177.995000 12.885000 178.195000 ;
        RECT 12.685000 178.395000 12.885000 178.595000 ;
        RECT 12.685000 178.795000 12.885000 178.995000 ;
        RECT 12.685000 179.195000 12.885000 179.395000 ;
        RECT 12.685000 179.595000 12.885000 179.795000 ;
        RECT 12.685000 179.995000 12.885000 180.195000 ;
        RECT 12.685000 180.395000 12.885000 180.595000 ;
        RECT 12.685000 180.795000 12.885000 180.995000 ;
        RECT 12.685000 181.195000 12.885000 181.395000 ;
        RECT 12.685000 181.595000 12.885000 181.795000 ;
        RECT 12.685000 181.995000 12.885000 182.195000 ;
        RECT 12.685000 182.395000 12.885000 182.595000 ;
        RECT 12.685000 182.795000 12.885000 182.995000 ;
        RECT 12.685000 183.195000 12.885000 183.395000 ;
        RECT 12.685000 183.595000 12.885000 183.795000 ;
        RECT 12.685000 183.995000 12.885000 184.195000 ;
        RECT 12.685000 184.395000 12.885000 184.595000 ;
        RECT 12.685000 184.795000 12.885000 184.995000 ;
        RECT 12.685000 185.195000 12.885000 185.395000 ;
        RECT 12.685000 185.595000 12.885000 185.795000 ;
        RECT 12.685000 185.995000 12.885000 186.195000 ;
        RECT 12.685000 186.395000 12.885000 186.595000 ;
        RECT 12.685000 186.795000 12.885000 186.995000 ;
        RECT 12.685000 187.195000 12.885000 187.395000 ;
        RECT 12.685000 187.595000 12.885000 187.795000 ;
        RECT 12.685000 187.995000 12.885000 188.195000 ;
        RECT 12.685000 188.395000 12.885000 188.595000 ;
        RECT 12.685000 188.795000 12.885000 188.995000 ;
        RECT 12.685000 189.195000 12.885000 189.395000 ;
        RECT 12.685000 189.595000 12.885000 189.795000 ;
        RECT 12.685000 189.995000 12.885000 190.195000 ;
        RECT 12.685000 190.395000 12.885000 190.595000 ;
        RECT 12.685000 190.795000 12.885000 190.995000 ;
        RECT 12.685000 191.195000 12.885000 191.395000 ;
        RECT 12.685000 191.595000 12.885000 191.795000 ;
        RECT 12.685000 191.995000 12.885000 192.195000 ;
        RECT 12.685000 192.395000 12.885000 192.595000 ;
        RECT 12.685000 192.795000 12.885000 192.995000 ;
        RECT 12.685000 193.195000 12.885000 193.395000 ;
        RECT 12.685000 193.595000 12.885000 193.795000 ;
        RECT 12.685000 193.995000 12.885000 194.195000 ;
        RECT 12.685000 194.395000 12.885000 194.595000 ;
        RECT 12.685000 194.795000 12.885000 194.995000 ;
        RECT 12.685000 195.200000 12.885000 195.400000 ;
        RECT 12.685000 195.605000 12.885000 195.805000 ;
        RECT 12.685000 196.010000 12.885000 196.210000 ;
        RECT 12.685000 196.415000 12.885000 196.615000 ;
        RECT 12.685000 196.820000 12.885000 197.020000 ;
        RECT 12.685000 197.225000 12.885000 197.425000 ;
        RECT 12.685000 197.630000 12.885000 197.830000 ;
        RECT 12.685000 198.035000 12.885000 198.235000 ;
        RECT 12.685000 198.440000 12.885000 198.640000 ;
        RECT 12.685000 198.845000 12.885000 199.045000 ;
        RECT 12.685000 199.250000 12.885000 199.450000 ;
        RECT 12.685000 199.655000 12.885000 199.855000 ;
        RECT 12.765000  25.910000 12.965000  26.110000 ;
        RECT 12.765000  26.340000 12.965000  26.540000 ;
        RECT 12.765000  26.770000 12.965000  26.970000 ;
        RECT 12.765000  27.200000 12.965000  27.400000 ;
        RECT 12.765000  27.630000 12.965000  27.830000 ;
        RECT 12.765000  28.060000 12.965000  28.260000 ;
        RECT 12.765000  28.490000 12.965000  28.690000 ;
        RECT 12.765000  28.920000 12.965000  29.120000 ;
        RECT 12.765000  29.350000 12.965000  29.550000 ;
        RECT 12.765000  29.780000 12.965000  29.980000 ;
        RECT 12.765000  30.210000 12.965000  30.410000 ;
        RECT 13.085000 175.995000 13.285000 176.195000 ;
        RECT 13.085000 176.395000 13.285000 176.595000 ;
        RECT 13.085000 176.795000 13.285000 176.995000 ;
        RECT 13.085000 177.195000 13.285000 177.395000 ;
        RECT 13.085000 177.595000 13.285000 177.795000 ;
        RECT 13.085000 177.995000 13.285000 178.195000 ;
        RECT 13.085000 178.395000 13.285000 178.595000 ;
        RECT 13.085000 178.795000 13.285000 178.995000 ;
        RECT 13.085000 179.195000 13.285000 179.395000 ;
        RECT 13.085000 179.595000 13.285000 179.795000 ;
        RECT 13.085000 179.995000 13.285000 180.195000 ;
        RECT 13.085000 180.395000 13.285000 180.595000 ;
        RECT 13.085000 180.795000 13.285000 180.995000 ;
        RECT 13.085000 181.195000 13.285000 181.395000 ;
        RECT 13.085000 181.595000 13.285000 181.795000 ;
        RECT 13.085000 181.995000 13.285000 182.195000 ;
        RECT 13.085000 182.395000 13.285000 182.595000 ;
        RECT 13.085000 182.795000 13.285000 182.995000 ;
        RECT 13.085000 183.195000 13.285000 183.395000 ;
        RECT 13.085000 183.595000 13.285000 183.795000 ;
        RECT 13.085000 183.995000 13.285000 184.195000 ;
        RECT 13.085000 184.395000 13.285000 184.595000 ;
        RECT 13.085000 184.795000 13.285000 184.995000 ;
        RECT 13.085000 185.195000 13.285000 185.395000 ;
        RECT 13.085000 185.595000 13.285000 185.795000 ;
        RECT 13.085000 185.995000 13.285000 186.195000 ;
        RECT 13.085000 186.395000 13.285000 186.595000 ;
        RECT 13.085000 186.795000 13.285000 186.995000 ;
        RECT 13.085000 187.195000 13.285000 187.395000 ;
        RECT 13.085000 187.595000 13.285000 187.795000 ;
        RECT 13.085000 187.995000 13.285000 188.195000 ;
        RECT 13.085000 188.395000 13.285000 188.595000 ;
        RECT 13.085000 188.795000 13.285000 188.995000 ;
        RECT 13.085000 189.195000 13.285000 189.395000 ;
        RECT 13.085000 189.595000 13.285000 189.795000 ;
        RECT 13.085000 189.995000 13.285000 190.195000 ;
        RECT 13.085000 190.395000 13.285000 190.595000 ;
        RECT 13.085000 190.795000 13.285000 190.995000 ;
        RECT 13.085000 191.195000 13.285000 191.395000 ;
        RECT 13.085000 191.595000 13.285000 191.795000 ;
        RECT 13.085000 191.995000 13.285000 192.195000 ;
        RECT 13.085000 192.395000 13.285000 192.595000 ;
        RECT 13.085000 192.795000 13.285000 192.995000 ;
        RECT 13.085000 193.195000 13.285000 193.395000 ;
        RECT 13.085000 193.595000 13.285000 193.795000 ;
        RECT 13.085000 193.995000 13.285000 194.195000 ;
        RECT 13.085000 194.395000 13.285000 194.595000 ;
        RECT 13.085000 194.795000 13.285000 194.995000 ;
        RECT 13.085000 195.200000 13.285000 195.400000 ;
        RECT 13.085000 195.605000 13.285000 195.805000 ;
        RECT 13.085000 196.010000 13.285000 196.210000 ;
        RECT 13.085000 196.415000 13.285000 196.615000 ;
        RECT 13.085000 196.820000 13.285000 197.020000 ;
        RECT 13.085000 197.225000 13.285000 197.425000 ;
        RECT 13.085000 197.630000 13.285000 197.830000 ;
        RECT 13.085000 198.035000 13.285000 198.235000 ;
        RECT 13.085000 198.440000 13.285000 198.640000 ;
        RECT 13.085000 198.845000 13.285000 199.045000 ;
        RECT 13.085000 199.250000 13.285000 199.450000 ;
        RECT 13.085000 199.655000 13.285000 199.855000 ;
        RECT 13.170000  25.910000 13.370000  26.110000 ;
        RECT 13.170000  26.340000 13.370000  26.540000 ;
        RECT 13.170000  26.770000 13.370000  26.970000 ;
        RECT 13.170000  27.200000 13.370000  27.400000 ;
        RECT 13.170000  27.630000 13.370000  27.830000 ;
        RECT 13.170000  28.060000 13.370000  28.260000 ;
        RECT 13.170000  28.490000 13.370000  28.690000 ;
        RECT 13.170000  28.920000 13.370000  29.120000 ;
        RECT 13.170000  29.350000 13.370000  29.550000 ;
        RECT 13.170000  29.780000 13.370000  29.980000 ;
        RECT 13.170000  30.210000 13.370000  30.410000 ;
        RECT 13.575000  25.910000 13.775000  26.110000 ;
        RECT 13.575000  26.340000 13.775000  26.540000 ;
        RECT 13.575000  26.770000 13.775000  26.970000 ;
        RECT 13.575000  27.200000 13.775000  27.400000 ;
        RECT 13.575000  27.630000 13.775000  27.830000 ;
        RECT 13.575000  28.060000 13.775000  28.260000 ;
        RECT 13.575000  28.490000 13.775000  28.690000 ;
        RECT 13.575000  28.920000 13.775000  29.120000 ;
        RECT 13.575000  29.350000 13.775000  29.550000 ;
        RECT 13.575000  29.780000 13.775000  29.980000 ;
        RECT 13.575000  30.210000 13.775000  30.410000 ;
        RECT 13.695000 197.250000 13.895000 197.450000 ;
        RECT 13.695000 197.650000 13.895000 197.850000 ;
        RECT 13.695000 198.050000 13.895000 198.250000 ;
        RECT 13.695000 198.450000 13.895000 198.650000 ;
        RECT 13.695000 198.850000 13.895000 199.050000 ;
        RECT 13.695000 199.250000 13.895000 199.450000 ;
        RECT 13.695000 199.650000 13.895000 199.850000 ;
        RECT 13.825000 196.295000 14.025000 196.495000 ;
        RECT 13.825000 196.705000 14.025000 196.905000 ;
        RECT 13.980000  25.910000 14.180000  26.110000 ;
        RECT 13.980000  26.340000 14.180000  26.540000 ;
        RECT 13.980000  26.770000 14.180000  26.970000 ;
        RECT 13.980000  27.200000 14.180000  27.400000 ;
        RECT 13.980000  27.630000 14.180000  27.830000 ;
        RECT 13.980000  28.060000 14.180000  28.260000 ;
        RECT 13.980000  28.490000 14.180000  28.690000 ;
        RECT 13.980000  28.920000 14.180000  29.120000 ;
        RECT 13.980000  29.350000 14.180000  29.550000 ;
        RECT 13.980000  29.780000 14.180000  29.980000 ;
        RECT 13.980000  30.210000 14.180000  30.410000 ;
        RECT 14.100000 197.250000 14.300000 197.450000 ;
        RECT 14.100000 197.650000 14.300000 197.850000 ;
        RECT 14.100000 198.050000 14.300000 198.250000 ;
        RECT 14.100000 198.450000 14.300000 198.650000 ;
        RECT 14.100000 198.850000 14.300000 199.050000 ;
        RECT 14.100000 199.250000 14.300000 199.450000 ;
        RECT 14.100000 199.650000 14.300000 199.850000 ;
        RECT 14.385000  25.910000 14.585000  26.110000 ;
        RECT 14.385000  26.340000 14.585000  26.540000 ;
        RECT 14.385000  26.770000 14.585000  26.970000 ;
        RECT 14.385000  27.200000 14.585000  27.400000 ;
        RECT 14.385000  27.630000 14.585000  27.830000 ;
        RECT 14.385000  28.060000 14.585000  28.260000 ;
        RECT 14.385000  28.490000 14.585000  28.690000 ;
        RECT 14.385000  28.920000 14.585000  29.120000 ;
        RECT 14.385000  29.350000 14.585000  29.550000 ;
        RECT 14.385000  29.780000 14.585000  29.980000 ;
        RECT 14.385000  30.210000 14.585000  30.410000 ;
        RECT 14.505000 197.250000 14.705000 197.450000 ;
        RECT 14.505000 197.650000 14.705000 197.850000 ;
        RECT 14.505000 198.050000 14.705000 198.250000 ;
        RECT 14.505000 198.450000 14.705000 198.650000 ;
        RECT 14.505000 198.850000 14.705000 199.050000 ;
        RECT 14.505000 199.250000 14.705000 199.450000 ;
        RECT 14.505000 199.650000 14.705000 199.850000 ;
        RECT 14.790000  25.910000 14.990000  26.110000 ;
        RECT 14.790000  26.340000 14.990000  26.540000 ;
        RECT 14.790000  26.770000 14.990000  26.970000 ;
        RECT 14.790000  27.200000 14.990000  27.400000 ;
        RECT 14.790000  27.630000 14.990000  27.830000 ;
        RECT 14.790000  28.060000 14.990000  28.260000 ;
        RECT 14.790000  28.490000 14.990000  28.690000 ;
        RECT 14.790000  28.920000 14.990000  29.120000 ;
        RECT 14.790000  29.350000 14.990000  29.550000 ;
        RECT 14.790000  29.780000 14.990000  29.980000 ;
        RECT 14.790000  30.210000 14.990000  30.410000 ;
        RECT 14.910000 197.250000 15.110000 197.450000 ;
        RECT 14.910000 197.650000 15.110000 197.850000 ;
        RECT 14.910000 198.050000 15.110000 198.250000 ;
        RECT 14.910000 198.450000 15.110000 198.650000 ;
        RECT 14.910000 198.850000 15.110000 199.050000 ;
        RECT 14.910000 199.250000 15.110000 199.450000 ;
        RECT 14.910000 199.650000 15.110000 199.850000 ;
        RECT 15.195000  25.910000 15.395000  26.110000 ;
        RECT 15.195000  26.340000 15.395000  26.540000 ;
        RECT 15.195000  26.770000 15.395000  26.970000 ;
        RECT 15.195000  27.200000 15.395000  27.400000 ;
        RECT 15.195000  27.630000 15.395000  27.830000 ;
        RECT 15.195000  28.060000 15.395000  28.260000 ;
        RECT 15.195000  28.490000 15.395000  28.690000 ;
        RECT 15.195000  28.920000 15.395000  29.120000 ;
        RECT 15.195000  29.350000 15.395000  29.550000 ;
        RECT 15.195000  29.780000 15.395000  29.980000 ;
        RECT 15.195000  30.210000 15.395000  30.410000 ;
        RECT 15.315000 197.250000 15.515000 197.450000 ;
        RECT 15.315000 197.650000 15.515000 197.850000 ;
        RECT 15.315000 198.050000 15.515000 198.250000 ;
        RECT 15.315000 198.450000 15.515000 198.650000 ;
        RECT 15.315000 198.850000 15.515000 199.050000 ;
        RECT 15.315000 199.250000 15.515000 199.450000 ;
        RECT 15.315000 199.650000 15.515000 199.850000 ;
        RECT 15.600000  25.910000 15.800000  26.110000 ;
        RECT 15.600000  26.340000 15.800000  26.540000 ;
        RECT 15.600000  26.770000 15.800000  26.970000 ;
        RECT 15.600000  27.200000 15.800000  27.400000 ;
        RECT 15.600000  27.630000 15.800000  27.830000 ;
        RECT 15.600000  28.060000 15.800000  28.260000 ;
        RECT 15.600000  28.490000 15.800000  28.690000 ;
        RECT 15.600000  28.920000 15.800000  29.120000 ;
        RECT 15.600000  29.350000 15.800000  29.550000 ;
        RECT 15.600000  29.780000 15.800000  29.980000 ;
        RECT 15.600000  30.210000 15.800000  30.410000 ;
        RECT 15.720000 197.250000 15.920000 197.450000 ;
        RECT 15.720000 197.650000 15.920000 197.850000 ;
        RECT 15.720000 198.050000 15.920000 198.250000 ;
        RECT 15.720000 198.450000 15.920000 198.650000 ;
        RECT 15.720000 198.850000 15.920000 199.050000 ;
        RECT 15.720000 199.250000 15.920000 199.450000 ;
        RECT 15.720000 199.650000 15.920000 199.850000 ;
        RECT 16.005000  25.910000 16.205000  26.110000 ;
        RECT 16.005000  26.340000 16.205000  26.540000 ;
        RECT 16.005000  26.770000 16.205000  26.970000 ;
        RECT 16.005000  27.200000 16.205000  27.400000 ;
        RECT 16.005000  27.630000 16.205000  27.830000 ;
        RECT 16.005000  28.060000 16.205000  28.260000 ;
        RECT 16.005000  28.490000 16.205000  28.690000 ;
        RECT 16.005000  28.920000 16.205000  29.120000 ;
        RECT 16.005000  29.350000 16.205000  29.550000 ;
        RECT 16.005000  29.780000 16.205000  29.980000 ;
        RECT 16.005000  30.210000 16.205000  30.410000 ;
        RECT 16.125000 197.250000 16.325000 197.450000 ;
        RECT 16.125000 197.650000 16.325000 197.850000 ;
        RECT 16.125000 198.050000 16.325000 198.250000 ;
        RECT 16.125000 198.450000 16.325000 198.650000 ;
        RECT 16.125000 198.850000 16.325000 199.050000 ;
        RECT 16.125000 199.250000 16.325000 199.450000 ;
        RECT 16.125000 199.650000 16.325000 199.850000 ;
        RECT 16.410000  25.910000 16.610000  26.110000 ;
        RECT 16.410000  26.340000 16.610000  26.540000 ;
        RECT 16.410000  26.770000 16.610000  26.970000 ;
        RECT 16.410000  27.200000 16.610000  27.400000 ;
        RECT 16.410000  27.630000 16.610000  27.830000 ;
        RECT 16.410000  28.060000 16.610000  28.260000 ;
        RECT 16.410000  28.490000 16.610000  28.690000 ;
        RECT 16.410000  28.920000 16.610000  29.120000 ;
        RECT 16.410000  29.350000 16.610000  29.550000 ;
        RECT 16.410000  29.780000 16.610000  29.980000 ;
        RECT 16.410000  30.210000 16.610000  30.410000 ;
        RECT 16.530000 197.250000 16.730000 197.450000 ;
        RECT 16.530000 197.650000 16.730000 197.850000 ;
        RECT 16.530000 198.050000 16.730000 198.250000 ;
        RECT 16.530000 198.450000 16.730000 198.650000 ;
        RECT 16.530000 198.850000 16.730000 199.050000 ;
        RECT 16.530000 199.250000 16.730000 199.450000 ;
        RECT 16.530000 199.650000 16.730000 199.850000 ;
        RECT 16.815000  25.910000 17.015000  26.110000 ;
        RECT 16.815000  26.340000 17.015000  26.540000 ;
        RECT 16.815000  26.770000 17.015000  26.970000 ;
        RECT 16.815000  27.200000 17.015000  27.400000 ;
        RECT 16.815000  27.630000 17.015000  27.830000 ;
        RECT 16.815000  28.060000 17.015000  28.260000 ;
        RECT 16.815000  28.490000 17.015000  28.690000 ;
        RECT 16.815000  28.920000 17.015000  29.120000 ;
        RECT 16.815000  29.350000 17.015000  29.550000 ;
        RECT 16.815000  29.780000 17.015000  29.980000 ;
        RECT 16.815000  30.210000 17.015000  30.410000 ;
        RECT 16.935000 197.250000 17.135000 197.450000 ;
        RECT 16.935000 197.650000 17.135000 197.850000 ;
        RECT 16.935000 198.050000 17.135000 198.250000 ;
        RECT 16.935000 198.450000 17.135000 198.650000 ;
        RECT 16.935000 198.850000 17.135000 199.050000 ;
        RECT 16.935000 199.250000 17.135000 199.450000 ;
        RECT 16.935000 199.650000 17.135000 199.850000 ;
        RECT 17.220000  25.910000 17.420000  26.110000 ;
        RECT 17.220000  26.340000 17.420000  26.540000 ;
        RECT 17.220000  26.770000 17.420000  26.970000 ;
        RECT 17.220000  27.200000 17.420000  27.400000 ;
        RECT 17.220000  27.630000 17.420000  27.830000 ;
        RECT 17.220000  28.060000 17.420000  28.260000 ;
        RECT 17.220000  28.490000 17.420000  28.690000 ;
        RECT 17.220000  28.920000 17.420000  29.120000 ;
        RECT 17.220000  29.350000 17.420000  29.550000 ;
        RECT 17.220000  29.780000 17.420000  29.980000 ;
        RECT 17.220000  30.210000 17.420000  30.410000 ;
        RECT 17.340000 197.250000 17.540000 197.450000 ;
        RECT 17.340000 197.650000 17.540000 197.850000 ;
        RECT 17.340000 198.050000 17.540000 198.250000 ;
        RECT 17.340000 198.450000 17.540000 198.650000 ;
        RECT 17.340000 198.850000 17.540000 199.050000 ;
        RECT 17.340000 199.250000 17.540000 199.450000 ;
        RECT 17.340000 199.650000 17.540000 199.850000 ;
        RECT 17.625000  25.910000 17.825000  26.110000 ;
        RECT 17.625000  26.340000 17.825000  26.540000 ;
        RECT 17.625000  26.770000 17.825000  26.970000 ;
        RECT 17.625000  27.200000 17.825000  27.400000 ;
        RECT 17.625000  27.630000 17.825000  27.830000 ;
        RECT 17.625000  28.060000 17.825000  28.260000 ;
        RECT 17.625000  28.490000 17.825000  28.690000 ;
        RECT 17.625000  28.920000 17.825000  29.120000 ;
        RECT 17.625000  29.350000 17.825000  29.550000 ;
        RECT 17.625000  29.780000 17.825000  29.980000 ;
        RECT 17.625000  30.210000 17.825000  30.410000 ;
        RECT 17.745000 197.250000 17.945000 197.450000 ;
        RECT 17.745000 197.650000 17.945000 197.850000 ;
        RECT 17.745000 198.050000 17.945000 198.250000 ;
        RECT 17.745000 198.450000 17.945000 198.650000 ;
        RECT 17.745000 198.850000 17.945000 199.050000 ;
        RECT 17.745000 199.250000 17.945000 199.450000 ;
        RECT 17.745000 199.650000 17.945000 199.850000 ;
        RECT 18.030000  25.910000 18.230000  26.110000 ;
        RECT 18.030000  26.340000 18.230000  26.540000 ;
        RECT 18.030000  26.770000 18.230000  26.970000 ;
        RECT 18.030000  27.200000 18.230000  27.400000 ;
        RECT 18.030000  27.630000 18.230000  27.830000 ;
        RECT 18.030000  28.060000 18.230000  28.260000 ;
        RECT 18.030000  28.490000 18.230000  28.690000 ;
        RECT 18.030000  28.920000 18.230000  29.120000 ;
        RECT 18.030000  29.350000 18.230000  29.550000 ;
        RECT 18.030000  29.780000 18.230000  29.980000 ;
        RECT 18.030000  30.210000 18.230000  30.410000 ;
        RECT 18.150000 197.250000 18.350000 197.450000 ;
        RECT 18.150000 197.650000 18.350000 197.850000 ;
        RECT 18.150000 198.050000 18.350000 198.250000 ;
        RECT 18.150000 198.450000 18.350000 198.650000 ;
        RECT 18.150000 198.850000 18.350000 199.050000 ;
        RECT 18.150000 199.250000 18.350000 199.450000 ;
        RECT 18.150000 199.650000 18.350000 199.850000 ;
        RECT 18.435000  25.910000 18.635000  26.110000 ;
        RECT 18.435000  26.340000 18.635000  26.540000 ;
        RECT 18.435000  26.770000 18.635000  26.970000 ;
        RECT 18.435000  27.200000 18.635000  27.400000 ;
        RECT 18.435000  27.630000 18.635000  27.830000 ;
        RECT 18.435000  28.060000 18.635000  28.260000 ;
        RECT 18.435000  28.490000 18.635000  28.690000 ;
        RECT 18.435000  28.920000 18.635000  29.120000 ;
        RECT 18.435000  29.350000 18.635000  29.550000 ;
        RECT 18.435000  29.780000 18.635000  29.980000 ;
        RECT 18.435000  30.210000 18.635000  30.410000 ;
        RECT 18.555000 197.250000 18.755000 197.450000 ;
        RECT 18.555000 197.650000 18.755000 197.850000 ;
        RECT 18.555000 198.050000 18.755000 198.250000 ;
        RECT 18.555000 198.450000 18.755000 198.650000 ;
        RECT 18.555000 198.850000 18.755000 199.050000 ;
        RECT 18.555000 199.250000 18.755000 199.450000 ;
        RECT 18.555000 199.650000 18.755000 199.850000 ;
        RECT 18.840000  25.910000 19.040000  26.110000 ;
        RECT 18.840000  26.340000 19.040000  26.540000 ;
        RECT 18.840000  26.770000 19.040000  26.970000 ;
        RECT 18.840000  27.200000 19.040000  27.400000 ;
        RECT 18.840000  27.630000 19.040000  27.830000 ;
        RECT 18.840000  28.060000 19.040000  28.260000 ;
        RECT 18.840000  28.490000 19.040000  28.690000 ;
        RECT 18.840000  28.920000 19.040000  29.120000 ;
        RECT 18.840000  29.350000 19.040000  29.550000 ;
        RECT 18.840000  29.780000 19.040000  29.980000 ;
        RECT 18.840000  30.210000 19.040000  30.410000 ;
        RECT 18.960000 197.250000 19.160000 197.450000 ;
        RECT 18.960000 197.650000 19.160000 197.850000 ;
        RECT 18.960000 198.050000 19.160000 198.250000 ;
        RECT 18.960000 198.450000 19.160000 198.650000 ;
        RECT 18.960000 198.850000 19.160000 199.050000 ;
        RECT 18.960000 199.250000 19.160000 199.450000 ;
        RECT 18.960000 199.650000 19.160000 199.850000 ;
        RECT 19.245000  25.910000 19.445000  26.110000 ;
        RECT 19.245000  26.340000 19.445000  26.540000 ;
        RECT 19.245000  26.770000 19.445000  26.970000 ;
        RECT 19.245000  27.200000 19.445000  27.400000 ;
        RECT 19.245000  27.630000 19.445000  27.830000 ;
        RECT 19.245000  28.060000 19.445000  28.260000 ;
        RECT 19.245000  28.490000 19.445000  28.690000 ;
        RECT 19.245000  28.920000 19.445000  29.120000 ;
        RECT 19.245000  29.350000 19.445000  29.550000 ;
        RECT 19.245000  29.780000 19.445000  29.980000 ;
        RECT 19.245000  30.210000 19.445000  30.410000 ;
        RECT 19.365000 197.250000 19.565000 197.450000 ;
        RECT 19.365000 197.650000 19.565000 197.850000 ;
        RECT 19.365000 198.050000 19.565000 198.250000 ;
        RECT 19.365000 198.450000 19.565000 198.650000 ;
        RECT 19.365000 198.850000 19.565000 199.050000 ;
        RECT 19.365000 199.250000 19.565000 199.450000 ;
        RECT 19.365000 199.650000 19.565000 199.850000 ;
        RECT 19.650000  25.910000 19.850000  26.110000 ;
        RECT 19.650000  26.340000 19.850000  26.540000 ;
        RECT 19.650000  26.770000 19.850000  26.970000 ;
        RECT 19.650000  27.200000 19.850000  27.400000 ;
        RECT 19.650000  27.630000 19.850000  27.830000 ;
        RECT 19.650000  28.060000 19.850000  28.260000 ;
        RECT 19.650000  28.490000 19.850000  28.690000 ;
        RECT 19.650000  28.920000 19.850000  29.120000 ;
        RECT 19.650000  29.350000 19.850000  29.550000 ;
        RECT 19.650000  29.780000 19.850000  29.980000 ;
        RECT 19.650000  30.210000 19.850000  30.410000 ;
        RECT 19.770000 197.250000 19.970000 197.450000 ;
        RECT 19.770000 197.650000 19.970000 197.850000 ;
        RECT 19.770000 198.050000 19.970000 198.250000 ;
        RECT 19.770000 198.450000 19.970000 198.650000 ;
        RECT 19.770000 198.850000 19.970000 199.050000 ;
        RECT 19.770000 199.250000 19.970000 199.450000 ;
        RECT 19.770000 199.650000 19.970000 199.850000 ;
        RECT 20.055000  25.910000 20.255000  26.110000 ;
        RECT 20.055000  26.340000 20.255000  26.540000 ;
        RECT 20.055000  26.770000 20.255000  26.970000 ;
        RECT 20.055000  27.200000 20.255000  27.400000 ;
        RECT 20.055000  27.630000 20.255000  27.830000 ;
        RECT 20.055000  28.060000 20.255000  28.260000 ;
        RECT 20.055000  28.490000 20.255000  28.690000 ;
        RECT 20.055000  28.920000 20.255000  29.120000 ;
        RECT 20.055000  29.350000 20.255000  29.550000 ;
        RECT 20.055000  29.780000 20.255000  29.980000 ;
        RECT 20.055000  30.210000 20.255000  30.410000 ;
        RECT 20.175000 197.250000 20.375000 197.450000 ;
        RECT 20.175000 197.650000 20.375000 197.850000 ;
        RECT 20.175000 198.050000 20.375000 198.250000 ;
        RECT 20.175000 198.450000 20.375000 198.650000 ;
        RECT 20.175000 198.850000 20.375000 199.050000 ;
        RECT 20.175000 199.250000 20.375000 199.450000 ;
        RECT 20.175000 199.650000 20.375000 199.850000 ;
        RECT 20.460000  25.910000 20.660000  26.110000 ;
        RECT 20.460000  26.340000 20.660000  26.540000 ;
        RECT 20.460000  26.770000 20.660000  26.970000 ;
        RECT 20.460000  27.200000 20.660000  27.400000 ;
        RECT 20.460000  27.630000 20.660000  27.830000 ;
        RECT 20.460000  28.060000 20.660000  28.260000 ;
        RECT 20.460000  28.490000 20.660000  28.690000 ;
        RECT 20.460000  28.920000 20.660000  29.120000 ;
        RECT 20.460000  29.350000 20.660000  29.550000 ;
        RECT 20.460000  29.780000 20.660000  29.980000 ;
        RECT 20.460000  30.210000 20.660000  30.410000 ;
        RECT 20.580000 197.250000 20.780000 197.450000 ;
        RECT 20.580000 197.650000 20.780000 197.850000 ;
        RECT 20.580000 198.050000 20.780000 198.250000 ;
        RECT 20.580000 198.450000 20.780000 198.650000 ;
        RECT 20.580000 198.850000 20.780000 199.050000 ;
        RECT 20.580000 199.250000 20.780000 199.450000 ;
        RECT 20.580000 199.650000 20.780000 199.850000 ;
        RECT 20.865000  25.910000 21.065000  26.110000 ;
        RECT 20.865000  26.340000 21.065000  26.540000 ;
        RECT 20.865000  26.770000 21.065000  26.970000 ;
        RECT 20.865000  27.200000 21.065000  27.400000 ;
        RECT 20.865000  27.630000 21.065000  27.830000 ;
        RECT 20.865000  28.060000 21.065000  28.260000 ;
        RECT 20.865000  28.490000 21.065000  28.690000 ;
        RECT 20.865000  28.920000 21.065000  29.120000 ;
        RECT 20.865000  29.350000 21.065000  29.550000 ;
        RECT 20.865000  29.780000 21.065000  29.980000 ;
        RECT 20.865000  30.210000 21.065000  30.410000 ;
        RECT 20.985000 197.250000 21.185000 197.450000 ;
        RECT 20.985000 197.650000 21.185000 197.850000 ;
        RECT 20.985000 198.050000 21.185000 198.250000 ;
        RECT 20.985000 198.450000 21.185000 198.650000 ;
        RECT 20.985000 198.850000 21.185000 199.050000 ;
        RECT 20.985000 199.250000 21.185000 199.450000 ;
        RECT 20.985000 199.650000 21.185000 199.850000 ;
        RECT 21.270000  25.910000 21.470000  26.110000 ;
        RECT 21.270000  26.340000 21.470000  26.540000 ;
        RECT 21.270000  26.770000 21.470000  26.970000 ;
        RECT 21.270000  27.200000 21.470000  27.400000 ;
        RECT 21.270000  27.630000 21.470000  27.830000 ;
        RECT 21.270000  28.060000 21.470000  28.260000 ;
        RECT 21.270000  28.490000 21.470000  28.690000 ;
        RECT 21.270000  28.920000 21.470000  29.120000 ;
        RECT 21.270000  29.350000 21.470000  29.550000 ;
        RECT 21.270000  29.780000 21.470000  29.980000 ;
        RECT 21.270000  30.210000 21.470000  30.410000 ;
        RECT 21.390000 197.250000 21.590000 197.450000 ;
        RECT 21.390000 197.650000 21.590000 197.850000 ;
        RECT 21.390000 198.050000 21.590000 198.250000 ;
        RECT 21.390000 198.450000 21.590000 198.650000 ;
        RECT 21.390000 198.850000 21.590000 199.050000 ;
        RECT 21.390000 199.250000 21.590000 199.450000 ;
        RECT 21.390000 199.650000 21.590000 199.850000 ;
        RECT 21.675000  25.910000 21.875000  26.110000 ;
        RECT 21.675000  26.340000 21.875000  26.540000 ;
        RECT 21.675000  26.770000 21.875000  26.970000 ;
        RECT 21.675000  27.200000 21.875000  27.400000 ;
        RECT 21.675000  27.630000 21.875000  27.830000 ;
        RECT 21.675000  28.060000 21.875000  28.260000 ;
        RECT 21.675000  28.490000 21.875000  28.690000 ;
        RECT 21.675000  28.920000 21.875000  29.120000 ;
        RECT 21.675000  29.350000 21.875000  29.550000 ;
        RECT 21.675000  29.780000 21.875000  29.980000 ;
        RECT 21.675000  30.210000 21.875000  30.410000 ;
        RECT 21.795000 197.250000 21.995000 197.450000 ;
        RECT 21.795000 197.650000 21.995000 197.850000 ;
        RECT 21.795000 198.050000 21.995000 198.250000 ;
        RECT 21.795000 198.450000 21.995000 198.650000 ;
        RECT 21.795000 198.850000 21.995000 199.050000 ;
        RECT 21.795000 199.250000 21.995000 199.450000 ;
        RECT 21.795000 199.650000 21.995000 199.850000 ;
        RECT 22.080000  25.910000 22.280000  26.110000 ;
        RECT 22.080000  26.340000 22.280000  26.540000 ;
        RECT 22.080000  26.770000 22.280000  26.970000 ;
        RECT 22.080000  27.200000 22.280000  27.400000 ;
        RECT 22.080000  27.630000 22.280000  27.830000 ;
        RECT 22.080000  28.060000 22.280000  28.260000 ;
        RECT 22.080000  28.490000 22.280000  28.690000 ;
        RECT 22.080000  28.920000 22.280000  29.120000 ;
        RECT 22.080000  29.350000 22.280000  29.550000 ;
        RECT 22.080000  29.780000 22.280000  29.980000 ;
        RECT 22.080000  30.210000 22.280000  30.410000 ;
        RECT 22.200000 197.250000 22.400000 197.450000 ;
        RECT 22.200000 197.650000 22.400000 197.850000 ;
        RECT 22.200000 198.050000 22.400000 198.250000 ;
        RECT 22.200000 198.450000 22.400000 198.650000 ;
        RECT 22.200000 198.850000 22.400000 199.050000 ;
        RECT 22.200000 199.250000 22.400000 199.450000 ;
        RECT 22.200000 199.650000 22.400000 199.850000 ;
        RECT 22.485000  25.910000 22.685000  26.110000 ;
        RECT 22.485000  26.340000 22.685000  26.540000 ;
        RECT 22.485000  26.770000 22.685000  26.970000 ;
        RECT 22.485000  27.200000 22.685000  27.400000 ;
        RECT 22.485000  27.630000 22.685000  27.830000 ;
        RECT 22.485000  28.060000 22.685000  28.260000 ;
        RECT 22.485000  28.490000 22.685000  28.690000 ;
        RECT 22.485000  28.920000 22.685000  29.120000 ;
        RECT 22.485000  29.350000 22.685000  29.550000 ;
        RECT 22.485000  29.780000 22.685000  29.980000 ;
        RECT 22.485000  30.210000 22.685000  30.410000 ;
        RECT 22.605000 197.250000 22.805000 197.450000 ;
        RECT 22.605000 197.650000 22.805000 197.850000 ;
        RECT 22.605000 198.050000 22.805000 198.250000 ;
        RECT 22.605000 198.450000 22.805000 198.650000 ;
        RECT 22.605000 198.850000 22.805000 199.050000 ;
        RECT 22.605000 199.250000 22.805000 199.450000 ;
        RECT 22.605000 199.650000 22.805000 199.850000 ;
        RECT 22.890000  25.910000 23.090000  26.110000 ;
        RECT 22.890000  26.340000 23.090000  26.540000 ;
        RECT 22.890000  26.770000 23.090000  26.970000 ;
        RECT 22.890000  27.200000 23.090000  27.400000 ;
        RECT 22.890000  27.630000 23.090000  27.830000 ;
        RECT 22.890000  28.060000 23.090000  28.260000 ;
        RECT 22.890000  28.490000 23.090000  28.690000 ;
        RECT 22.890000  28.920000 23.090000  29.120000 ;
        RECT 22.890000  29.350000 23.090000  29.550000 ;
        RECT 22.890000  29.780000 23.090000  29.980000 ;
        RECT 22.890000  30.210000 23.090000  30.410000 ;
        RECT 23.010000 197.250000 23.210000 197.450000 ;
        RECT 23.010000 197.650000 23.210000 197.850000 ;
        RECT 23.010000 198.050000 23.210000 198.250000 ;
        RECT 23.010000 198.450000 23.210000 198.650000 ;
        RECT 23.010000 198.850000 23.210000 199.050000 ;
        RECT 23.010000 199.250000 23.210000 199.450000 ;
        RECT 23.010000 199.650000 23.210000 199.850000 ;
        RECT 23.295000  25.910000 23.495000  26.110000 ;
        RECT 23.295000  26.340000 23.495000  26.540000 ;
        RECT 23.295000  26.770000 23.495000  26.970000 ;
        RECT 23.295000  27.200000 23.495000  27.400000 ;
        RECT 23.295000  27.630000 23.495000  27.830000 ;
        RECT 23.295000  28.060000 23.495000  28.260000 ;
        RECT 23.295000  28.490000 23.495000  28.690000 ;
        RECT 23.295000  28.920000 23.495000  29.120000 ;
        RECT 23.295000  29.350000 23.495000  29.550000 ;
        RECT 23.295000  29.780000 23.495000  29.980000 ;
        RECT 23.295000  30.210000 23.495000  30.410000 ;
        RECT 23.415000 197.250000 23.615000 197.450000 ;
        RECT 23.415000 197.650000 23.615000 197.850000 ;
        RECT 23.415000 198.050000 23.615000 198.250000 ;
        RECT 23.415000 198.450000 23.615000 198.650000 ;
        RECT 23.415000 198.850000 23.615000 199.050000 ;
        RECT 23.415000 199.250000 23.615000 199.450000 ;
        RECT 23.415000 199.650000 23.615000 199.850000 ;
        RECT 23.700000  25.910000 23.900000  26.110000 ;
        RECT 23.700000  26.340000 23.900000  26.540000 ;
        RECT 23.700000  26.770000 23.900000  26.970000 ;
        RECT 23.700000  27.200000 23.900000  27.400000 ;
        RECT 23.700000  27.630000 23.900000  27.830000 ;
        RECT 23.700000  28.060000 23.900000  28.260000 ;
        RECT 23.700000  28.490000 23.900000  28.690000 ;
        RECT 23.700000  28.920000 23.900000  29.120000 ;
        RECT 23.700000  29.350000 23.900000  29.550000 ;
        RECT 23.700000  29.780000 23.900000  29.980000 ;
        RECT 23.700000  30.210000 23.900000  30.410000 ;
        RECT 23.820000 197.250000 24.020000 197.450000 ;
        RECT 23.820000 197.650000 24.020000 197.850000 ;
        RECT 23.820000 198.050000 24.020000 198.250000 ;
        RECT 23.820000 198.450000 24.020000 198.650000 ;
        RECT 23.820000 198.850000 24.020000 199.050000 ;
        RECT 23.820000 199.250000 24.020000 199.450000 ;
        RECT 23.820000 199.650000 24.020000 199.850000 ;
        RECT 24.105000  25.910000 24.305000  26.110000 ;
        RECT 24.105000  26.340000 24.305000  26.540000 ;
        RECT 24.105000  26.770000 24.305000  26.970000 ;
        RECT 24.105000  27.200000 24.305000  27.400000 ;
        RECT 24.105000  27.630000 24.305000  27.830000 ;
        RECT 24.105000  28.060000 24.305000  28.260000 ;
        RECT 24.105000  28.490000 24.305000  28.690000 ;
        RECT 24.105000  28.920000 24.305000  29.120000 ;
        RECT 24.105000  29.350000 24.305000  29.550000 ;
        RECT 24.105000  29.780000 24.305000  29.980000 ;
        RECT 24.105000  30.210000 24.305000  30.410000 ;
        RECT 24.225000 197.250000 24.425000 197.450000 ;
        RECT 24.225000 197.650000 24.425000 197.850000 ;
        RECT 24.225000 198.050000 24.425000 198.250000 ;
        RECT 24.225000 198.450000 24.425000 198.650000 ;
        RECT 24.225000 198.850000 24.425000 199.050000 ;
        RECT 24.225000 199.250000 24.425000 199.450000 ;
        RECT 24.225000 199.650000 24.425000 199.850000 ;
        RECT 24.630000 197.250000 24.830000 197.450000 ;
        RECT 24.630000 197.650000 24.830000 197.850000 ;
        RECT 24.630000 198.050000 24.830000 198.250000 ;
        RECT 24.630000 198.450000 24.830000 198.650000 ;
        RECT 24.630000 198.850000 24.830000 199.050000 ;
        RECT 24.630000 199.250000 24.830000 199.450000 ;
        RECT 24.630000 199.650000 24.830000 199.850000 ;
        RECT 25.035000 197.250000 25.235000 197.450000 ;
        RECT 25.035000 197.650000 25.235000 197.850000 ;
        RECT 25.035000 198.050000 25.235000 198.250000 ;
        RECT 25.035000 198.450000 25.235000 198.650000 ;
        RECT 25.035000 198.850000 25.235000 199.050000 ;
        RECT 25.035000 199.250000 25.235000 199.450000 ;
        RECT 25.035000 199.650000 25.235000 199.850000 ;
        RECT 25.440000 197.250000 25.640000 197.450000 ;
        RECT 25.440000 197.650000 25.640000 197.850000 ;
        RECT 25.440000 198.050000 25.640000 198.250000 ;
        RECT 25.440000 198.450000 25.640000 198.650000 ;
        RECT 25.440000 198.850000 25.640000 199.050000 ;
        RECT 25.440000 199.250000 25.640000 199.450000 ;
        RECT 25.440000 199.650000 25.640000 199.850000 ;
        RECT 25.845000 197.250000 26.045000 197.450000 ;
        RECT 25.845000 197.650000 26.045000 197.850000 ;
        RECT 25.845000 198.050000 26.045000 198.250000 ;
        RECT 25.845000 198.450000 26.045000 198.650000 ;
        RECT 25.845000 198.850000 26.045000 199.050000 ;
        RECT 25.845000 199.250000 26.045000 199.450000 ;
        RECT 25.845000 199.650000 26.045000 199.850000 ;
        RECT 26.250000 197.250000 26.450000 197.450000 ;
        RECT 26.250000 197.650000 26.450000 197.850000 ;
        RECT 26.250000 198.050000 26.450000 198.250000 ;
        RECT 26.250000 198.450000 26.450000 198.650000 ;
        RECT 26.250000 198.850000 26.450000 199.050000 ;
        RECT 26.250000 199.250000 26.450000 199.450000 ;
        RECT 26.250000 199.650000 26.450000 199.850000 ;
        RECT 26.655000 197.250000 26.855000 197.450000 ;
        RECT 26.655000 197.650000 26.855000 197.850000 ;
        RECT 26.655000 198.050000 26.855000 198.250000 ;
        RECT 26.655000 198.450000 26.855000 198.650000 ;
        RECT 26.655000 198.850000 26.855000 199.050000 ;
        RECT 26.655000 199.250000 26.855000 199.450000 ;
        RECT 26.655000 199.650000 26.855000 199.850000 ;
        RECT 27.060000 197.250000 27.260000 197.450000 ;
        RECT 27.060000 197.650000 27.260000 197.850000 ;
        RECT 27.060000 198.050000 27.260000 198.250000 ;
        RECT 27.060000 198.450000 27.260000 198.650000 ;
        RECT 27.060000 198.850000 27.260000 199.050000 ;
        RECT 27.060000 199.250000 27.260000 199.450000 ;
        RECT 27.060000 199.650000 27.260000 199.850000 ;
        RECT 27.460000 197.250000 27.660000 197.450000 ;
        RECT 27.460000 197.650000 27.660000 197.850000 ;
        RECT 27.460000 198.050000 27.660000 198.250000 ;
        RECT 27.460000 198.450000 27.660000 198.650000 ;
        RECT 27.460000 198.850000 27.660000 199.050000 ;
        RECT 27.460000 199.250000 27.660000 199.450000 ;
        RECT 27.460000 199.650000 27.660000 199.850000 ;
        RECT 27.860000 197.250000 28.060000 197.450000 ;
        RECT 27.860000 197.650000 28.060000 197.850000 ;
        RECT 27.860000 198.050000 28.060000 198.250000 ;
        RECT 27.860000 198.450000 28.060000 198.650000 ;
        RECT 27.860000 198.850000 28.060000 199.050000 ;
        RECT 27.860000 199.250000 28.060000 199.450000 ;
        RECT 27.860000 199.650000 28.060000 199.850000 ;
        RECT 28.260000 197.250000 28.460000 197.450000 ;
        RECT 28.260000 197.650000 28.460000 197.850000 ;
        RECT 28.260000 198.050000 28.460000 198.250000 ;
        RECT 28.260000 198.450000 28.460000 198.650000 ;
        RECT 28.260000 198.850000 28.460000 199.050000 ;
        RECT 28.260000 199.250000 28.460000 199.450000 ;
        RECT 28.260000 199.650000 28.460000 199.850000 ;
        RECT 28.660000 197.250000 28.860000 197.450000 ;
        RECT 28.660000 197.650000 28.860000 197.850000 ;
        RECT 28.660000 198.050000 28.860000 198.250000 ;
        RECT 28.660000 198.450000 28.860000 198.650000 ;
        RECT 28.660000 198.850000 28.860000 199.050000 ;
        RECT 28.660000 199.250000 28.860000 199.450000 ;
        RECT 28.660000 199.650000 28.860000 199.850000 ;
        RECT 29.060000 197.250000 29.260000 197.450000 ;
        RECT 29.060000 197.650000 29.260000 197.850000 ;
        RECT 29.060000 198.050000 29.260000 198.250000 ;
        RECT 29.060000 198.450000 29.260000 198.650000 ;
        RECT 29.060000 198.850000 29.260000 199.050000 ;
        RECT 29.060000 199.250000 29.260000 199.450000 ;
        RECT 29.060000 199.650000 29.260000 199.850000 ;
        RECT 29.460000 197.250000 29.660000 197.450000 ;
        RECT 29.460000 197.650000 29.660000 197.850000 ;
        RECT 29.460000 198.050000 29.660000 198.250000 ;
        RECT 29.460000 198.450000 29.660000 198.650000 ;
        RECT 29.460000 198.850000 29.660000 199.050000 ;
        RECT 29.460000 199.250000 29.660000 199.450000 ;
        RECT 29.460000 199.650000 29.660000 199.850000 ;
        RECT 29.860000 197.250000 30.060000 197.450000 ;
        RECT 29.860000 197.650000 30.060000 197.850000 ;
        RECT 29.860000 198.050000 30.060000 198.250000 ;
        RECT 29.860000 198.450000 30.060000 198.650000 ;
        RECT 29.860000 198.850000 30.060000 199.050000 ;
        RECT 29.860000 199.250000 30.060000 199.450000 ;
        RECT 29.860000 199.650000 30.060000 199.850000 ;
        RECT 30.260000 197.250000 30.460000 197.450000 ;
        RECT 30.260000 197.650000 30.460000 197.850000 ;
        RECT 30.260000 198.050000 30.460000 198.250000 ;
        RECT 30.260000 198.450000 30.460000 198.650000 ;
        RECT 30.260000 198.850000 30.460000 199.050000 ;
        RECT 30.260000 199.250000 30.460000 199.450000 ;
        RECT 30.260000 199.650000 30.460000 199.850000 ;
        RECT 30.660000 197.250000 30.860000 197.450000 ;
        RECT 30.660000 197.650000 30.860000 197.850000 ;
        RECT 30.660000 198.050000 30.860000 198.250000 ;
        RECT 30.660000 198.450000 30.860000 198.650000 ;
        RECT 30.660000 198.850000 30.860000 199.050000 ;
        RECT 30.660000 199.250000 30.860000 199.450000 ;
        RECT 30.660000 199.650000 30.860000 199.850000 ;
        RECT 31.060000 197.250000 31.260000 197.450000 ;
        RECT 31.060000 197.650000 31.260000 197.850000 ;
        RECT 31.060000 198.050000 31.260000 198.250000 ;
        RECT 31.060000 198.450000 31.260000 198.650000 ;
        RECT 31.060000 198.850000 31.260000 199.050000 ;
        RECT 31.060000 199.250000 31.260000 199.450000 ;
        RECT 31.060000 199.650000 31.260000 199.850000 ;
        RECT 31.460000 197.250000 31.660000 197.450000 ;
        RECT 31.460000 197.650000 31.660000 197.850000 ;
        RECT 31.460000 198.050000 31.660000 198.250000 ;
        RECT 31.460000 198.450000 31.660000 198.650000 ;
        RECT 31.460000 198.850000 31.660000 199.050000 ;
        RECT 31.460000 199.250000 31.660000 199.450000 ;
        RECT 31.460000 199.650000 31.660000 199.850000 ;
        RECT 31.860000 197.250000 32.060000 197.450000 ;
        RECT 31.860000 197.650000 32.060000 197.850000 ;
        RECT 31.860000 198.050000 32.060000 198.250000 ;
        RECT 31.860000 198.450000 32.060000 198.650000 ;
        RECT 31.860000 198.850000 32.060000 199.050000 ;
        RECT 31.860000 199.250000 32.060000 199.450000 ;
        RECT 31.860000 199.650000 32.060000 199.850000 ;
        RECT 32.260000 197.250000 32.460000 197.450000 ;
        RECT 32.260000 197.650000 32.460000 197.850000 ;
        RECT 32.260000 198.050000 32.460000 198.250000 ;
        RECT 32.260000 198.450000 32.460000 198.650000 ;
        RECT 32.260000 198.850000 32.460000 199.050000 ;
        RECT 32.260000 199.250000 32.460000 199.450000 ;
        RECT 32.260000 199.650000 32.460000 199.850000 ;
        RECT 32.660000 197.250000 32.860000 197.450000 ;
        RECT 32.660000 197.650000 32.860000 197.850000 ;
        RECT 32.660000 198.050000 32.860000 198.250000 ;
        RECT 32.660000 198.450000 32.860000 198.650000 ;
        RECT 32.660000 198.850000 32.860000 199.050000 ;
        RECT 32.660000 199.250000 32.860000 199.450000 ;
        RECT 32.660000 199.650000 32.860000 199.850000 ;
        RECT 33.060000 197.250000 33.260000 197.450000 ;
        RECT 33.060000 197.650000 33.260000 197.850000 ;
        RECT 33.060000 198.050000 33.260000 198.250000 ;
        RECT 33.060000 198.450000 33.260000 198.650000 ;
        RECT 33.060000 198.850000 33.260000 199.050000 ;
        RECT 33.060000 199.250000 33.260000 199.450000 ;
        RECT 33.060000 199.650000 33.260000 199.850000 ;
        RECT 33.460000 197.250000 33.660000 197.450000 ;
        RECT 33.460000 197.650000 33.660000 197.850000 ;
        RECT 33.460000 198.050000 33.660000 198.250000 ;
        RECT 33.460000 198.450000 33.660000 198.650000 ;
        RECT 33.460000 198.850000 33.660000 199.050000 ;
        RECT 33.460000 199.250000 33.660000 199.450000 ;
        RECT 33.460000 199.650000 33.660000 199.850000 ;
        RECT 33.860000 197.250000 34.060000 197.450000 ;
        RECT 33.860000 197.650000 34.060000 197.850000 ;
        RECT 33.860000 198.050000 34.060000 198.250000 ;
        RECT 33.860000 198.450000 34.060000 198.650000 ;
        RECT 33.860000 198.850000 34.060000 199.050000 ;
        RECT 33.860000 199.250000 34.060000 199.450000 ;
        RECT 33.860000 199.650000 34.060000 199.850000 ;
        RECT 34.260000 197.250000 34.460000 197.450000 ;
        RECT 34.260000 197.650000 34.460000 197.850000 ;
        RECT 34.260000 198.050000 34.460000 198.250000 ;
        RECT 34.260000 198.450000 34.460000 198.650000 ;
        RECT 34.260000 198.850000 34.460000 199.050000 ;
        RECT 34.260000 199.250000 34.460000 199.450000 ;
        RECT 34.260000 199.650000 34.460000 199.850000 ;
        RECT 34.660000 197.250000 34.860000 197.450000 ;
        RECT 34.660000 197.650000 34.860000 197.850000 ;
        RECT 34.660000 198.050000 34.860000 198.250000 ;
        RECT 34.660000 198.450000 34.860000 198.650000 ;
        RECT 34.660000 198.850000 34.860000 199.050000 ;
        RECT 34.660000 199.250000 34.860000 199.450000 ;
        RECT 34.660000 199.650000 34.860000 199.850000 ;
        RECT 35.060000 197.250000 35.260000 197.450000 ;
        RECT 35.060000 197.650000 35.260000 197.850000 ;
        RECT 35.060000 198.050000 35.260000 198.250000 ;
        RECT 35.060000 198.450000 35.260000 198.650000 ;
        RECT 35.060000 198.850000 35.260000 199.050000 ;
        RECT 35.060000 199.250000 35.260000 199.450000 ;
        RECT 35.060000 199.650000 35.260000 199.850000 ;
        RECT 35.460000 197.250000 35.660000 197.450000 ;
        RECT 35.460000 197.650000 35.660000 197.850000 ;
        RECT 35.460000 198.050000 35.660000 198.250000 ;
        RECT 35.460000 198.450000 35.660000 198.650000 ;
        RECT 35.460000 198.850000 35.660000 199.050000 ;
        RECT 35.460000 199.250000 35.660000 199.450000 ;
        RECT 35.460000 199.650000 35.660000 199.850000 ;
        RECT 35.860000 197.250000 36.060000 197.450000 ;
        RECT 35.860000 197.650000 36.060000 197.850000 ;
        RECT 35.860000 198.050000 36.060000 198.250000 ;
        RECT 35.860000 198.450000 36.060000 198.650000 ;
        RECT 35.860000 198.850000 36.060000 199.050000 ;
        RECT 35.860000 199.250000 36.060000 199.450000 ;
        RECT 35.860000 199.650000 36.060000 199.850000 ;
        RECT 36.260000 197.250000 36.460000 197.450000 ;
        RECT 36.260000 197.650000 36.460000 197.850000 ;
        RECT 36.260000 198.050000 36.460000 198.250000 ;
        RECT 36.260000 198.450000 36.460000 198.650000 ;
        RECT 36.260000 198.850000 36.460000 199.050000 ;
        RECT 36.260000 199.250000 36.460000 199.450000 ;
        RECT 36.260000 199.650000 36.460000 199.850000 ;
        RECT 36.660000 197.250000 36.860000 197.450000 ;
        RECT 36.660000 197.650000 36.860000 197.850000 ;
        RECT 36.660000 198.050000 36.860000 198.250000 ;
        RECT 36.660000 198.450000 36.860000 198.650000 ;
        RECT 36.660000 198.850000 36.860000 199.050000 ;
        RECT 36.660000 199.250000 36.860000 199.450000 ;
        RECT 36.660000 199.650000 36.860000 199.850000 ;
        RECT 37.060000 197.250000 37.260000 197.450000 ;
        RECT 37.060000 197.650000 37.260000 197.850000 ;
        RECT 37.060000 198.050000 37.260000 198.250000 ;
        RECT 37.060000 198.450000 37.260000 198.650000 ;
        RECT 37.060000 198.850000 37.260000 199.050000 ;
        RECT 37.060000 199.250000 37.260000 199.450000 ;
        RECT 37.060000 199.650000 37.260000 199.850000 ;
        RECT 37.460000 197.250000 37.660000 197.450000 ;
        RECT 37.460000 197.650000 37.660000 197.850000 ;
        RECT 37.460000 198.050000 37.660000 198.250000 ;
        RECT 37.460000 198.450000 37.660000 198.650000 ;
        RECT 37.460000 198.850000 37.660000 199.050000 ;
        RECT 37.460000 199.250000 37.660000 199.450000 ;
        RECT 37.460000 199.650000 37.660000 199.850000 ;
        RECT 37.860000 197.250000 38.060000 197.450000 ;
        RECT 37.860000 197.650000 38.060000 197.850000 ;
        RECT 37.860000 198.050000 38.060000 198.250000 ;
        RECT 37.860000 198.450000 38.060000 198.650000 ;
        RECT 37.860000 198.850000 38.060000 199.050000 ;
        RECT 37.860000 199.250000 38.060000 199.450000 ;
        RECT 37.860000 199.650000 38.060000 199.850000 ;
        RECT 38.260000 197.250000 38.460000 197.450000 ;
        RECT 38.260000 197.650000 38.460000 197.850000 ;
        RECT 38.260000 198.050000 38.460000 198.250000 ;
        RECT 38.260000 198.450000 38.460000 198.650000 ;
        RECT 38.260000 198.850000 38.460000 199.050000 ;
        RECT 38.260000 199.250000 38.460000 199.450000 ;
        RECT 38.260000 199.650000 38.460000 199.850000 ;
        RECT 38.660000 197.250000 38.860000 197.450000 ;
        RECT 38.660000 197.650000 38.860000 197.850000 ;
        RECT 38.660000 198.050000 38.860000 198.250000 ;
        RECT 38.660000 198.450000 38.860000 198.650000 ;
        RECT 38.660000 198.850000 38.860000 199.050000 ;
        RECT 38.660000 199.250000 38.860000 199.450000 ;
        RECT 38.660000 199.650000 38.860000 199.850000 ;
        RECT 39.060000 197.250000 39.260000 197.450000 ;
        RECT 39.060000 197.650000 39.260000 197.850000 ;
        RECT 39.060000 198.050000 39.260000 198.250000 ;
        RECT 39.060000 198.450000 39.260000 198.650000 ;
        RECT 39.060000 198.850000 39.260000 199.050000 ;
        RECT 39.060000 199.250000 39.260000 199.450000 ;
        RECT 39.060000 199.650000 39.260000 199.850000 ;
        RECT 39.460000 197.250000 39.660000 197.450000 ;
        RECT 39.460000 197.650000 39.660000 197.850000 ;
        RECT 39.460000 198.050000 39.660000 198.250000 ;
        RECT 39.460000 198.450000 39.660000 198.650000 ;
        RECT 39.460000 198.850000 39.660000 199.050000 ;
        RECT 39.460000 199.250000 39.660000 199.450000 ;
        RECT 39.460000 199.650000 39.660000 199.850000 ;
        RECT 39.860000 197.250000 40.060000 197.450000 ;
        RECT 39.860000 197.650000 40.060000 197.850000 ;
        RECT 39.860000 198.050000 40.060000 198.250000 ;
        RECT 39.860000 198.450000 40.060000 198.650000 ;
        RECT 39.860000 198.850000 40.060000 199.050000 ;
        RECT 39.860000 199.250000 40.060000 199.450000 ;
        RECT 39.860000 199.650000 40.060000 199.850000 ;
        RECT 40.260000 197.250000 40.460000 197.450000 ;
        RECT 40.260000 197.650000 40.460000 197.850000 ;
        RECT 40.260000 198.050000 40.460000 198.250000 ;
        RECT 40.260000 198.450000 40.460000 198.650000 ;
        RECT 40.260000 198.850000 40.460000 199.050000 ;
        RECT 40.260000 199.250000 40.460000 199.450000 ;
        RECT 40.260000 199.650000 40.460000 199.850000 ;
        RECT 40.660000 197.250000 40.860000 197.450000 ;
        RECT 40.660000 197.650000 40.860000 197.850000 ;
        RECT 40.660000 198.050000 40.860000 198.250000 ;
        RECT 40.660000 198.450000 40.860000 198.650000 ;
        RECT 40.660000 198.850000 40.860000 199.050000 ;
        RECT 40.660000 199.250000 40.860000 199.450000 ;
        RECT 40.660000 199.650000 40.860000 199.850000 ;
        RECT 41.060000 197.250000 41.260000 197.450000 ;
        RECT 41.060000 197.650000 41.260000 197.850000 ;
        RECT 41.060000 198.050000 41.260000 198.250000 ;
        RECT 41.060000 198.450000 41.260000 198.650000 ;
        RECT 41.060000 198.850000 41.260000 199.050000 ;
        RECT 41.060000 199.250000 41.260000 199.450000 ;
        RECT 41.060000 199.650000 41.260000 199.850000 ;
        RECT 41.460000 197.250000 41.660000 197.450000 ;
        RECT 41.460000 197.650000 41.660000 197.850000 ;
        RECT 41.460000 198.050000 41.660000 198.250000 ;
        RECT 41.460000 198.450000 41.660000 198.650000 ;
        RECT 41.460000 198.850000 41.660000 199.050000 ;
        RECT 41.460000 199.250000 41.660000 199.450000 ;
        RECT 41.460000 199.650000 41.660000 199.850000 ;
        RECT 41.860000 197.250000 42.060000 197.450000 ;
        RECT 41.860000 197.650000 42.060000 197.850000 ;
        RECT 41.860000 198.050000 42.060000 198.250000 ;
        RECT 41.860000 198.450000 42.060000 198.650000 ;
        RECT 41.860000 198.850000 42.060000 199.050000 ;
        RECT 41.860000 199.250000 42.060000 199.450000 ;
        RECT 41.860000 199.650000 42.060000 199.850000 ;
        RECT 42.260000 197.250000 42.460000 197.450000 ;
        RECT 42.260000 197.650000 42.460000 197.850000 ;
        RECT 42.260000 198.050000 42.460000 198.250000 ;
        RECT 42.260000 198.450000 42.460000 198.650000 ;
        RECT 42.260000 198.850000 42.460000 199.050000 ;
        RECT 42.260000 199.250000 42.460000 199.450000 ;
        RECT 42.260000 199.650000 42.460000 199.850000 ;
        RECT 42.660000 197.250000 42.860000 197.450000 ;
        RECT 42.660000 197.650000 42.860000 197.850000 ;
        RECT 42.660000 198.050000 42.860000 198.250000 ;
        RECT 42.660000 198.450000 42.860000 198.650000 ;
        RECT 42.660000 198.850000 42.860000 199.050000 ;
        RECT 42.660000 199.250000 42.860000 199.450000 ;
        RECT 42.660000 199.650000 42.860000 199.850000 ;
        RECT 43.060000 197.250000 43.260000 197.450000 ;
        RECT 43.060000 197.650000 43.260000 197.850000 ;
        RECT 43.060000 198.050000 43.260000 198.250000 ;
        RECT 43.060000 198.450000 43.260000 198.650000 ;
        RECT 43.060000 198.850000 43.260000 199.050000 ;
        RECT 43.060000 199.250000 43.260000 199.450000 ;
        RECT 43.060000 199.650000 43.260000 199.850000 ;
        RECT 43.460000 197.250000 43.660000 197.450000 ;
        RECT 43.460000 197.650000 43.660000 197.850000 ;
        RECT 43.460000 198.050000 43.660000 198.250000 ;
        RECT 43.460000 198.450000 43.660000 198.650000 ;
        RECT 43.460000 198.850000 43.660000 199.050000 ;
        RECT 43.460000 199.250000 43.660000 199.450000 ;
        RECT 43.460000 199.650000 43.660000 199.850000 ;
        RECT 43.860000 197.250000 44.060000 197.450000 ;
        RECT 43.860000 197.650000 44.060000 197.850000 ;
        RECT 43.860000 198.050000 44.060000 198.250000 ;
        RECT 43.860000 198.450000 44.060000 198.650000 ;
        RECT 43.860000 198.850000 44.060000 199.050000 ;
        RECT 43.860000 199.250000 44.060000 199.450000 ;
        RECT 43.860000 199.650000 44.060000 199.850000 ;
        RECT 44.260000 197.250000 44.460000 197.450000 ;
        RECT 44.260000 197.650000 44.460000 197.850000 ;
        RECT 44.260000 198.050000 44.460000 198.250000 ;
        RECT 44.260000 198.450000 44.460000 198.650000 ;
        RECT 44.260000 198.850000 44.460000 199.050000 ;
        RECT 44.260000 199.250000 44.460000 199.450000 ;
        RECT 44.260000 199.650000 44.460000 199.850000 ;
        RECT 44.660000 197.250000 44.860000 197.450000 ;
        RECT 44.660000 197.650000 44.860000 197.850000 ;
        RECT 44.660000 198.050000 44.860000 198.250000 ;
        RECT 44.660000 198.450000 44.860000 198.650000 ;
        RECT 44.660000 198.850000 44.860000 199.050000 ;
        RECT 44.660000 199.250000 44.860000 199.450000 ;
        RECT 44.660000 199.650000 44.860000 199.850000 ;
        RECT 45.060000 197.250000 45.260000 197.450000 ;
        RECT 45.060000 197.650000 45.260000 197.850000 ;
        RECT 45.060000 198.050000 45.260000 198.250000 ;
        RECT 45.060000 198.450000 45.260000 198.650000 ;
        RECT 45.060000 198.850000 45.260000 199.050000 ;
        RECT 45.060000 199.250000 45.260000 199.450000 ;
        RECT 45.060000 199.650000 45.260000 199.850000 ;
        RECT 45.460000 197.250000 45.660000 197.450000 ;
        RECT 45.460000 197.650000 45.660000 197.850000 ;
        RECT 45.460000 198.050000 45.660000 198.250000 ;
        RECT 45.460000 198.450000 45.660000 198.650000 ;
        RECT 45.460000 198.850000 45.660000 199.050000 ;
        RECT 45.460000 199.250000 45.660000 199.450000 ;
        RECT 45.460000 199.650000 45.660000 199.850000 ;
        RECT 45.860000 197.250000 46.060000 197.450000 ;
        RECT 45.860000 197.650000 46.060000 197.850000 ;
        RECT 45.860000 198.050000 46.060000 198.250000 ;
        RECT 45.860000 198.450000 46.060000 198.650000 ;
        RECT 45.860000 198.850000 46.060000 199.050000 ;
        RECT 45.860000 199.250000 46.060000 199.450000 ;
        RECT 45.860000 199.650000 46.060000 199.850000 ;
        RECT 46.260000 197.250000 46.460000 197.450000 ;
        RECT 46.260000 197.650000 46.460000 197.850000 ;
        RECT 46.260000 198.050000 46.460000 198.250000 ;
        RECT 46.260000 198.450000 46.460000 198.650000 ;
        RECT 46.260000 198.850000 46.460000 199.050000 ;
        RECT 46.260000 199.250000 46.460000 199.450000 ;
        RECT 46.260000 199.650000 46.460000 199.850000 ;
        RECT 46.660000 197.250000 46.860000 197.450000 ;
        RECT 46.660000 197.650000 46.860000 197.850000 ;
        RECT 46.660000 198.050000 46.860000 198.250000 ;
        RECT 46.660000 198.450000 46.860000 198.650000 ;
        RECT 46.660000 198.850000 46.860000 199.050000 ;
        RECT 46.660000 199.250000 46.860000 199.450000 ;
        RECT 46.660000 199.650000 46.860000 199.850000 ;
        RECT 47.060000 197.250000 47.260000 197.450000 ;
        RECT 47.060000 197.650000 47.260000 197.850000 ;
        RECT 47.060000 198.050000 47.260000 198.250000 ;
        RECT 47.060000 198.450000 47.260000 198.650000 ;
        RECT 47.060000 198.850000 47.260000 199.050000 ;
        RECT 47.060000 199.250000 47.260000 199.450000 ;
        RECT 47.060000 199.650000 47.260000 199.850000 ;
        RECT 47.460000 197.250000 47.660000 197.450000 ;
        RECT 47.460000 197.650000 47.660000 197.850000 ;
        RECT 47.460000 198.050000 47.660000 198.250000 ;
        RECT 47.460000 198.450000 47.660000 198.650000 ;
        RECT 47.460000 198.850000 47.660000 199.050000 ;
        RECT 47.460000 199.250000 47.660000 199.450000 ;
        RECT 47.460000 199.650000 47.660000 199.850000 ;
        RECT 47.860000 197.250000 48.060000 197.450000 ;
        RECT 47.860000 197.650000 48.060000 197.850000 ;
        RECT 47.860000 198.050000 48.060000 198.250000 ;
        RECT 47.860000 198.450000 48.060000 198.650000 ;
        RECT 47.860000 198.850000 48.060000 199.050000 ;
        RECT 47.860000 199.250000 48.060000 199.450000 ;
        RECT 47.860000 199.650000 48.060000 199.850000 ;
        RECT 48.260000 197.250000 48.460000 197.450000 ;
        RECT 48.260000 197.650000 48.460000 197.850000 ;
        RECT 48.260000 198.050000 48.460000 198.250000 ;
        RECT 48.260000 198.450000 48.460000 198.650000 ;
        RECT 48.260000 198.850000 48.460000 199.050000 ;
        RECT 48.260000 199.250000 48.460000 199.450000 ;
        RECT 48.260000 199.650000 48.460000 199.850000 ;
        RECT 48.660000 197.250000 48.860000 197.450000 ;
        RECT 48.660000 197.650000 48.860000 197.850000 ;
        RECT 48.660000 198.050000 48.860000 198.250000 ;
        RECT 48.660000 198.450000 48.860000 198.650000 ;
        RECT 48.660000 198.850000 48.860000 199.050000 ;
        RECT 48.660000 199.250000 48.860000 199.450000 ;
        RECT 48.660000 199.650000 48.860000 199.850000 ;
        RECT 49.060000 197.250000 49.260000 197.450000 ;
        RECT 49.060000 197.650000 49.260000 197.850000 ;
        RECT 49.060000 198.050000 49.260000 198.250000 ;
        RECT 49.060000 198.450000 49.260000 198.650000 ;
        RECT 49.060000 198.850000 49.260000 199.050000 ;
        RECT 49.060000 199.250000 49.260000 199.450000 ;
        RECT 49.060000 199.650000 49.260000 199.850000 ;
        RECT 49.460000 197.250000 49.660000 197.450000 ;
        RECT 49.460000 197.650000 49.660000 197.850000 ;
        RECT 49.460000 198.050000 49.660000 198.250000 ;
        RECT 49.460000 198.450000 49.660000 198.650000 ;
        RECT 49.460000 198.850000 49.660000 199.050000 ;
        RECT 49.460000 199.250000 49.660000 199.450000 ;
        RECT 49.460000 199.650000 49.660000 199.850000 ;
        RECT 49.860000 197.250000 50.060000 197.450000 ;
        RECT 49.860000 197.650000 50.060000 197.850000 ;
        RECT 49.860000 198.050000 50.060000 198.250000 ;
        RECT 49.860000 198.450000 50.060000 198.650000 ;
        RECT 49.860000 198.850000 50.060000 199.050000 ;
        RECT 49.860000 199.250000 50.060000 199.450000 ;
        RECT 49.860000 199.650000 50.060000 199.850000 ;
        RECT 50.260000 197.250000 50.460000 197.450000 ;
        RECT 50.260000 197.650000 50.460000 197.850000 ;
        RECT 50.260000 198.050000 50.460000 198.250000 ;
        RECT 50.260000 198.450000 50.460000 198.650000 ;
        RECT 50.260000 198.850000 50.460000 199.050000 ;
        RECT 50.260000 199.250000 50.460000 199.450000 ;
        RECT 50.260000 199.650000 50.460000 199.850000 ;
        RECT 50.480000  25.910000 50.680000  26.110000 ;
        RECT 50.480000  26.340000 50.680000  26.540000 ;
        RECT 50.480000  26.770000 50.680000  26.970000 ;
        RECT 50.480000  27.200000 50.680000  27.400000 ;
        RECT 50.480000  27.630000 50.680000  27.830000 ;
        RECT 50.480000  28.060000 50.680000  28.260000 ;
        RECT 50.480000  28.490000 50.680000  28.690000 ;
        RECT 50.480000  28.920000 50.680000  29.120000 ;
        RECT 50.480000  29.350000 50.680000  29.550000 ;
        RECT 50.480000  29.780000 50.680000  29.980000 ;
        RECT 50.480000  30.210000 50.680000  30.410000 ;
        RECT 50.660000 197.250000 50.860000 197.450000 ;
        RECT 50.660000 197.650000 50.860000 197.850000 ;
        RECT 50.660000 198.050000 50.860000 198.250000 ;
        RECT 50.660000 198.450000 50.860000 198.650000 ;
        RECT 50.660000 198.850000 50.860000 199.050000 ;
        RECT 50.660000 199.250000 50.860000 199.450000 ;
        RECT 50.660000 199.650000 50.860000 199.850000 ;
        RECT 50.890000  25.910000 51.090000  26.110000 ;
        RECT 50.890000  26.340000 51.090000  26.540000 ;
        RECT 50.890000  26.770000 51.090000  26.970000 ;
        RECT 50.890000  27.200000 51.090000  27.400000 ;
        RECT 50.890000  27.630000 51.090000  27.830000 ;
        RECT 50.890000  28.060000 51.090000  28.260000 ;
        RECT 50.890000  28.490000 51.090000  28.690000 ;
        RECT 50.890000  28.920000 51.090000  29.120000 ;
        RECT 50.890000  29.350000 51.090000  29.550000 ;
        RECT 50.890000  29.780000 51.090000  29.980000 ;
        RECT 50.890000  30.210000 51.090000  30.410000 ;
        RECT 51.060000 197.250000 51.260000 197.450000 ;
        RECT 51.060000 197.650000 51.260000 197.850000 ;
        RECT 51.060000 198.050000 51.260000 198.250000 ;
        RECT 51.060000 198.450000 51.260000 198.650000 ;
        RECT 51.060000 198.850000 51.260000 199.050000 ;
        RECT 51.060000 199.250000 51.260000 199.450000 ;
        RECT 51.060000 199.650000 51.260000 199.850000 ;
        RECT 51.300000  25.910000 51.500000  26.110000 ;
        RECT 51.300000  26.340000 51.500000  26.540000 ;
        RECT 51.300000  26.770000 51.500000  26.970000 ;
        RECT 51.300000  27.200000 51.500000  27.400000 ;
        RECT 51.300000  27.630000 51.500000  27.830000 ;
        RECT 51.300000  28.060000 51.500000  28.260000 ;
        RECT 51.300000  28.490000 51.500000  28.690000 ;
        RECT 51.300000  28.920000 51.500000  29.120000 ;
        RECT 51.300000  29.350000 51.500000  29.550000 ;
        RECT 51.300000  29.780000 51.500000  29.980000 ;
        RECT 51.300000  30.210000 51.500000  30.410000 ;
        RECT 51.460000 197.250000 51.660000 197.450000 ;
        RECT 51.460000 197.650000 51.660000 197.850000 ;
        RECT 51.460000 198.050000 51.660000 198.250000 ;
        RECT 51.460000 198.450000 51.660000 198.650000 ;
        RECT 51.460000 198.850000 51.660000 199.050000 ;
        RECT 51.460000 199.250000 51.660000 199.450000 ;
        RECT 51.460000 199.650000 51.660000 199.850000 ;
        RECT 51.710000  25.910000 51.910000  26.110000 ;
        RECT 51.710000  26.340000 51.910000  26.540000 ;
        RECT 51.710000  26.770000 51.910000  26.970000 ;
        RECT 51.710000  27.200000 51.910000  27.400000 ;
        RECT 51.710000  27.630000 51.910000  27.830000 ;
        RECT 51.710000  28.060000 51.910000  28.260000 ;
        RECT 51.710000  28.490000 51.910000  28.690000 ;
        RECT 51.710000  28.920000 51.910000  29.120000 ;
        RECT 51.710000  29.350000 51.910000  29.550000 ;
        RECT 51.710000  29.780000 51.910000  29.980000 ;
        RECT 51.710000  30.210000 51.910000  30.410000 ;
        RECT 51.860000 197.250000 52.060000 197.450000 ;
        RECT 51.860000 197.650000 52.060000 197.850000 ;
        RECT 51.860000 198.050000 52.060000 198.250000 ;
        RECT 51.860000 198.450000 52.060000 198.650000 ;
        RECT 51.860000 198.850000 52.060000 199.050000 ;
        RECT 51.860000 199.250000 52.060000 199.450000 ;
        RECT 51.860000 199.650000 52.060000 199.850000 ;
        RECT 52.120000  25.910000 52.320000  26.110000 ;
        RECT 52.120000  26.340000 52.320000  26.540000 ;
        RECT 52.120000  26.770000 52.320000  26.970000 ;
        RECT 52.120000  27.200000 52.320000  27.400000 ;
        RECT 52.120000  27.630000 52.320000  27.830000 ;
        RECT 52.120000  28.060000 52.320000  28.260000 ;
        RECT 52.120000  28.490000 52.320000  28.690000 ;
        RECT 52.120000  28.920000 52.320000  29.120000 ;
        RECT 52.120000  29.350000 52.320000  29.550000 ;
        RECT 52.120000  29.780000 52.320000  29.980000 ;
        RECT 52.120000  30.210000 52.320000  30.410000 ;
        RECT 52.260000 197.250000 52.460000 197.450000 ;
        RECT 52.260000 197.650000 52.460000 197.850000 ;
        RECT 52.260000 198.050000 52.460000 198.250000 ;
        RECT 52.260000 198.450000 52.460000 198.650000 ;
        RECT 52.260000 198.850000 52.460000 199.050000 ;
        RECT 52.260000 199.250000 52.460000 199.450000 ;
        RECT 52.260000 199.650000 52.460000 199.850000 ;
        RECT 52.530000  25.910000 52.730000  26.110000 ;
        RECT 52.530000  26.340000 52.730000  26.540000 ;
        RECT 52.530000  26.770000 52.730000  26.970000 ;
        RECT 52.530000  27.200000 52.730000  27.400000 ;
        RECT 52.530000  27.630000 52.730000  27.830000 ;
        RECT 52.530000  28.060000 52.730000  28.260000 ;
        RECT 52.530000  28.490000 52.730000  28.690000 ;
        RECT 52.530000  28.920000 52.730000  29.120000 ;
        RECT 52.530000  29.350000 52.730000  29.550000 ;
        RECT 52.530000  29.780000 52.730000  29.980000 ;
        RECT 52.530000  30.210000 52.730000  30.410000 ;
        RECT 52.660000 197.250000 52.860000 197.450000 ;
        RECT 52.660000 197.650000 52.860000 197.850000 ;
        RECT 52.660000 198.050000 52.860000 198.250000 ;
        RECT 52.660000 198.450000 52.860000 198.650000 ;
        RECT 52.660000 198.850000 52.860000 199.050000 ;
        RECT 52.660000 199.250000 52.860000 199.450000 ;
        RECT 52.660000 199.650000 52.860000 199.850000 ;
        RECT 52.940000  25.910000 53.140000  26.110000 ;
        RECT 52.940000  26.340000 53.140000  26.540000 ;
        RECT 52.940000  26.770000 53.140000  26.970000 ;
        RECT 52.940000  27.200000 53.140000  27.400000 ;
        RECT 52.940000  27.630000 53.140000  27.830000 ;
        RECT 52.940000  28.060000 53.140000  28.260000 ;
        RECT 52.940000  28.490000 53.140000  28.690000 ;
        RECT 52.940000  28.920000 53.140000  29.120000 ;
        RECT 52.940000  29.350000 53.140000  29.550000 ;
        RECT 52.940000  29.780000 53.140000  29.980000 ;
        RECT 52.940000  30.210000 53.140000  30.410000 ;
        RECT 53.060000 197.250000 53.260000 197.450000 ;
        RECT 53.060000 197.650000 53.260000 197.850000 ;
        RECT 53.060000 198.050000 53.260000 198.250000 ;
        RECT 53.060000 198.450000 53.260000 198.650000 ;
        RECT 53.060000 198.850000 53.260000 199.050000 ;
        RECT 53.060000 199.250000 53.260000 199.450000 ;
        RECT 53.060000 199.650000 53.260000 199.850000 ;
        RECT 53.345000  25.910000 53.545000  26.110000 ;
        RECT 53.345000  26.340000 53.545000  26.540000 ;
        RECT 53.345000  26.770000 53.545000  26.970000 ;
        RECT 53.345000  27.200000 53.545000  27.400000 ;
        RECT 53.345000  27.630000 53.545000  27.830000 ;
        RECT 53.345000  28.060000 53.545000  28.260000 ;
        RECT 53.345000  28.490000 53.545000  28.690000 ;
        RECT 53.345000  28.920000 53.545000  29.120000 ;
        RECT 53.345000  29.350000 53.545000  29.550000 ;
        RECT 53.345000  29.780000 53.545000  29.980000 ;
        RECT 53.345000  30.210000 53.545000  30.410000 ;
        RECT 53.460000 197.250000 53.660000 197.450000 ;
        RECT 53.460000 197.650000 53.660000 197.850000 ;
        RECT 53.460000 198.050000 53.660000 198.250000 ;
        RECT 53.460000 198.450000 53.660000 198.650000 ;
        RECT 53.460000 198.850000 53.660000 199.050000 ;
        RECT 53.460000 199.250000 53.660000 199.450000 ;
        RECT 53.460000 199.650000 53.660000 199.850000 ;
        RECT 53.750000  25.910000 53.950000  26.110000 ;
        RECT 53.750000  26.340000 53.950000  26.540000 ;
        RECT 53.750000  26.770000 53.950000  26.970000 ;
        RECT 53.750000  27.200000 53.950000  27.400000 ;
        RECT 53.750000  27.630000 53.950000  27.830000 ;
        RECT 53.750000  28.060000 53.950000  28.260000 ;
        RECT 53.750000  28.490000 53.950000  28.690000 ;
        RECT 53.750000  28.920000 53.950000  29.120000 ;
        RECT 53.750000  29.350000 53.950000  29.550000 ;
        RECT 53.750000  29.780000 53.950000  29.980000 ;
        RECT 53.750000  30.210000 53.950000  30.410000 ;
        RECT 53.860000 197.250000 54.060000 197.450000 ;
        RECT 53.860000 197.650000 54.060000 197.850000 ;
        RECT 53.860000 198.050000 54.060000 198.250000 ;
        RECT 53.860000 198.450000 54.060000 198.650000 ;
        RECT 53.860000 198.850000 54.060000 199.050000 ;
        RECT 53.860000 199.250000 54.060000 199.450000 ;
        RECT 53.860000 199.650000 54.060000 199.850000 ;
        RECT 54.155000  25.910000 54.355000  26.110000 ;
        RECT 54.155000  26.340000 54.355000  26.540000 ;
        RECT 54.155000  26.770000 54.355000  26.970000 ;
        RECT 54.155000  27.200000 54.355000  27.400000 ;
        RECT 54.155000  27.630000 54.355000  27.830000 ;
        RECT 54.155000  28.060000 54.355000  28.260000 ;
        RECT 54.155000  28.490000 54.355000  28.690000 ;
        RECT 54.155000  28.920000 54.355000  29.120000 ;
        RECT 54.155000  29.350000 54.355000  29.550000 ;
        RECT 54.155000  29.780000 54.355000  29.980000 ;
        RECT 54.155000  30.210000 54.355000  30.410000 ;
        RECT 54.260000 197.250000 54.460000 197.450000 ;
        RECT 54.260000 197.650000 54.460000 197.850000 ;
        RECT 54.260000 198.050000 54.460000 198.250000 ;
        RECT 54.260000 198.450000 54.460000 198.650000 ;
        RECT 54.260000 198.850000 54.460000 199.050000 ;
        RECT 54.260000 199.250000 54.460000 199.450000 ;
        RECT 54.260000 199.650000 54.460000 199.850000 ;
        RECT 54.560000  25.910000 54.760000  26.110000 ;
        RECT 54.560000  26.340000 54.760000  26.540000 ;
        RECT 54.560000  26.770000 54.760000  26.970000 ;
        RECT 54.560000  27.200000 54.760000  27.400000 ;
        RECT 54.560000  27.630000 54.760000  27.830000 ;
        RECT 54.560000  28.060000 54.760000  28.260000 ;
        RECT 54.560000  28.490000 54.760000  28.690000 ;
        RECT 54.560000  28.920000 54.760000  29.120000 ;
        RECT 54.560000  29.350000 54.760000  29.550000 ;
        RECT 54.560000  29.780000 54.760000  29.980000 ;
        RECT 54.560000  30.210000 54.760000  30.410000 ;
        RECT 54.660000 197.250000 54.860000 197.450000 ;
        RECT 54.660000 197.650000 54.860000 197.850000 ;
        RECT 54.660000 198.050000 54.860000 198.250000 ;
        RECT 54.660000 198.450000 54.860000 198.650000 ;
        RECT 54.660000 198.850000 54.860000 199.050000 ;
        RECT 54.660000 199.250000 54.860000 199.450000 ;
        RECT 54.660000 199.650000 54.860000 199.850000 ;
        RECT 54.965000  25.910000 55.165000  26.110000 ;
        RECT 54.965000  26.340000 55.165000  26.540000 ;
        RECT 54.965000  26.770000 55.165000  26.970000 ;
        RECT 54.965000  27.200000 55.165000  27.400000 ;
        RECT 54.965000  27.630000 55.165000  27.830000 ;
        RECT 54.965000  28.060000 55.165000  28.260000 ;
        RECT 54.965000  28.490000 55.165000  28.690000 ;
        RECT 54.965000  28.920000 55.165000  29.120000 ;
        RECT 54.965000  29.350000 55.165000  29.550000 ;
        RECT 54.965000  29.780000 55.165000  29.980000 ;
        RECT 54.965000  30.210000 55.165000  30.410000 ;
        RECT 55.060000 197.250000 55.260000 197.450000 ;
        RECT 55.060000 197.650000 55.260000 197.850000 ;
        RECT 55.060000 198.050000 55.260000 198.250000 ;
        RECT 55.060000 198.450000 55.260000 198.650000 ;
        RECT 55.060000 198.850000 55.260000 199.050000 ;
        RECT 55.060000 199.250000 55.260000 199.450000 ;
        RECT 55.060000 199.650000 55.260000 199.850000 ;
        RECT 55.370000  25.910000 55.570000  26.110000 ;
        RECT 55.370000  26.340000 55.570000  26.540000 ;
        RECT 55.370000  26.770000 55.570000  26.970000 ;
        RECT 55.370000  27.200000 55.570000  27.400000 ;
        RECT 55.370000  27.630000 55.570000  27.830000 ;
        RECT 55.370000  28.060000 55.570000  28.260000 ;
        RECT 55.370000  28.490000 55.570000  28.690000 ;
        RECT 55.370000  28.920000 55.570000  29.120000 ;
        RECT 55.370000  29.350000 55.570000  29.550000 ;
        RECT 55.370000  29.780000 55.570000  29.980000 ;
        RECT 55.370000  30.210000 55.570000  30.410000 ;
        RECT 55.460000 197.250000 55.660000 197.450000 ;
        RECT 55.460000 197.650000 55.660000 197.850000 ;
        RECT 55.460000 198.050000 55.660000 198.250000 ;
        RECT 55.460000 198.450000 55.660000 198.650000 ;
        RECT 55.460000 198.850000 55.660000 199.050000 ;
        RECT 55.460000 199.250000 55.660000 199.450000 ;
        RECT 55.460000 199.650000 55.660000 199.850000 ;
        RECT 55.775000  25.910000 55.975000  26.110000 ;
        RECT 55.775000  26.340000 55.975000  26.540000 ;
        RECT 55.775000  26.770000 55.975000  26.970000 ;
        RECT 55.775000  27.200000 55.975000  27.400000 ;
        RECT 55.775000  27.630000 55.975000  27.830000 ;
        RECT 55.775000  28.060000 55.975000  28.260000 ;
        RECT 55.775000  28.490000 55.975000  28.690000 ;
        RECT 55.775000  28.920000 55.975000  29.120000 ;
        RECT 55.775000  29.350000 55.975000  29.550000 ;
        RECT 55.775000  29.780000 55.975000  29.980000 ;
        RECT 55.775000  30.210000 55.975000  30.410000 ;
        RECT 55.860000 197.250000 56.060000 197.450000 ;
        RECT 55.860000 197.650000 56.060000 197.850000 ;
        RECT 55.860000 198.050000 56.060000 198.250000 ;
        RECT 55.860000 198.450000 56.060000 198.650000 ;
        RECT 55.860000 198.850000 56.060000 199.050000 ;
        RECT 55.860000 199.250000 56.060000 199.450000 ;
        RECT 55.860000 199.650000 56.060000 199.850000 ;
        RECT 56.180000  25.910000 56.380000  26.110000 ;
        RECT 56.180000  26.340000 56.380000  26.540000 ;
        RECT 56.180000  26.770000 56.380000  26.970000 ;
        RECT 56.180000  27.200000 56.380000  27.400000 ;
        RECT 56.180000  27.630000 56.380000  27.830000 ;
        RECT 56.180000  28.060000 56.380000  28.260000 ;
        RECT 56.180000  28.490000 56.380000  28.690000 ;
        RECT 56.180000  28.920000 56.380000  29.120000 ;
        RECT 56.180000  29.350000 56.380000  29.550000 ;
        RECT 56.180000  29.780000 56.380000  29.980000 ;
        RECT 56.180000  30.210000 56.380000  30.410000 ;
        RECT 56.260000 197.250000 56.460000 197.450000 ;
        RECT 56.260000 197.650000 56.460000 197.850000 ;
        RECT 56.260000 198.050000 56.460000 198.250000 ;
        RECT 56.260000 198.450000 56.460000 198.650000 ;
        RECT 56.260000 198.850000 56.460000 199.050000 ;
        RECT 56.260000 199.250000 56.460000 199.450000 ;
        RECT 56.260000 199.650000 56.460000 199.850000 ;
        RECT 56.585000  25.910000 56.785000  26.110000 ;
        RECT 56.585000  26.340000 56.785000  26.540000 ;
        RECT 56.585000  26.770000 56.785000  26.970000 ;
        RECT 56.585000  27.200000 56.785000  27.400000 ;
        RECT 56.585000  27.630000 56.785000  27.830000 ;
        RECT 56.585000  28.060000 56.785000  28.260000 ;
        RECT 56.585000  28.490000 56.785000  28.690000 ;
        RECT 56.585000  28.920000 56.785000  29.120000 ;
        RECT 56.585000  29.350000 56.785000  29.550000 ;
        RECT 56.585000  29.780000 56.785000  29.980000 ;
        RECT 56.585000  30.210000 56.785000  30.410000 ;
        RECT 56.660000 197.250000 56.860000 197.450000 ;
        RECT 56.660000 197.650000 56.860000 197.850000 ;
        RECT 56.660000 198.050000 56.860000 198.250000 ;
        RECT 56.660000 198.450000 56.860000 198.650000 ;
        RECT 56.660000 198.850000 56.860000 199.050000 ;
        RECT 56.660000 199.250000 56.860000 199.450000 ;
        RECT 56.660000 199.650000 56.860000 199.850000 ;
        RECT 56.990000  25.910000 57.190000  26.110000 ;
        RECT 56.990000  26.340000 57.190000  26.540000 ;
        RECT 56.990000  26.770000 57.190000  26.970000 ;
        RECT 56.990000  27.200000 57.190000  27.400000 ;
        RECT 56.990000  27.630000 57.190000  27.830000 ;
        RECT 56.990000  28.060000 57.190000  28.260000 ;
        RECT 56.990000  28.490000 57.190000  28.690000 ;
        RECT 56.990000  28.920000 57.190000  29.120000 ;
        RECT 56.990000  29.350000 57.190000  29.550000 ;
        RECT 56.990000  29.780000 57.190000  29.980000 ;
        RECT 56.990000  30.210000 57.190000  30.410000 ;
        RECT 57.060000 197.250000 57.260000 197.450000 ;
        RECT 57.060000 197.650000 57.260000 197.850000 ;
        RECT 57.060000 198.050000 57.260000 198.250000 ;
        RECT 57.060000 198.450000 57.260000 198.650000 ;
        RECT 57.060000 198.850000 57.260000 199.050000 ;
        RECT 57.060000 199.250000 57.260000 199.450000 ;
        RECT 57.060000 199.650000 57.260000 199.850000 ;
        RECT 57.395000  25.910000 57.595000  26.110000 ;
        RECT 57.395000  26.340000 57.595000  26.540000 ;
        RECT 57.395000  26.770000 57.595000  26.970000 ;
        RECT 57.395000  27.200000 57.595000  27.400000 ;
        RECT 57.395000  27.630000 57.595000  27.830000 ;
        RECT 57.395000  28.060000 57.595000  28.260000 ;
        RECT 57.395000  28.490000 57.595000  28.690000 ;
        RECT 57.395000  28.920000 57.595000  29.120000 ;
        RECT 57.395000  29.350000 57.595000  29.550000 ;
        RECT 57.395000  29.780000 57.595000  29.980000 ;
        RECT 57.395000  30.210000 57.595000  30.410000 ;
        RECT 57.460000 197.250000 57.660000 197.450000 ;
        RECT 57.460000 197.650000 57.660000 197.850000 ;
        RECT 57.460000 198.050000 57.660000 198.250000 ;
        RECT 57.460000 198.450000 57.660000 198.650000 ;
        RECT 57.460000 198.850000 57.660000 199.050000 ;
        RECT 57.460000 199.250000 57.660000 199.450000 ;
        RECT 57.460000 199.650000 57.660000 199.850000 ;
        RECT 57.800000  25.910000 58.000000  26.110000 ;
        RECT 57.800000  26.340000 58.000000  26.540000 ;
        RECT 57.800000  26.770000 58.000000  26.970000 ;
        RECT 57.800000  27.200000 58.000000  27.400000 ;
        RECT 57.800000  27.630000 58.000000  27.830000 ;
        RECT 57.800000  28.060000 58.000000  28.260000 ;
        RECT 57.800000  28.490000 58.000000  28.690000 ;
        RECT 57.800000  28.920000 58.000000  29.120000 ;
        RECT 57.800000  29.350000 58.000000  29.550000 ;
        RECT 57.800000  29.780000 58.000000  29.980000 ;
        RECT 57.800000  30.210000 58.000000  30.410000 ;
        RECT 57.860000 197.250000 58.060000 197.450000 ;
        RECT 57.860000 197.650000 58.060000 197.850000 ;
        RECT 57.860000 198.050000 58.060000 198.250000 ;
        RECT 57.860000 198.450000 58.060000 198.650000 ;
        RECT 57.860000 198.850000 58.060000 199.050000 ;
        RECT 57.860000 199.250000 58.060000 199.450000 ;
        RECT 57.860000 199.650000 58.060000 199.850000 ;
        RECT 58.205000  25.910000 58.405000  26.110000 ;
        RECT 58.205000  26.340000 58.405000  26.540000 ;
        RECT 58.205000  26.770000 58.405000  26.970000 ;
        RECT 58.205000  27.200000 58.405000  27.400000 ;
        RECT 58.205000  27.630000 58.405000  27.830000 ;
        RECT 58.205000  28.060000 58.405000  28.260000 ;
        RECT 58.205000  28.490000 58.405000  28.690000 ;
        RECT 58.205000  28.920000 58.405000  29.120000 ;
        RECT 58.205000  29.350000 58.405000  29.550000 ;
        RECT 58.205000  29.780000 58.405000  29.980000 ;
        RECT 58.205000  30.210000 58.405000  30.410000 ;
        RECT 58.260000 197.250000 58.460000 197.450000 ;
        RECT 58.260000 197.650000 58.460000 197.850000 ;
        RECT 58.260000 198.050000 58.460000 198.250000 ;
        RECT 58.260000 198.450000 58.460000 198.650000 ;
        RECT 58.260000 198.850000 58.460000 199.050000 ;
        RECT 58.260000 199.250000 58.460000 199.450000 ;
        RECT 58.260000 199.650000 58.460000 199.850000 ;
        RECT 58.610000  25.910000 58.810000  26.110000 ;
        RECT 58.610000  26.340000 58.810000  26.540000 ;
        RECT 58.610000  26.770000 58.810000  26.970000 ;
        RECT 58.610000  27.200000 58.810000  27.400000 ;
        RECT 58.610000  27.630000 58.810000  27.830000 ;
        RECT 58.610000  28.060000 58.810000  28.260000 ;
        RECT 58.610000  28.490000 58.810000  28.690000 ;
        RECT 58.610000  28.920000 58.810000  29.120000 ;
        RECT 58.610000  29.350000 58.810000  29.550000 ;
        RECT 58.610000  29.780000 58.810000  29.980000 ;
        RECT 58.610000  30.210000 58.810000  30.410000 ;
        RECT 58.660000 197.250000 58.860000 197.450000 ;
        RECT 58.660000 197.650000 58.860000 197.850000 ;
        RECT 58.660000 198.050000 58.860000 198.250000 ;
        RECT 58.660000 198.450000 58.860000 198.650000 ;
        RECT 58.660000 198.850000 58.860000 199.050000 ;
        RECT 58.660000 199.250000 58.860000 199.450000 ;
        RECT 58.660000 199.650000 58.860000 199.850000 ;
        RECT 59.015000  25.910000 59.215000  26.110000 ;
        RECT 59.015000  26.340000 59.215000  26.540000 ;
        RECT 59.015000  26.770000 59.215000  26.970000 ;
        RECT 59.015000  27.200000 59.215000  27.400000 ;
        RECT 59.015000  27.630000 59.215000  27.830000 ;
        RECT 59.015000  28.060000 59.215000  28.260000 ;
        RECT 59.015000  28.490000 59.215000  28.690000 ;
        RECT 59.015000  28.920000 59.215000  29.120000 ;
        RECT 59.015000  29.350000 59.215000  29.550000 ;
        RECT 59.015000  29.780000 59.215000  29.980000 ;
        RECT 59.015000  30.210000 59.215000  30.410000 ;
        RECT 59.060000 197.250000 59.260000 197.450000 ;
        RECT 59.060000 197.650000 59.260000 197.850000 ;
        RECT 59.060000 198.050000 59.260000 198.250000 ;
        RECT 59.060000 198.450000 59.260000 198.650000 ;
        RECT 59.060000 198.850000 59.260000 199.050000 ;
        RECT 59.060000 199.250000 59.260000 199.450000 ;
        RECT 59.060000 199.650000 59.260000 199.850000 ;
        RECT 59.420000  25.910000 59.620000  26.110000 ;
        RECT 59.420000  26.340000 59.620000  26.540000 ;
        RECT 59.420000  26.770000 59.620000  26.970000 ;
        RECT 59.420000  27.200000 59.620000  27.400000 ;
        RECT 59.420000  27.630000 59.620000  27.830000 ;
        RECT 59.420000  28.060000 59.620000  28.260000 ;
        RECT 59.420000  28.490000 59.620000  28.690000 ;
        RECT 59.420000  28.920000 59.620000  29.120000 ;
        RECT 59.420000  29.350000 59.620000  29.550000 ;
        RECT 59.420000  29.780000 59.620000  29.980000 ;
        RECT 59.420000  30.210000 59.620000  30.410000 ;
        RECT 59.460000 197.250000 59.660000 197.450000 ;
        RECT 59.460000 197.650000 59.660000 197.850000 ;
        RECT 59.460000 198.050000 59.660000 198.250000 ;
        RECT 59.460000 198.450000 59.660000 198.650000 ;
        RECT 59.460000 198.850000 59.660000 199.050000 ;
        RECT 59.460000 199.250000 59.660000 199.450000 ;
        RECT 59.460000 199.650000 59.660000 199.850000 ;
        RECT 59.825000  25.910000 60.025000  26.110000 ;
        RECT 59.825000  26.340000 60.025000  26.540000 ;
        RECT 59.825000  26.770000 60.025000  26.970000 ;
        RECT 59.825000  27.200000 60.025000  27.400000 ;
        RECT 59.825000  27.630000 60.025000  27.830000 ;
        RECT 59.825000  28.060000 60.025000  28.260000 ;
        RECT 59.825000  28.490000 60.025000  28.690000 ;
        RECT 59.825000  28.920000 60.025000  29.120000 ;
        RECT 59.825000  29.350000 60.025000  29.550000 ;
        RECT 59.825000  29.780000 60.025000  29.980000 ;
        RECT 59.825000  30.210000 60.025000  30.410000 ;
        RECT 59.860000 197.250000 60.060000 197.450000 ;
        RECT 59.860000 197.650000 60.060000 197.850000 ;
        RECT 59.860000 198.050000 60.060000 198.250000 ;
        RECT 59.860000 198.450000 60.060000 198.650000 ;
        RECT 59.860000 198.850000 60.060000 199.050000 ;
        RECT 59.860000 199.250000 60.060000 199.450000 ;
        RECT 59.860000 199.650000 60.060000 199.850000 ;
        RECT 60.230000  25.910000 60.430000  26.110000 ;
        RECT 60.230000  26.340000 60.430000  26.540000 ;
        RECT 60.230000  26.770000 60.430000  26.970000 ;
        RECT 60.230000  27.200000 60.430000  27.400000 ;
        RECT 60.230000  27.630000 60.430000  27.830000 ;
        RECT 60.230000  28.060000 60.430000  28.260000 ;
        RECT 60.230000  28.490000 60.430000  28.690000 ;
        RECT 60.230000  28.920000 60.430000  29.120000 ;
        RECT 60.230000  29.350000 60.430000  29.550000 ;
        RECT 60.230000  29.780000 60.430000  29.980000 ;
        RECT 60.230000  30.210000 60.430000  30.410000 ;
        RECT 60.260000 197.250000 60.460000 197.450000 ;
        RECT 60.260000 197.650000 60.460000 197.850000 ;
        RECT 60.260000 198.050000 60.460000 198.250000 ;
        RECT 60.260000 198.450000 60.460000 198.650000 ;
        RECT 60.260000 198.850000 60.460000 199.050000 ;
        RECT 60.260000 199.250000 60.460000 199.450000 ;
        RECT 60.260000 199.650000 60.460000 199.850000 ;
        RECT 60.635000  25.910000 60.835000  26.110000 ;
        RECT 60.635000  26.340000 60.835000  26.540000 ;
        RECT 60.635000  26.770000 60.835000  26.970000 ;
        RECT 60.635000  27.200000 60.835000  27.400000 ;
        RECT 60.635000  27.630000 60.835000  27.830000 ;
        RECT 60.635000  28.060000 60.835000  28.260000 ;
        RECT 60.635000  28.490000 60.835000  28.690000 ;
        RECT 60.635000  28.920000 60.835000  29.120000 ;
        RECT 60.635000  29.350000 60.835000  29.550000 ;
        RECT 60.635000  29.780000 60.835000  29.980000 ;
        RECT 60.635000  30.210000 60.835000  30.410000 ;
        RECT 60.660000 197.250000 60.860000 197.450000 ;
        RECT 60.660000 197.650000 60.860000 197.850000 ;
        RECT 60.660000 198.050000 60.860000 198.250000 ;
        RECT 60.660000 198.450000 60.860000 198.650000 ;
        RECT 60.660000 198.850000 60.860000 199.050000 ;
        RECT 60.660000 199.250000 60.860000 199.450000 ;
        RECT 60.660000 199.650000 60.860000 199.850000 ;
        RECT 60.910000 196.295000 61.110000 196.495000 ;
        RECT 60.910000 196.705000 61.110000 196.905000 ;
        RECT 61.040000  25.910000 61.240000  26.110000 ;
        RECT 61.040000  26.340000 61.240000  26.540000 ;
        RECT 61.040000  26.770000 61.240000  26.970000 ;
        RECT 61.040000  27.200000 61.240000  27.400000 ;
        RECT 61.040000  27.630000 61.240000  27.830000 ;
        RECT 61.040000  28.060000 61.240000  28.260000 ;
        RECT 61.040000  28.490000 61.240000  28.690000 ;
        RECT 61.040000  28.920000 61.240000  29.120000 ;
        RECT 61.040000  29.350000 61.240000  29.550000 ;
        RECT 61.040000  29.780000 61.240000  29.980000 ;
        RECT 61.040000  30.210000 61.240000  30.410000 ;
        RECT 61.060000 197.250000 61.260000 197.450000 ;
        RECT 61.060000 197.650000 61.260000 197.850000 ;
        RECT 61.060000 198.050000 61.260000 198.250000 ;
        RECT 61.060000 198.450000 61.260000 198.650000 ;
        RECT 61.060000 198.850000 61.260000 199.050000 ;
        RECT 61.060000 199.250000 61.260000 199.450000 ;
        RECT 61.060000 199.650000 61.260000 199.850000 ;
        RECT 61.445000  25.910000 61.645000  26.110000 ;
        RECT 61.445000  26.340000 61.645000  26.540000 ;
        RECT 61.445000  26.770000 61.645000  26.970000 ;
        RECT 61.445000  27.200000 61.645000  27.400000 ;
        RECT 61.445000  27.630000 61.645000  27.830000 ;
        RECT 61.445000  28.060000 61.645000  28.260000 ;
        RECT 61.445000  28.490000 61.645000  28.690000 ;
        RECT 61.445000  28.920000 61.645000  29.120000 ;
        RECT 61.445000  29.350000 61.645000  29.550000 ;
        RECT 61.445000  29.780000 61.645000  29.980000 ;
        RECT 61.445000  30.210000 61.645000  30.410000 ;
        RECT 61.590000 175.995000 61.790000 176.195000 ;
        RECT 61.590000 176.395000 61.790000 176.595000 ;
        RECT 61.590000 176.795000 61.790000 176.995000 ;
        RECT 61.590000 177.195000 61.790000 177.395000 ;
        RECT 61.590000 177.595000 61.790000 177.795000 ;
        RECT 61.590000 177.995000 61.790000 178.195000 ;
        RECT 61.590000 178.395000 61.790000 178.595000 ;
        RECT 61.590000 178.795000 61.790000 178.995000 ;
        RECT 61.590000 179.195000 61.790000 179.395000 ;
        RECT 61.590000 179.595000 61.790000 179.795000 ;
        RECT 61.590000 179.995000 61.790000 180.195000 ;
        RECT 61.590000 180.395000 61.790000 180.595000 ;
        RECT 61.590000 180.795000 61.790000 180.995000 ;
        RECT 61.590000 181.195000 61.790000 181.395000 ;
        RECT 61.590000 181.595000 61.790000 181.795000 ;
        RECT 61.590000 181.995000 61.790000 182.195000 ;
        RECT 61.590000 182.395000 61.790000 182.595000 ;
        RECT 61.590000 182.795000 61.790000 182.995000 ;
        RECT 61.590000 183.195000 61.790000 183.395000 ;
        RECT 61.590000 183.595000 61.790000 183.795000 ;
        RECT 61.590000 183.995000 61.790000 184.195000 ;
        RECT 61.590000 184.395000 61.790000 184.595000 ;
        RECT 61.590000 184.795000 61.790000 184.995000 ;
        RECT 61.590000 185.195000 61.790000 185.395000 ;
        RECT 61.590000 185.595000 61.790000 185.795000 ;
        RECT 61.590000 185.995000 61.790000 186.195000 ;
        RECT 61.590000 186.395000 61.790000 186.595000 ;
        RECT 61.590000 186.795000 61.790000 186.995000 ;
        RECT 61.590000 187.195000 61.790000 187.395000 ;
        RECT 61.590000 187.595000 61.790000 187.795000 ;
        RECT 61.590000 187.995000 61.790000 188.195000 ;
        RECT 61.590000 188.395000 61.790000 188.595000 ;
        RECT 61.590000 188.795000 61.790000 188.995000 ;
        RECT 61.590000 189.195000 61.790000 189.395000 ;
        RECT 61.590000 189.595000 61.790000 189.795000 ;
        RECT 61.590000 189.995000 61.790000 190.195000 ;
        RECT 61.590000 190.395000 61.790000 190.595000 ;
        RECT 61.590000 190.795000 61.790000 190.995000 ;
        RECT 61.590000 191.195000 61.790000 191.395000 ;
        RECT 61.590000 191.595000 61.790000 191.795000 ;
        RECT 61.590000 191.995000 61.790000 192.195000 ;
        RECT 61.590000 192.395000 61.790000 192.595000 ;
        RECT 61.590000 192.795000 61.790000 192.995000 ;
        RECT 61.590000 193.195000 61.790000 193.395000 ;
        RECT 61.590000 193.595000 61.790000 193.795000 ;
        RECT 61.590000 193.995000 61.790000 194.195000 ;
        RECT 61.590000 194.395000 61.790000 194.595000 ;
        RECT 61.590000 194.795000 61.790000 194.995000 ;
        RECT 61.590000 195.200000 61.790000 195.400000 ;
        RECT 61.590000 195.605000 61.790000 195.805000 ;
        RECT 61.590000 196.010000 61.790000 196.210000 ;
        RECT 61.590000 196.415000 61.790000 196.615000 ;
        RECT 61.590000 196.820000 61.790000 197.020000 ;
        RECT 61.590000 197.225000 61.790000 197.425000 ;
        RECT 61.590000 197.630000 61.790000 197.830000 ;
        RECT 61.590000 198.035000 61.790000 198.235000 ;
        RECT 61.590000 198.440000 61.790000 198.640000 ;
        RECT 61.590000 198.845000 61.790000 199.045000 ;
        RECT 61.590000 199.250000 61.790000 199.450000 ;
        RECT 61.590000 199.655000 61.790000 199.855000 ;
        RECT 61.850000  25.910000 62.050000  26.110000 ;
        RECT 61.850000  26.340000 62.050000  26.540000 ;
        RECT 61.850000  26.770000 62.050000  26.970000 ;
        RECT 61.850000  27.200000 62.050000  27.400000 ;
        RECT 61.850000  27.630000 62.050000  27.830000 ;
        RECT 61.850000  28.060000 62.050000  28.260000 ;
        RECT 61.850000  28.490000 62.050000  28.690000 ;
        RECT 61.850000  28.920000 62.050000  29.120000 ;
        RECT 61.850000  29.350000 62.050000  29.550000 ;
        RECT 61.850000  29.780000 62.050000  29.980000 ;
        RECT 61.850000  30.210000 62.050000  30.410000 ;
        RECT 61.990000 175.995000 62.190000 176.195000 ;
        RECT 61.990000 176.395000 62.190000 176.595000 ;
        RECT 61.990000 176.795000 62.190000 176.995000 ;
        RECT 61.990000 177.195000 62.190000 177.395000 ;
        RECT 61.990000 177.595000 62.190000 177.795000 ;
        RECT 61.990000 177.995000 62.190000 178.195000 ;
        RECT 61.990000 178.395000 62.190000 178.595000 ;
        RECT 61.990000 178.795000 62.190000 178.995000 ;
        RECT 61.990000 179.195000 62.190000 179.395000 ;
        RECT 61.990000 179.595000 62.190000 179.795000 ;
        RECT 61.990000 179.995000 62.190000 180.195000 ;
        RECT 61.990000 180.395000 62.190000 180.595000 ;
        RECT 61.990000 180.795000 62.190000 180.995000 ;
        RECT 61.990000 181.195000 62.190000 181.395000 ;
        RECT 61.990000 181.595000 62.190000 181.795000 ;
        RECT 61.990000 181.995000 62.190000 182.195000 ;
        RECT 61.990000 182.395000 62.190000 182.595000 ;
        RECT 61.990000 182.795000 62.190000 182.995000 ;
        RECT 61.990000 183.195000 62.190000 183.395000 ;
        RECT 61.990000 183.595000 62.190000 183.795000 ;
        RECT 61.990000 183.995000 62.190000 184.195000 ;
        RECT 61.990000 184.395000 62.190000 184.595000 ;
        RECT 61.990000 184.795000 62.190000 184.995000 ;
        RECT 61.990000 185.195000 62.190000 185.395000 ;
        RECT 61.990000 185.595000 62.190000 185.795000 ;
        RECT 61.990000 185.995000 62.190000 186.195000 ;
        RECT 61.990000 186.395000 62.190000 186.595000 ;
        RECT 61.990000 186.795000 62.190000 186.995000 ;
        RECT 61.990000 187.195000 62.190000 187.395000 ;
        RECT 61.990000 187.595000 62.190000 187.795000 ;
        RECT 61.990000 187.995000 62.190000 188.195000 ;
        RECT 61.990000 188.395000 62.190000 188.595000 ;
        RECT 61.990000 188.795000 62.190000 188.995000 ;
        RECT 61.990000 189.195000 62.190000 189.395000 ;
        RECT 61.990000 189.595000 62.190000 189.795000 ;
        RECT 61.990000 189.995000 62.190000 190.195000 ;
        RECT 61.990000 190.395000 62.190000 190.595000 ;
        RECT 61.990000 190.795000 62.190000 190.995000 ;
        RECT 61.990000 191.195000 62.190000 191.395000 ;
        RECT 61.990000 191.595000 62.190000 191.795000 ;
        RECT 61.990000 191.995000 62.190000 192.195000 ;
        RECT 61.990000 192.395000 62.190000 192.595000 ;
        RECT 61.990000 192.795000 62.190000 192.995000 ;
        RECT 61.990000 193.195000 62.190000 193.395000 ;
        RECT 61.990000 193.595000 62.190000 193.795000 ;
        RECT 61.990000 193.995000 62.190000 194.195000 ;
        RECT 61.990000 194.395000 62.190000 194.595000 ;
        RECT 61.990000 194.795000 62.190000 194.995000 ;
        RECT 61.990000 195.200000 62.190000 195.400000 ;
        RECT 61.990000 195.605000 62.190000 195.805000 ;
        RECT 61.990000 196.010000 62.190000 196.210000 ;
        RECT 61.990000 196.415000 62.190000 196.615000 ;
        RECT 61.990000 196.820000 62.190000 197.020000 ;
        RECT 61.990000 197.225000 62.190000 197.425000 ;
        RECT 61.990000 197.630000 62.190000 197.830000 ;
        RECT 61.990000 198.035000 62.190000 198.235000 ;
        RECT 61.990000 198.440000 62.190000 198.640000 ;
        RECT 61.990000 198.845000 62.190000 199.045000 ;
        RECT 61.990000 199.250000 62.190000 199.450000 ;
        RECT 61.990000 199.655000 62.190000 199.855000 ;
        RECT 62.255000  25.910000 62.455000  26.110000 ;
        RECT 62.255000  26.340000 62.455000  26.540000 ;
        RECT 62.255000  26.770000 62.455000  26.970000 ;
        RECT 62.255000  27.200000 62.455000  27.400000 ;
        RECT 62.255000  27.630000 62.455000  27.830000 ;
        RECT 62.255000  28.060000 62.455000  28.260000 ;
        RECT 62.255000  28.490000 62.455000  28.690000 ;
        RECT 62.255000  28.920000 62.455000  29.120000 ;
        RECT 62.255000  29.350000 62.455000  29.550000 ;
        RECT 62.255000  29.780000 62.455000  29.980000 ;
        RECT 62.255000  30.210000 62.455000  30.410000 ;
        RECT 62.390000 175.995000 62.590000 176.195000 ;
        RECT 62.390000 176.395000 62.590000 176.595000 ;
        RECT 62.390000 176.795000 62.590000 176.995000 ;
        RECT 62.390000 177.195000 62.590000 177.395000 ;
        RECT 62.390000 177.595000 62.590000 177.795000 ;
        RECT 62.390000 177.995000 62.590000 178.195000 ;
        RECT 62.390000 178.395000 62.590000 178.595000 ;
        RECT 62.390000 178.795000 62.590000 178.995000 ;
        RECT 62.390000 179.195000 62.590000 179.395000 ;
        RECT 62.390000 179.595000 62.590000 179.795000 ;
        RECT 62.390000 179.995000 62.590000 180.195000 ;
        RECT 62.390000 180.395000 62.590000 180.595000 ;
        RECT 62.390000 180.795000 62.590000 180.995000 ;
        RECT 62.390000 181.195000 62.590000 181.395000 ;
        RECT 62.390000 181.595000 62.590000 181.795000 ;
        RECT 62.390000 181.995000 62.590000 182.195000 ;
        RECT 62.390000 182.395000 62.590000 182.595000 ;
        RECT 62.390000 182.795000 62.590000 182.995000 ;
        RECT 62.390000 183.195000 62.590000 183.395000 ;
        RECT 62.390000 183.595000 62.590000 183.795000 ;
        RECT 62.390000 183.995000 62.590000 184.195000 ;
        RECT 62.390000 184.395000 62.590000 184.595000 ;
        RECT 62.390000 184.795000 62.590000 184.995000 ;
        RECT 62.390000 185.195000 62.590000 185.395000 ;
        RECT 62.390000 185.595000 62.590000 185.795000 ;
        RECT 62.390000 185.995000 62.590000 186.195000 ;
        RECT 62.390000 186.395000 62.590000 186.595000 ;
        RECT 62.390000 186.795000 62.590000 186.995000 ;
        RECT 62.390000 187.195000 62.590000 187.395000 ;
        RECT 62.390000 187.595000 62.590000 187.795000 ;
        RECT 62.390000 187.995000 62.590000 188.195000 ;
        RECT 62.390000 188.395000 62.590000 188.595000 ;
        RECT 62.390000 188.795000 62.590000 188.995000 ;
        RECT 62.390000 189.195000 62.590000 189.395000 ;
        RECT 62.390000 189.595000 62.590000 189.795000 ;
        RECT 62.390000 189.995000 62.590000 190.195000 ;
        RECT 62.390000 190.395000 62.590000 190.595000 ;
        RECT 62.390000 190.795000 62.590000 190.995000 ;
        RECT 62.390000 191.195000 62.590000 191.395000 ;
        RECT 62.390000 191.595000 62.590000 191.795000 ;
        RECT 62.390000 191.995000 62.590000 192.195000 ;
        RECT 62.390000 192.395000 62.590000 192.595000 ;
        RECT 62.390000 192.795000 62.590000 192.995000 ;
        RECT 62.390000 193.195000 62.590000 193.395000 ;
        RECT 62.390000 193.595000 62.590000 193.795000 ;
        RECT 62.390000 193.995000 62.590000 194.195000 ;
        RECT 62.390000 194.395000 62.590000 194.595000 ;
        RECT 62.390000 194.795000 62.590000 194.995000 ;
        RECT 62.390000 195.200000 62.590000 195.400000 ;
        RECT 62.390000 195.605000 62.590000 195.805000 ;
        RECT 62.390000 196.010000 62.590000 196.210000 ;
        RECT 62.390000 196.415000 62.590000 196.615000 ;
        RECT 62.390000 196.820000 62.590000 197.020000 ;
        RECT 62.390000 197.225000 62.590000 197.425000 ;
        RECT 62.390000 197.630000 62.590000 197.830000 ;
        RECT 62.390000 198.035000 62.590000 198.235000 ;
        RECT 62.390000 198.440000 62.590000 198.640000 ;
        RECT 62.390000 198.845000 62.590000 199.045000 ;
        RECT 62.390000 199.250000 62.590000 199.450000 ;
        RECT 62.390000 199.655000 62.590000 199.855000 ;
        RECT 62.660000  25.910000 62.860000  26.110000 ;
        RECT 62.660000  26.340000 62.860000  26.540000 ;
        RECT 62.660000  26.770000 62.860000  26.970000 ;
        RECT 62.660000  27.200000 62.860000  27.400000 ;
        RECT 62.660000  27.630000 62.860000  27.830000 ;
        RECT 62.660000  28.060000 62.860000  28.260000 ;
        RECT 62.660000  28.490000 62.860000  28.690000 ;
        RECT 62.660000  28.920000 62.860000  29.120000 ;
        RECT 62.660000  29.350000 62.860000  29.550000 ;
        RECT 62.660000  29.780000 62.860000  29.980000 ;
        RECT 62.660000  30.210000 62.860000  30.410000 ;
        RECT 62.790000 175.995000 62.990000 176.195000 ;
        RECT 62.790000 176.395000 62.990000 176.595000 ;
        RECT 62.790000 176.795000 62.990000 176.995000 ;
        RECT 62.790000 177.195000 62.990000 177.395000 ;
        RECT 62.790000 177.595000 62.990000 177.795000 ;
        RECT 62.790000 177.995000 62.990000 178.195000 ;
        RECT 62.790000 178.395000 62.990000 178.595000 ;
        RECT 62.790000 178.795000 62.990000 178.995000 ;
        RECT 62.790000 179.195000 62.990000 179.395000 ;
        RECT 62.790000 179.595000 62.990000 179.795000 ;
        RECT 62.790000 179.995000 62.990000 180.195000 ;
        RECT 62.790000 180.395000 62.990000 180.595000 ;
        RECT 62.790000 180.795000 62.990000 180.995000 ;
        RECT 62.790000 181.195000 62.990000 181.395000 ;
        RECT 62.790000 181.595000 62.990000 181.795000 ;
        RECT 62.790000 181.995000 62.990000 182.195000 ;
        RECT 62.790000 182.395000 62.990000 182.595000 ;
        RECT 62.790000 182.795000 62.990000 182.995000 ;
        RECT 62.790000 183.195000 62.990000 183.395000 ;
        RECT 62.790000 183.595000 62.990000 183.795000 ;
        RECT 62.790000 183.995000 62.990000 184.195000 ;
        RECT 62.790000 184.395000 62.990000 184.595000 ;
        RECT 62.790000 184.795000 62.990000 184.995000 ;
        RECT 62.790000 185.195000 62.990000 185.395000 ;
        RECT 62.790000 185.595000 62.990000 185.795000 ;
        RECT 62.790000 185.995000 62.990000 186.195000 ;
        RECT 62.790000 186.395000 62.990000 186.595000 ;
        RECT 62.790000 186.795000 62.990000 186.995000 ;
        RECT 62.790000 187.195000 62.990000 187.395000 ;
        RECT 62.790000 187.595000 62.990000 187.795000 ;
        RECT 62.790000 187.995000 62.990000 188.195000 ;
        RECT 62.790000 188.395000 62.990000 188.595000 ;
        RECT 62.790000 188.795000 62.990000 188.995000 ;
        RECT 62.790000 189.195000 62.990000 189.395000 ;
        RECT 62.790000 189.595000 62.990000 189.795000 ;
        RECT 62.790000 189.995000 62.990000 190.195000 ;
        RECT 62.790000 190.395000 62.990000 190.595000 ;
        RECT 62.790000 190.795000 62.990000 190.995000 ;
        RECT 62.790000 191.195000 62.990000 191.395000 ;
        RECT 62.790000 191.595000 62.990000 191.795000 ;
        RECT 62.790000 191.995000 62.990000 192.195000 ;
        RECT 62.790000 192.395000 62.990000 192.595000 ;
        RECT 62.790000 192.795000 62.990000 192.995000 ;
        RECT 62.790000 193.195000 62.990000 193.395000 ;
        RECT 62.790000 193.595000 62.990000 193.795000 ;
        RECT 62.790000 193.995000 62.990000 194.195000 ;
        RECT 62.790000 194.395000 62.990000 194.595000 ;
        RECT 62.790000 194.795000 62.990000 194.995000 ;
        RECT 62.790000 195.200000 62.990000 195.400000 ;
        RECT 62.790000 195.605000 62.990000 195.805000 ;
        RECT 62.790000 196.010000 62.990000 196.210000 ;
        RECT 62.790000 196.415000 62.990000 196.615000 ;
        RECT 62.790000 196.820000 62.990000 197.020000 ;
        RECT 62.790000 197.225000 62.990000 197.425000 ;
        RECT 62.790000 197.630000 62.990000 197.830000 ;
        RECT 62.790000 198.035000 62.990000 198.235000 ;
        RECT 62.790000 198.440000 62.990000 198.640000 ;
        RECT 62.790000 198.845000 62.990000 199.045000 ;
        RECT 62.790000 199.250000 62.990000 199.450000 ;
        RECT 62.790000 199.655000 62.990000 199.855000 ;
        RECT 63.065000  25.910000 63.265000  26.110000 ;
        RECT 63.065000  26.340000 63.265000  26.540000 ;
        RECT 63.065000  26.770000 63.265000  26.970000 ;
        RECT 63.065000  27.200000 63.265000  27.400000 ;
        RECT 63.065000  27.630000 63.265000  27.830000 ;
        RECT 63.065000  28.060000 63.265000  28.260000 ;
        RECT 63.065000  28.490000 63.265000  28.690000 ;
        RECT 63.065000  28.920000 63.265000  29.120000 ;
        RECT 63.065000  29.350000 63.265000  29.550000 ;
        RECT 63.065000  29.780000 63.265000  29.980000 ;
        RECT 63.065000  30.210000 63.265000  30.410000 ;
        RECT 63.190000 175.995000 63.390000 176.195000 ;
        RECT 63.190000 176.395000 63.390000 176.595000 ;
        RECT 63.190000 176.795000 63.390000 176.995000 ;
        RECT 63.190000 177.195000 63.390000 177.395000 ;
        RECT 63.190000 177.595000 63.390000 177.795000 ;
        RECT 63.190000 177.995000 63.390000 178.195000 ;
        RECT 63.190000 178.395000 63.390000 178.595000 ;
        RECT 63.190000 178.795000 63.390000 178.995000 ;
        RECT 63.190000 179.195000 63.390000 179.395000 ;
        RECT 63.190000 179.595000 63.390000 179.795000 ;
        RECT 63.190000 179.995000 63.390000 180.195000 ;
        RECT 63.190000 180.395000 63.390000 180.595000 ;
        RECT 63.190000 180.795000 63.390000 180.995000 ;
        RECT 63.190000 181.195000 63.390000 181.395000 ;
        RECT 63.190000 181.595000 63.390000 181.795000 ;
        RECT 63.190000 181.995000 63.390000 182.195000 ;
        RECT 63.190000 182.395000 63.390000 182.595000 ;
        RECT 63.190000 182.795000 63.390000 182.995000 ;
        RECT 63.190000 183.195000 63.390000 183.395000 ;
        RECT 63.190000 183.595000 63.390000 183.795000 ;
        RECT 63.190000 183.995000 63.390000 184.195000 ;
        RECT 63.190000 184.395000 63.390000 184.595000 ;
        RECT 63.190000 184.795000 63.390000 184.995000 ;
        RECT 63.190000 185.195000 63.390000 185.395000 ;
        RECT 63.190000 185.595000 63.390000 185.795000 ;
        RECT 63.190000 185.995000 63.390000 186.195000 ;
        RECT 63.190000 186.395000 63.390000 186.595000 ;
        RECT 63.190000 186.795000 63.390000 186.995000 ;
        RECT 63.190000 187.195000 63.390000 187.395000 ;
        RECT 63.190000 187.595000 63.390000 187.795000 ;
        RECT 63.190000 187.995000 63.390000 188.195000 ;
        RECT 63.190000 188.395000 63.390000 188.595000 ;
        RECT 63.190000 188.795000 63.390000 188.995000 ;
        RECT 63.190000 189.195000 63.390000 189.395000 ;
        RECT 63.190000 189.595000 63.390000 189.795000 ;
        RECT 63.190000 189.995000 63.390000 190.195000 ;
        RECT 63.190000 190.395000 63.390000 190.595000 ;
        RECT 63.190000 190.795000 63.390000 190.995000 ;
        RECT 63.190000 191.195000 63.390000 191.395000 ;
        RECT 63.190000 191.595000 63.390000 191.795000 ;
        RECT 63.190000 191.995000 63.390000 192.195000 ;
        RECT 63.190000 192.395000 63.390000 192.595000 ;
        RECT 63.190000 192.795000 63.390000 192.995000 ;
        RECT 63.190000 193.195000 63.390000 193.395000 ;
        RECT 63.190000 193.595000 63.390000 193.795000 ;
        RECT 63.190000 193.995000 63.390000 194.195000 ;
        RECT 63.190000 194.395000 63.390000 194.595000 ;
        RECT 63.190000 194.795000 63.390000 194.995000 ;
        RECT 63.190000 195.200000 63.390000 195.400000 ;
        RECT 63.190000 195.605000 63.390000 195.805000 ;
        RECT 63.190000 196.010000 63.390000 196.210000 ;
        RECT 63.190000 196.415000 63.390000 196.615000 ;
        RECT 63.190000 196.820000 63.390000 197.020000 ;
        RECT 63.190000 197.225000 63.390000 197.425000 ;
        RECT 63.190000 197.630000 63.390000 197.830000 ;
        RECT 63.190000 198.035000 63.390000 198.235000 ;
        RECT 63.190000 198.440000 63.390000 198.640000 ;
        RECT 63.190000 198.845000 63.390000 199.045000 ;
        RECT 63.190000 199.250000 63.390000 199.450000 ;
        RECT 63.190000 199.655000 63.390000 199.855000 ;
        RECT 63.470000  25.910000 63.670000  26.110000 ;
        RECT 63.470000  26.340000 63.670000  26.540000 ;
        RECT 63.470000  26.770000 63.670000  26.970000 ;
        RECT 63.470000  27.200000 63.670000  27.400000 ;
        RECT 63.470000  27.630000 63.670000  27.830000 ;
        RECT 63.470000  28.060000 63.670000  28.260000 ;
        RECT 63.470000  28.490000 63.670000  28.690000 ;
        RECT 63.470000  28.920000 63.670000  29.120000 ;
        RECT 63.470000  29.350000 63.670000  29.550000 ;
        RECT 63.470000  29.780000 63.670000  29.980000 ;
        RECT 63.470000  30.210000 63.670000  30.410000 ;
        RECT 63.590000 175.995000 63.790000 176.195000 ;
        RECT 63.590000 176.395000 63.790000 176.595000 ;
        RECT 63.590000 176.795000 63.790000 176.995000 ;
        RECT 63.590000 177.195000 63.790000 177.395000 ;
        RECT 63.590000 177.595000 63.790000 177.795000 ;
        RECT 63.590000 177.995000 63.790000 178.195000 ;
        RECT 63.590000 178.395000 63.790000 178.595000 ;
        RECT 63.590000 178.795000 63.790000 178.995000 ;
        RECT 63.590000 179.195000 63.790000 179.395000 ;
        RECT 63.590000 179.595000 63.790000 179.795000 ;
        RECT 63.590000 179.995000 63.790000 180.195000 ;
        RECT 63.590000 180.395000 63.790000 180.595000 ;
        RECT 63.590000 180.795000 63.790000 180.995000 ;
        RECT 63.590000 181.195000 63.790000 181.395000 ;
        RECT 63.590000 181.595000 63.790000 181.795000 ;
        RECT 63.590000 181.995000 63.790000 182.195000 ;
        RECT 63.590000 182.395000 63.790000 182.595000 ;
        RECT 63.590000 182.795000 63.790000 182.995000 ;
        RECT 63.590000 183.195000 63.790000 183.395000 ;
        RECT 63.590000 183.595000 63.790000 183.795000 ;
        RECT 63.590000 183.995000 63.790000 184.195000 ;
        RECT 63.590000 184.395000 63.790000 184.595000 ;
        RECT 63.590000 184.795000 63.790000 184.995000 ;
        RECT 63.590000 185.195000 63.790000 185.395000 ;
        RECT 63.590000 185.595000 63.790000 185.795000 ;
        RECT 63.590000 185.995000 63.790000 186.195000 ;
        RECT 63.590000 186.395000 63.790000 186.595000 ;
        RECT 63.590000 186.795000 63.790000 186.995000 ;
        RECT 63.590000 187.195000 63.790000 187.395000 ;
        RECT 63.590000 187.595000 63.790000 187.795000 ;
        RECT 63.590000 187.995000 63.790000 188.195000 ;
        RECT 63.590000 188.395000 63.790000 188.595000 ;
        RECT 63.590000 188.795000 63.790000 188.995000 ;
        RECT 63.590000 189.195000 63.790000 189.395000 ;
        RECT 63.590000 189.595000 63.790000 189.795000 ;
        RECT 63.590000 189.995000 63.790000 190.195000 ;
        RECT 63.590000 190.395000 63.790000 190.595000 ;
        RECT 63.590000 190.795000 63.790000 190.995000 ;
        RECT 63.590000 191.195000 63.790000 191.395000 ;
        RECT 63.590000 191.595000 63.790000 191.795000 ;
        RECT 63.590000 191.995000 63.790000 192.195000 ;
        RECT 63.590000 192.395000 63.790000 192.595000 ;
        RECT 63.590000 192.795000 63.790000 192.995000 ;
        RECT 63.590000 193.195000 63.790000 193.395000 ;
        RECT 63.590000 193.595000 63.790000 193.795000 ;
        RECT 63.590000 193.995000 63.790000 194.195000 ;
        RECT 63.590000 194.395000 63.790000 194.595000 ;
        RECT 63.590000 194.795000 63.790000 194.995000 ;
        RECT 63.590000 195.200000 63.790000 195.400000 ;
        RECT 63.590000 195.605000 63.790000 195.805000 ;
        RECT 63.590000 196.010000 63.790000 196.210000 ;
        RECT 63.590000 196.415000 63.790000 196.615000 ;
        RECT 63.590000 196.820000 63.790000 197.020000 ;
        RECT 63.590000 197.225000 63.790000 197.425000 ;
        RECT 63.590000 197.630000 63.790000 197.830000 ;
        RECT 63.590000 198.035000 63.790000 198.235000 ;
        RECT 63.590000 198.440000 63.790000 198.640000 ;
        RECT 63.590000 198.845000 63.790000 199.045000 ;
        RECT 63.590000 199.250000 63.790000 199.450000 ;
        RECT 63.590000 199.655000 63.790000 199.855000 ;
        RECT 63.875000  25.910000 64.075000  26.110000 ;
        RECT 63.875000  26.340000 64.075000  26.540000 ;
        RECT 63.875000  26.770000 64.075000  26.970000 ;
        RECT 63.875000  27.200000 64.075000  27.400000 ;
        RECT 63.875000  27.630000 64.075000  27.830000 ;
        RECT 63.875000  28.060000 64.075000  28.260000 ;
        RECT 63.875000  28.490000 64.075000  28.690000 ;
        RECT 63.875000  28.920000 64.075000  29.120000 ;
        RECT 63.875000  29.350000 64.075000  29.550000 ;
        RECT 63.875000  29.780000 64.075000  29.980000 ;
        RECT 63.875000  30.210000 64.075000  30.410000 ;
        RECT 63.990000 175.995000 64.190000 176.195000 ;
        RECT 63.990000 176.395000 64.190000 176.595000 ;
        RECT 63.990000 176.795000 64.190000 176.995000 ;
        RECT 63.990000 177.195000 64.190000 177.395000 ;
        RECT 63.990000 177.595000 64.190000 177.795000 ;
        RECT 63.990000 177.995000 64.190000 178.195000 ;
        RECT 63.990000 178.395000 64.190000 178.595000 ;
        RECT 63.990000 178.795000 64.190000 178.995000 ;
        RECT 63.990000 179.195000 64.190000 179.395000 ;
        RECT 63.990000 179.595000 64.190000 179.795000 ;
        RECT 63.990000 179.995000 64.190000 180.195000 ;
        RECT 63.990000 180.395000 64.190000 180.595000 ;
        RECT 63.990000 180.795000 64.190000 180.995000 ;
        RECT 63.990000 181.195000 64.190000 181.395000 ;
        RECT 63.990000 181.595000 64.190000 181.795000 ;
        RECT 63.990000 181.995000 64.190000 182.195000 ;
        RECT 63.990000 182.395000 64.190000 182.595000 ;
        RECT 63.990000 182.795000 64.190000 182.995000 ;
        RECT 63.990000 183.195000 64.190000 183.395000 ;
        RECT 63.990000 183.595000 64.190000 183.795000 ;
        RECT 63.990000 183.995000 64.190000 184.195000 ;
        RECT 63.990000 184.395000 64.190000 184.595000 ;
        RECT 63.990000 184.795000 64.190000 184.995000 ;
        RECT 63.990000 185.195000 64.190000 185.395000 ;
        RECT 63.990000 185.595000 64.190000 185.795000 ;
        RECT 63.990000 185.995000 64.190000 186.195000 ;
        RECT 63.990000 186.395000 64.190000 186.595000 ;
        RECT 63.990000 186.795000 64.190000 186.995000 ;
        RECT 63.990000 187.195000 64.190000 187.395000 ;
        RECT 63.990000 187.595000 64.190000 187.795000 ;
        RECT 63.990000 187.995000 64.190000 188.195000 ;
        RECT 63.990000 188.395000 64.190000 188.595000 ;
        RECT 63.990000 188.795000 64.190000 188.995000 ;
        RECT 63.990000 189.195000 64.190000 189.395000 ;
        RECT 63.990000 189.595000 64.190000 189.795000 ;
        RECT 63.990000 189.995000 64.190000 190.195000 ;
        RECT 63.990000 190.395000 64.190000 190.595000 ;
        RECT 63.990000 190.795000 64.190000 190.995000 ;
        RECT 63.990000 191.195000 64.190000 191.395000 ;
        RECT 63.990000 191.595000 64.190000 191.795000 ;
        RECT 63.990000 191.995000 64.190000 192.195000 ;
        RECT 63.990000 192.395000 64.190000 192.595000 ;
        RECT 63.990000 192.795000 64.190000 192.995000 ;
        RECT 63.990000 193.195000 64.190000 193.395000 ;
        RECT 63.990000 193.595000 64.190000 193.795000 ;
        RECT 63.990000 193.995000 64.190000 194.195000 ;
        RECT 63.990000 194.395000 64.190000 194.595000 ;
        RECT 63.990000 194.795000 64.190000 194.995000 ;
        RECT 63.990000 195.200000 64.190000 195.400000 ;
        RECT 63.990000 195.605000 64.190000 195.805000 ;
        RECT 63.990000 196.010000 64.190000 196.210000 ;
        RECT 63.990000 196.415000 64.190000 196.615000 ;
        RECT 63.990000 196.820000 64.190000 197.020000 ;
        RECT 63.990000 197.225000 64.190000 197.425000 ;
        RECT 63.990000 197.630000 64.190000 197.830000 ;
        RECT 63.990000 198.035000 64.190000 198.235000 ;
        RECT 63.990000 198.440000 64.190000 198.640000 ;
        RECT 63.990000 198.845000 64.190000 199.045000 ;
        RECT 63.990000 199.250000 64.190000 199.450000 ;
        RECT 63.990000 199.655000 64.190000 199.855000 ;
        RECT 64.280000  25.910000 64.480000  26.110000 ;
        RECT 64.280000  26.340000 64.480000  26.540000 ;
        RECT 64.280000  26.770000 64.480000  26.970000 ;
        RECT 64.280000  27.200000 64.480000  27.400000 ;
        RECT 64.280000  27.630000 64.480000  27.830000 ;
        RECT 64.280000  28.060000 64.480000  28.260000 ;
        RECT 64.280000  28.490000 64.480000  28.690000 ;
        RECT 64.280000  28.920000 64.480000  29.120000 ;
        RECT 64.280000  29.350000 64.480000  29.550000 ;
        RECT 64.280000  29.780000 64.480000  29.980000 ;
        RECT 64.280000  30.210000 64.480000  30.410000 ;
        RECT 64.390000 175.995000 64.590000 176.195000 ;
        RECT 64.390000 176.395000 64.590000 176.595000 ;
        RECT 64.390000 176.795000 64.590000 176.995000 ;
        RECT 64.390000 177.195000 64.590000 177.395000 ;
        RECT 64.390000 177.595000 64.590000 177.795000 ;
        RECT 64.390000 177.995000 64.590000 178.195000 ;
        RECT 64.390000 178.395000 64.590000 178.595000 ;
        RECT 64.390000 178.795000 64.590000 178.995000 ;
        RECT 64.390000 179.195000 64.590000 179.395000 ;
        RECT 64.390000 179.595000 64.590000 179.795000 ;
        RECT 64.390000 179.995000 64.590000 180.195000 ;
        RECT 64.390000 180.395000 64.590000 180.595000 ;
        RECT 64.390000 180.795000 64.590000 180.995000 ;
        RECT 64.390000 181.195000 64.590000 181.395000 ;
        RECT 64.390000 181.595000 64.590000 181.795000 ;
        RECT 64.390000 181.995000 64.590000 182.195000 ;
        RECT 64.390000 182.395000 64.590000 182.595000 ;
        RECT 64.390000 182.795000 64.590000 182.995000 ;
        RECT 64.390000 183.195000 64.590000 183.395000 ;
        RECT 64.390000 183.595000 64.590000 183.795000 ;
        RECT 64.390000 183.995000 64.590000 184.195000 ;
        RECT 64.390000 184.395000 64.590000 184.595000 ;
        RECT 64.390000 184.795000 64.590000 184.995000 ;
        RECT 64.390000 185.195000 64.590000 185.395000 ;
        RECT 64.390000 185.595000 64.590000 185.795000 ;
        RECT 64.390000 185.995000 64.590000 186.195000 ;
        RECT 64.390000 186.395000 64.590000 186.595000 ;
        RECT 64.390000 186.795000 64.590000 186.995000 ;
        RECT 64.390000 187.195000 64.590000 187.395000 ;
        RECT 64.390000 187.595000 64.590000 187.795000 ;
        RECT 64.390000 187.995000 64.590000 188.195000 ;
        RECT 64.390000 188.395000 64.590000 188.595000 ;
        RECT 64.390000 188.795000 64.590000 188.995000 ;
        RECT 64.390000 189.195000 64.590000 189.395000 ;
        RECT 64.390000 189.595000 64.590000 189.795000 ;
        RECT 64.390000 189.995000 64.590000 190.195000 ;
        RECT 64.390000 190.395000 64.590000 190.595000 ;
        RECT 64.390000 190.795000 64.590000 190.995000 ;
        RECT 64.390000 191.195000 64.590000 191.395000 ;
        RECT 64.390000 191.595000 64.590000 191.795000 ;
        RECT 64.390000 191.995000 64.590000 192.195000 ;
        RECT 64.390000 192.395000 64.590000 192.595000 ;
        RECT 64.390000 192.795000 64.590000 192.995000 ;
        RECT 64.390000 193.195000 64.590000 193.395000 ;
        RECT 64.390000 193.595000 64.590000 193.795000 ;
        RECT 64.390000 193.995000 64.590000 194.195000 ;
        RECT 64.390000 194.395000 64.590000 194.595000 ;
        RECT 64.390000 194.795000 64.590000 194.995000 ;
        RECT 64.390000 195.200000 64.590000 195.400000 ;
        RECT 64.390000 195.605000 64.590000 195.805000 ;
        RECT 64.390000 196.010000 64.590000 196.210000 ;
        RECT 64.390000 196.415000 64.590000 196.615000 ;
        RECT 64.390000 196.820000 64.590000 197.020000 ;
        RECT 64.390000 197.225000 64.590000 197.425000 ;
        RECT 64.390000 197.630000 64.590000 197.830000 ;
        RECT 64.390000 198.035000 64.590000 198.235000 ;
        RECT 64.390000 198.440000 64.590000 198.640000 ;
        RECT 64.390000 198.845000 64.590000 199.045000 ;
        RECT 64.390000 199.250000 64.590000 199.450000 ;
        RECT 64.390000 199.655000 64.590000 199.855000 ;
        RECT 64.685000  25.910000 64.885000  26.110000 ;
        RECT 64.685000  26.340000 64.885000  26.540000 ;
        RECT 64.685000  26.770000 64.885000  26.970000 ;
        RECT 64.685000  27.200000 64.885000  27.400000 ;
        RECT 64.685000  27.630000 64.885000  27.830000 ;
        RECT 64.685000  28.060000 64.885000  28.260000 ;
        RECT 64.685000  28.490000 64.885000  28.690000 ;
        RECT 64.685000  28.920000 64.885000  29.120000 ;
        RECT 64.685000  29.350000 64.885000  29.550000 ;
        RECT 64.685000  29.780000 64.885000  29.980000 ;
        RECT 64.685000  30.210000 64.885000  30.410000 ;
        RECT 64.790000 175.995000 64.990000 176.195000 ;
        RECT 64.790000 176.395000 64.990000 176.595000 ;
        RECT 64.790000 176.795000 64.990000 176.995000 ;
        RECT 64.790000 177.195000 64.990000 177.395000 ;
        RECT 64.790000 177.595000 64.990000 177.795000 ;
        RECT 64.790000 177.995000 64.990000 178.195000 ;
        RECT 64.790000 178.395000 64.990000 178.595000 ;
        RECT 64.790000 178.795000 64.990000 178.995000 ;
        RECT 64.790000 179.195000 64.990000 179.395000 ;
        RECT 64.790000 179.595000 64.990000 179.795000 ;
        RECT 64.790000 179.995000 64.990000 180.195000 ;
        RECT 64.790000 180.395000 64.990000 180.595000 ;
        RECT 64.790000 180.795000 64.990000 180.995000 ;
        RECT 64.790000 181.195000 64.990000 181.395000 ;
        RECT 64.790000 181.595000 64.990000 181.795000 ;
        RECT 64.790000 181.995000 64.990000 182.195000 ;
        RECT 64.790000 182.395000 64.990000 182.595000 ;
        RECT 64.790000 182.795000 64.990000 182.995000 ;
        RECT 64.790000 183.195000 64.990000 183.395000 ;
        RECT 64.790000 183.595000 64.990000 183.795000 ;
        RECT 64.790000 183.995000 64.990000 184.195000 ;
        RECT 64.790000 184.395000 64.990000 184.595000 ;
        RECT 64.790000 184.795000 64.990000 184.995000 ;
        RECT 64.790000 185.195000 64.990000 185.395000 ;
        RECT 64.790000 185.595000 64.990000 185.795000 ;
        RECT 64.790000 185.995000 64.990000 186.195000 ;
        RECT 64.790000 186.395000 64.990000 186.595000 ;
        RECT 64.790000 186.795000 64.990000 186.995000 ;
        RECT 64.790000 187.195000 64.990000 187.395000 ;
        RECT 64.790000 187.595000 64.990000 187.795000 ;
        RECT 64.790000 187.995000 64.990000 188.195000 ;
        RECT 64.790000 188.395000 64.990000 188.595000 ;
        RECT 64.790000 188.795000 64.990000 188.995000 ;
        RECT 64.790000 189.195000 64.990000 189.395000 ;
        RECT 64.790000 189.595000 64.990000 189.795000 ;
        RECT 64.790000 189.995000 64.990000 190.195000 ;
        RECT 64.790000 190.395000 64.990000 190.595000 ;
        RECT 64.790000 190.795000 64.990000 190.995000 ;
        RECT 64.790000 191.195000 64.990000 191.395000 ;
        RECT 64.790000 191.595000 64.990000 191.795000 ;
        RECT 64.790000 191.995000 64.990000 192.195000 ;
        RECT 64.790000 192.395000 64.990000 192.595000 ;
        RECT 64.790000 192.795000 64.990000 192.995000 ;
        RECT 64.790000 193.195000 64.990000 193.395000 ;
        RECT 64.790000 193.595000 64.990000 193.795000 ;
        RECT 64.790000 193.995000 64.990000 194.195000 ;
        RECT 64.790000 194.395000 64.990000 194.595000 ;
        RECT 64.790000 194.795000 64.990000 194.995000 ;
        RECT 64.790000 195.200000 64.990000 195.400000 ;
        RECT 64.790000 195.605000 64.990000 195.805000 ;
        RECT 64.790000 196.010000 64.990000 196.210000 ;
        RECT 64.790000 196.415000 64.990000 196.615000 ;
        RECT 64.790000 196.820000 64.990000 197.020000 ;
        RECT 64.790000 197.225000 64.990000 197.425000 ;
        RECT 64.790000 197.630000 64.990000 197.830000 ;
        RECT 64.790000 198.035000 64.990000 198.235000 ;
        RECT 64.790000 198.440000 64.990000 198.640000 ;
        RECT 64.790000 198.845000 64.990000 199.045000 ;
        RECT 64.790000 199.250000 64.990000 199.450000 ;
        RECT 64.790000 199.655000 64.990000 199.855000 ;
        RECT 65.090000  25.910000 65.290000  26.110000 ;
        RECT 65.090000  26.340000 65.290000  26.540000 ;
        RECT 65.090000  26.770000 65.290000  26.970000 ;
        RECT 65.090000  27.200000 65.290000  27.400000 ;
        RECT 65.090000  27.630000 65.290000  27.830000 ;
        RECT 65.090000  28.060000 65.290000  28.260000 ;
        RECT 65.090000  28.490000 65.290000  28.690000 ;
        RECT 65.090000  28.920000 65.290000  29.120000 ;
        RECT 65.090000  29.350000 65.290000  29.550000 ;
        RECT 65.090000  29.780000 65.290000  29.980000 ;
        RECT 65.090000  30.210000 65.290000  30.410000 ;
        RECT 65.190000 175.995000 65.390000 176.195000 ;
        RECT 65.190000 176.395000 65.390000 176.595000 ;
        RECT 65.190000 176.795000 65.390000 176.995000 ;
        RECT 65.190000 177.195000 65.390000 177.395000 ;
        RECT 65.190000 177.595000 65.390000 177.795000 ;
        RECT 65.190000 177.995000 65.390000 178.195000 ;
        RECT 65.190000 178.395000 65.390000 178.595000 ;
        RECT 65.190000 178.795000 65.390000 178.995000 ;
        RECT 65.190000 179.195000 65.390000 179.395000 ;
        RECT 65.190000 179.595000 65.390000 179.795000 ;
        RECT 65.190000 179.995000 65.390000 180.195000 ;
        RECT 65.190000 180.395000 65.390000 180.595000 ;
        RECT 65.190000 180.795000 65.390000 180.995000 ;
        RECT 65.190000 181.195000 65.390000 181.395000 ;
        RECT 65.190000 181.595000 65.390000 181.795000 ;
        RECT 65.190000 181.995000 65.390000 182.195000 ;
        RECT 65.190000 182.395000 65.390000 182.595000 ;
        RECT 65.190000 182.795000 65.390000 182.995000 ;
        RECT 65.190000 183.195000 65.390000 183.395000 ;
        RECT 65.190000 183.595000 65.390000 183.795000 ;
        RECT 65.190000 183.995000 65.390000 184.195000 ;
        RECT 65.190000 184.395000 65.390000 184.595000 ;
        RECT 65.190000 184.795000 65.390000 184.995000 ;
        RECT 65.190000 185.195000 65.390000 185.395000 ;
        RECT 65.190000 185.595000 65.390000 185.795000 ;
        RECT 65.190000 185.995000 65.390000 186.195000 ;
        RECT 65.190000 186.395000 65.390000 186.595000 ;
        RECT 65.190000 186.795000 65.390000 186.995000 ;
        RECT 65.190000 187.195000 65.390000 187.395000 ;
        RECT 65.190000 187.595000 65.390000 187.795000 ;
        RECT 65.190000 187.995000 65.390000 188.195000 ;
        RECT 65.190000 188.395000 65.390000 188.595000 ;
        RECT 65.190000 188.795000 65.390000 188.995000 ;
        RECT 65.190000 189.195000 65.390000 189.395000 ;
        RECT 65.190000 189.595000 65.390000 189.795000 ;
        RECT 65.190000 189.995000 65.390000 190.195000 ;
        RECT 65.190000 190.395000 65.390000 190.595000 ;
        RECT 65.190000 190.795000 65.390000 190.995000 ;
        RECT 65.190000 191.195000 65.390000 191.395000 ;
        RECT 65.190000 191.595000 65.390000 191.795000 ;
        RECT 65.190000 191.995000 65.390000 192.195000 ;
        RECT 65.190000 192.395000 65.390000 192.595000 ;
        RECT 65.190000 192.795000 65.390000 192.995000 ;
        RECT 65.190000 193.195000 65.390000 193.395000 ;
        RECT 65.190000 193.595000 65.390000 193.795000 ;
        RECT 65.190000 193.995000 65.390000 194.195000 ;
        RECT 65.190000 194.395000 65.390000 194.595000 ;
        RECT 65.190000 194.795000 65.390000 194.995000 ;
        RECT 65.190000 195.200000 65.390000 195.400000 ;
        RECT 65.190000 195.605000 65.390000 195.805000 ;
        RECT 65.190000 196.010000 65.390000 196.210000 ;
        RECT 65.190000 196.415000 65.390000 196.615000 ;
        RECT 65.190000 196.820000 65.390000 197.020000 ;
        RECT 65.190000 197.225000 65.390000 197.425000 ;
        RECT 65.190000 197.630000 65.390000 197.830000 ;
        RECT 65.190000 198.035000 65.390000 198.235000 ;
        RECT 65.190000 198.440000 65.390000 198.640000 ;
        RECT 65.190000 198.845000 65.390000 199.045000 ;
        RECT 65.190000 199.250000 65.390000 199.450000 ;
        RECT 65.190000 199.655000 65.390000 199.855000 ;
        RECT 65.495000  25.910000 65.695000  26.110000 ;
        RECT 65.495000  26.340000 65.695000  26.540000 ;
        RECT 65.495000  26.770000 65.695000  26.970000 ;
        RECT 65.495000  27.200000 65.695000  27.400000 ;
        RECT 65.495000  27.630000 65.695000  27.830000 ;
        RECT 65.495000  28.060000 65.695000  28.260000 ;
        RECT 65.495000  28.490000 65.695000  28.690000 ;
        RECT 65.495000  28.920000 65.695000  29.120000 ;
        RECT 65.495000  29.350000 65.695000  29.550000 ;
        RECT 65.495000  29.780000 65.695000  29.980000 ;
        RECT 65.495000  30.210000 65.695000  30.410000 ;
        RECT 65.590000 175.995000 65.790000 176.195000 ;
        RECT 65.590000 176.395000 65.790000 176.595000 ;
        RECT 65.590000 176.795000 65.790000 176.995000 ;
        RECT 65.590000 177.195000 65.790000 177.395000 ;
        RECT 65.590000 177.595000 65.790000 177.795000 ;
        RECT 65.590000 177.995000 65.790000 178.195000 ;
        RECT 65.590000 178.395000 65.790000 178.595000 ;
        RECT 65.590000 178.795000 65.790000 178.995000 ;
        RECT 65.590000 179.195000 65.790000 179.395000 ;
        RECT 65.590000 179.595000 65.790000 179.795000 ;
        RECT 65.590000 179.995000 65.790000 180.195000 ;
        RECT 65.590000 180.395000 65.790000 180.595000 ;
        RECT 65.590000 180.795000 65.790000 180.995000 ;
        RECT 65.590000 181.195000 65.790000 181.395000 ;
        RECT 65.590000 181.595000 65.790000 181.795000 ;
        RECT 65.590000 181.995000 65.790000 182.195000 ;
        RECT 65.590000 182.395000 65.790000 182.595000 ;
        RECT 65.590000 182.795000 65.790000 182.995000 ;
        RECT 65.590000 183.195000 65.790000 183.395000 ;
        RECT 65.590000 183.595000 65.790000 183.795000 ;
        RECT 65.590000 183.995000 65.790000 184.195000 ;
        RECT 65.590000 184.395000 65.790000 184.595000 ;
        RECT 65.590000 184.795000 65.790000 184.995000 ;
        RECT 65.590000 185.195000 65.790000 185.395000 ;
        RECT 65.590000 185.595000 65.790000 185.795000 ;
        RECT 65.590000 185.995000 65.790000 186.195000 ;
        RECT 65.590000 186.395000 65.790000 186.595000 ;
        RECT 65.590000 186.795000 65.790000 186.995000 ;
        RECT 65.590000 187.195000 65.790000 187.395000 ;
        RECT 65.590000 187.595000 65.790000 187.795000 ;
        RECT 65.590000 187.995000 65.790000 188.195000 ;
        RECT 65.590000 188.395000 65.790000 188.595000 ;
        RECT 65.590000 188.795000 65.790000 188.995000 ;
        RECT 65.590000 189.195000 65.790000 189.395000 ;
        RECT 65.590000 189.595000 65.790000 189.795000 ;
        RECT 65.590000 189.995000 65.790000 190.195000 ;
        RECT 65.590000 190.395000 65.790000 190.595000 ;
        RECT 65.590000 190.795000 65.790000 190.995000 ;
        RECT 65.590000 191.195000 65.790000 191.395000 ;
        RECT 65.590000 191.595000 65.790000 191.795000 ;
        RECT 65.590000 191.995000 65.790000 192.195000 ;
        RECT 65.590000 192.395000 65.790000 192.595000 ;
        RECT 65.590000 192.795000 65.790000 192.995000 ;
        RECT 65.590000 193.195000 65.790000 193.395000 ;
        RECT 65.590000 193.595000 65.790000 193.795000 ;
        RECT 65.590000 193.995000 65.790000 194.195000 ;
        RECT 65.590000 194.395000 65.790000 194.595000 ;
        RECT 65.590000 194.795000 65.790000 194.995000 ;
        RECT 65.590000 195.200000 65.790000 195.400000 ;
        RECT 65.590000 195.605000 65.790000 195.805000 ;
        RECT 65.590000 196.010000 65.790000 196.210000 ;
        RECT 65.590000 196.415000 65.790000 196.615000 ;
        RECT 65.590000 196.820000 65.790000 197.020000 ;
        RECT 65.590000 197.225000 65.790000 197.425000 ;
        RECT 65.590000 197.630000 65.790000 197.830000 ;
        RECT 65.590000 198.035000 65.790000 198.235000 ;
        RECT 65.590000 198.440000 65.790000 198.640000 ;
        RECT 65.590000 198.845000 65.790000 199.045000 ;
        RECT 65.590000 199.250000 65.790000 199.450000 ;
        RECT 65.590000 199.655000 65.790000 199.855000 ;
        RECT 65.900000  25.910000 66.100000  26.110000 ;
        RECT 65.900000  26.340000 66.100000  26.540000 ;
        RECT 65.900000  26.770000 66.100000  26.970000 ;
        RECT 65.900000  27.200000 66.100000  27.400000 ;
        RECT 65.900000  27.630000 66.100000  27.830000 ;
        RECT 65.900000  28.060000 66.100000  28.260000 ;
        RECT 65.900000  28.490000 66.100000  28.690000 ;
        RECT 65.900000  28.920000 66.100000  29.120000 ;
        RECT 65.900000  29.350000 66.100000  29.550000 ;
        RECT 65.900000  29.780000 66.100000  29.980000 ;
        RECT 65.900000  30.210000 66.100000  30.410000 ;
        RECT 65.990000 175.995000 66.190000 176.195000 ;
        RECT 65.990000 176.395000 66.190000 176.595000 ;
        RECT 65.990000 176.795000 66.190000 176.995000 ;
        RECT 65.990000 177.195000 66.190000 177.395000 ;
        RECT 65.990000 177.595000 66.190000 177.795000 ;
        RECT 65.990000 177.995000 66.190000 178.195000 ;
        RECT 65.990000 178.395000 66.190000 178.595000 ;
        RECT 65.990000 178.795000 66.190000 178.995000 ;
        RECT 65.990000 179.195000 66.190000 179.395000 ;
        RECT 65.990000 179.595000 66.190000 179.795000 ;
        RECT 65.990000 179.995000 66.190000 180.195000 ;
        RECT 65.990000 180.395000 66.190000 180.595000 ;
        RECT 65.990000 180.795000 66.190000 180.995000 ;
        RECT 65.990000 181.195000 66.190000 181.395000 ;
        RECT 65.990000 181.595000 66.190000 181.795000 ;
        RECT 65.990000 181.995000 66.190000 182.195000 ;
        RECT 65.990000 182.395000 66.190000 182.595000 ;
        RECT 65.990000 182.795000 66.190000 182.995000 ;
        RECT 65.990000 183.195000 66.190000 183.395000 ;
        RECT 65.990000 183.595000 66.190000 183.795000 ;
        RECT 65.990000 183.995000 66.190000 184.195000 ;
        RECT 65.990000 184.395000 66.190000 184.595000 ;
        RECT 65.990000 184.795000 66.190000 184.995000 ;
        RECT 65.990000 185.195000 66.190000 185.395000 ;
        RECT 65.990000 185.595000 66.190000 185.795000 ;
        RECT 65.990000 185.995000 66.190000 186.195000 ;
        RECT 65.990000 186.395000 66.190000 186.595000 ;
        RECT 65.990000 186.795000 66.190000 186.995000 ;
        RECT 65.990000 187.195000 66.190000 187.395000 ;
        RECT 65.990000 187.595000 66.190000 187.795000 ;
        RECT 65.990000 187.995000 66.190000 188.195000 ;
        RECT 65.990000 188.395000 66.190000 188.595000 ;
        RECT 65.990000 188.795000 66.190000 188.995000 ;
        RECT 65.990000 189.195000 66.190000 189.395000 ;
        RECT 65.990000 189.595000 66.190000 189.795000 ;
        RECT 65.990000 189.995000 66.190000 190.195000 ;
        RECT 65.990000 190.395000 66.190000 190.595000 ;
        RECT 65.990000 190.795000 66.190000 190.995000 ;
        RECT 65.990000 191.195000 66.190000 191.395000 ;
        RECT 65.990000 191.595000 66.190000 191.795000 ;
        RECT 65.990000 191.995000 66.190000 192.195000 ;
        RECT 65.990000 192.395000 66.190000 192.595000 ;
        RECT 65.990000 192.795000 66.190000 192.995000 ;
        RECT 65.990000 193.195000 66.190000 193.395000 ;
        RECT 65.990000 193.595000 66.190000 193.795000 ;
        RECT 65.990000 193.995000 66.190000 194.195000 ;
        RECT 65.990000 194.395000 66.190000 194.595000 ;
        RECT 65.990000 194.795000 66.190000 194.995000 ;
        RECT 65.990000 195.200000 66.190000 195.400000 ;
        RECT 65.990000 195.605000 66.190000 195.805000 ;
        RECT 65.990000 196.010000 66.190000 196.210000 ;
        RECT 65.990000 196.415000 66.190000 196.615000 ;
        RECT 65.990000 196.820000 66.190000 197.020000 ;
        RECT 65.990000 197.225000 66.190000 197.425000 ;
        RECT 65.990000 197.630000 66.190000 197.830000 ;
        RECT 65.990000 198.035000 66.190000 198.235000 ;
        RECT 65.990000 198.440000 66.190000 198.640000 ;
        RECT 65.990000 198.845000 66.190000 199.045000 ;
        RECT 65.990000 199.250000 66.190000 199.450000 ;
        RECT 65.990000 199.655000 66.190000 199.855000 ;
        RECT 66.305000  25.910000 66.505000  26.110000 ;
        RECT 66.305000  26.340000 66.505000  26.540000 ;
        RECT 66.305000  26.770000 66.505000  26.970000 ;
        RECT 66.305000  27.200000 66.505000  27.400000 ;
        RECT 66.305000  27.630000 66.505000  27.830000 ;
        RECT 66.305000  28.060000 66.505000  28.260000 ;
        RECT 66.305000  28.490000 66.505000  28.690000 ;
        RECT 66.305000  28.920000 66.505000  29.120000 ;
        RECT 66.305000  29.350000 66.505000  29.550000 ;
        RECT 66.305000  29.780000 66.505000  29.980000 ;
        RECT 66.305000  30.210000 66.505000  30.410000 ;
        RECT 66.390000 175.995000 66.590000 176.195000 ;
        RECT 66.390000 176.395000 66.590000 176.595000 ;
        RECT 66.390000 176.795000 66.590000 176.995000 ;
        RECT 66.390000 177.195000 66.590000 177.395000 ;
        RECT 66.390000 177.595000 66.590000 177.795000 ;
        RECT 66.390000 177.995000 66.590000 178.195000 ;
        RECT 66.390000 178.395000 66.590000 178.595000 ;
        RECT 66.390000 178.795000 66.590000 178.995000 ;
        RECT 66.390000 179.195000 66.590000 179.395000 ;
        RECT 66.390000 179.595000 66.590000 179.795000 ;
        RECT 66.390000 179.995000 66.590000 180.195000 ;
        RECT 66.390000 180.395000 66.590000 180.595000 ;
        RECT 66.390000 180.795000 66.590000 180.995000 ;
        RECT 66.390000 181.195000 66.590000 181.395000 ;
        RECT 66.390000 181.595000 66.590000 181.795000 ;
        RECT 66.390000 181.995000 66.590000 182.195000 ;
        RECT 66.390000 182.395000 66.590000 182.595000 ;
        RECT 66.390000 182.795000 66.590000 182.995000 ;
        RECT 66.390000 183.195000 66.590000 183.395000 ;
        RECT 66.390000 183.595000 66.590000 183.795000 ;
        RECT 66.390000 183.995000 66.590000 184.195000 ;
        RECT 66.390000 184.395000 66.590000 184.595000 ;
        RECT 66.390000 184.795000 66.590000 184.995000 ;
        RECT 66.390000 185.195000 66.590000 185.395000 ;
        RECT 66.390000 185.595000 66.590000 185.795000 ;
        RECT 66.390000 185.995000 66.590000 186.195000 ;
        RECT 66.390000 186.395000 66.590000 186.595000 ;
        RECT 66.390000 186.795000 66.590000 186.995000 ;
        RECT 66.390000 187.195000 66.590000 187.395000 ;
        RECT 66.390000 187.595000 66.590000 187.795000 ;
        RECT 66.390000 187.995000 66.590000 188.195000 ;
        RECT 66.390000 188.395000 66.590000 188.595000 ;
        RECT 66.390000 188.795000 66.590000 188.995000 ;
        RECT 66.390000 189.195000 66.590000 189.395000 ;
        RECT 66.390000 189.595000 66.590000 189.795000 ;
        RECT 66.390000 189.995000 66.590000 190.195000 ;
        RECT 66.390000 190.395000 66.590000 190.595000 ;
        RECT 66.390000 190.795000 66.590000 190.995000 ;
        RECT 66.390000 191.195000 66.590000 191.395000 ;
        RECT 66.390000 191.595000 66.590000 191.795000 ;
        RECT 66.390000 191.995000 66.590000 192.195000 ;
        RECT 66.390000 192.395000 66.590000 192.595000 ;
        RECT 66.390000 192.795000 66.590000 192.995000 ;
        RECT 66.390000 193.195000 66.590000 193.395000 ;
        RECT 66.390000 193.595000 66.590000 193.795000 ;
        RECT 66.390000 193.995000 66.590000 194.195000 ;
        RECT 66.390000 194.395000 66.590000 194.595000 ;
        RECT 66.390000 194.795000 66.590000 194.995000 ;
        RECT 66.390000 195.200000 66.590000 195.400000 ;
        RECT 66.390000 195.605000 66.590000 195.805000 ;
        RECT 66.390000 196.010000 66.590000 196.210000 ;
        RECT 66.390000 196.415000 66.590000 196.615000 ;
        RECT 66.390000 196.820000 66.590000 197.020000 ;
        RECT 66.390000 197.225000 66.590000 197.425000 ;
        RECT 66.390000 197.630000 66.590000 197.830000 ;
        RECT 66.390000 198.035000 66.590000 198.235000 ;
        RECT 66.390000 198.440000 66.590000 198.640000 ;
        RECT 66.390000 198.845000 66.590000 199.045000 ;
        RECT 66.390000 199.250000 66.590000 199.450000 ;
        RECT 66.390000 199.655000 66.590000 199.855000 ;
        RECT 66.710000  25.910000 66.910000  26.110000 ;
        RECT 66.710000  26.340000 66.910000  26.540000 ;
        RECT 66.710000  26.770000 66.910000  26.970000 ;
        RECT 66.710000  27.200000 66.910000  27.400000 ;
        RECT 66.710000  27.630000 66.910000  27.830000 ;
        RECT 66.710000  28.060000 66.910000  28.260000 ;
        RECT 66.710000  28.490000 66.910000  28.690000 ;
        RECT 66.710000  28.920000 66.910000  29.120000 ;
        RECT 66.710000  29.350000 66.910000  29.550000 ;
        RECT 66.710000  29.780000 66.910000  29.980000 ;
        RECT 66.710000  30.210000 66.910000  30.410000 ;
        RECT 66.790000 175.995000 66.990000 176.195000 ;
        RECT 66.790000 176.395000 66.990000 176.595000 ;
        RECT 66.790000 176.795000 66.990000 176.995000 ;
        RECT 66.790000 177.195000 66.990000 177.395000 ;
        RECT 66.790000 177.595000 66.990000 177.795000 ;
        RECT 66.790000 177.995000 66.990000 178.195000 ;
        RECT 66.790000 178.395000 66.990000 178.595000 ;
        RECT 66.790000 178.795000 66.990000 178.995000 ;
        RECT 66.790000 179.195000 66.990000 179.395000 ;
        RECT 66.790000 179.595000 66.990000 179.795000 ;
        RECT 66.790000 179.995000 66.990000 180.195000 ;
        RECT 66.790000 180.395000 66.990000 180.595000 ;
        RECT 66.790000 180.795000 66.990000 180.995000 ;
        RECT 66.790000 181.195000 66.990000 181.395000 ;
        RECT 66.790000 181.595000 66.990000 181.795000 ;
        RECT 66.790000 181.995000 66.990000 182.195000 ;
        RECT 66.790000 182.395000 66.990000 182.595000 ;
        RECT 66.790000 182.795000 66.990000 182.995000 ;
        RECT 66.790000 183.195000 66.990000 183.395000 ;
        RECT 66.790000 183.595000 66.990000 183.795000 ;
        RECT 66.790000 183.995000 66.990000 184.195000 ;
        RECT 66.790000 184.395000 66.990000 184.595000 ;
        RECT 66.790000 184.795000 66.990000 184.995000 ;
        RECT 66.790000 185.195000 66.990000 185.395000 ;
        RECT 66.790000 185.595000 66.990000 185.795000 ;
        RECT 66.790000 185.995000 66.990000 186.195000 ;
        RECT 66.790000 186.395000 66.990000 186.595000 ;
        RECT 66.790000 186.795000 66.990000 186.995000 ;
        RECT 66.790000 187.195000 66.990000 187.395000 ;
        RECT 66.790000 187.595000 66.990000 187.795000 ;
        RECT 66.790000 187.995000 66.990000 188.195000 ;
        RECT 66.790000 188.395000 66.990000 188.595000 ;
        RECT 66.790000 188.795000 66.990000 188.995000 ;
        RECT 66.790000 189.195000 66.990000 189.395000 ;
        RECT 66.790000 189.595000 66.990000 189.795000 ;
        RECT 66.790000 189.995000 66.990000 190.195000 ;
        RECT 66.790000 190.395000 66.990000 190.595000 ;
        RECT 66.790000 190.795000 66.990000 190.995000 ;
        RECT 66.790000 191.195000 66.990000 191.395000 ;
        RECT 66.790000 191.595000 66.990000 191.795000 ;
        RECT 66.790000 191.995000 66.990000 192.195000 ;
        RECT 66.790000 192.395000 66.990000 192.595000 ;
        RECT 66.790000 192.795000 66.990000 192.995000 ;
        RECT 66.790000 193.195000 66.990000 193.395000 ;
        RECT 66.790000 193.595000 66.990000 193.795000 ;
        RECT 66.790000 193.995000 66.990000 194.195000 ;
        RECT 66.790000 194.395000 66.990000 194.595000 ;
        RECT 66.790000 194.795000 66.990000 194.995000 ;
        RECT 66.790000 195.200000 66.990000 195.400000 ;
        RECT 66.790000 195.605000 66.990000 195.805000 ;
        RECT 66.790000 196.010000 66.990000 196.210000 ;
        RECT 66.790000 196.415000 66.990000 196.615000 ;
        RECT 66.790000 196.820000 66.990000 197.020000 ;
        RECT 66.790000 197.225000 66.990000 197.425000 ;
        RECT 66.790000 197.630000 66.990000 197.830000 ;
        RECT 66.790000 198.035000 66.990000 198.235000 ;
        RECT 66.790000 198.440000 66.990000 198.640000 ;
        RECT 66.790000 198.845000 66.990000 199.045000 ;
        RECT 66.790000 199.250000 66.990000 199.450000 ;
        RECT 66.790000 199.655000 66.990000 199.855000 ;
        RECT 67.115000  25.910000 67.315000  26.110000 ;
        RECT 67.115000  26.340000 67.315000  26.540000 ;
        RECT 67.115000  26.770000 67.315000  26.970000 ;
        RECT 67.115000  27.200000 67.315000  27.400000 ;
        RECT 67.115000  27.630000 67.315000  27.830000 ;
        RECT 67.115000  28.060000 67.315000  28.260000 ;
        RECT 67.115000  28.490000 67.315000  28.690000 ;
        RECT 67.115000  28.920000 67.315000  29.120000 ;
        RECT 67.115000  29.350000 67.315000  29.550000 ;
        RECT 67.115000  29.780000 67.315000  29.980000 ;
        RECT 67.115000  30.210000 67.315000  30.410000 ;
        RECT 67.190000 175.995000 67.390000 176.195000 ;
        RECT 67.190000 176.395000 67.390000 176.595000 ;
        RECT 67.190000 176.795000 67.390000 176.995000 ;
        RECT 67.190000 177.195000 67.390000 177.395000 ;
        RECT 67.190000 177.595000 67.390000 177.795000 ;
        RECT 67.190000 177.995000 67.390000 178.195000 ;
        RECT 67.190000 178.395000 67.390000 178.595000 ;
        RECT 67.190000 178.795000 67.390000 178.995000 ;
        RECT 67.190000 179.195000 67.390000 179.395000 ;
        RECT 67.190000 179.595000 67.390000 179.795000 ;
        RECT 67.190000 179.995000 67.390000 180.195000 ;
        RECT 67.190000 180.395000 67.390000 180.595000 ;
        RECT 67.190000 180.795000 67.390000 180.995000 ;
        RECT 67.190000 181.195000 67.390000 181.395000 ;
        RECT 67.190000 181.595000 67.390000 181.795000 ;
        RECT 67.190000 181.995000 67.390000 182.195000 ;
        RECT 67.190000 182.395000 67.390000 182.595000 ;
        RECT 67.190000 182.795000 67.390000 182.995000 ;
        RECT 67.190000 183.195000 67.390000 183.395000 ;
        RECT 67.190000 183.595000 67.390000 183.795000 ;
        RECT 67.190000 183.995000 67.390000 184.195000 ;
        RECT 67.190000 184.395000 67.390000 184.595000 ;
        RECT 67.190000 184.795000 67.390000 184.995000 ;
        RECT 67.190000 185.195000 67.390000 185.395000 ;
        RECT 67.190000 185.595000 67.390000 185.795000 ;
        RECT 67.190000 185.995000 67.390000 186.195000 ;
        RECT 67.190000 186.395000 67.390000 186.595000 ;
        RECT 67.190000 186.795000 67.390000 186.995000 ;
        RECT 67.190000 187.195000 67.390000 187.395000 ;
        RECT 67.190000 187.595000 67.390000 187.795000 ;
        RECT 67.190000 187.995000 67.390000 188.195000 ;
        RECT 67.190000 188.395000 67.390000 188.595000 ;
        RECT 67.190000 188.795000 67.390000 188.995000 ;
        RECT 67.190000 189.195000 67.390000 189.395000 ;
        RECT 67.190000 189.595000 67.390000 189.795000 ;
        RECT 67.190000 189.995000 67.390000 190.195000 ;
        RECT 67.190000 190.395000 67.390000 190.595000 ;
        RECT 67.190000 190.795000 67.390000 190.995000 ;
        RECT 67.190000 191.195000 67.390000 191.395000 ;
        RECT 67.190000 191.595000 67.390000 191.795000 ;
        RECT 67.190000 191.995000 67.390000 192.195000 ;
        RECT 67.190000 192.395000 67.390000 192.595000 ;
        RECT 67.190000 192.795000 67.390000 192.995000 ;
        RECT 67.190000 193.195000 67.390000 193.395000 ;
        RECT 67.190000 193.595000 67.390000 193.795000 ;
        RECT 67.190000 193.995000 67.390000 194.195000 ;
        RECT 67.190000 194.395000 67.390000 194.595000 ;
        RECT 67.190000 194.795000 67.390000 194.995000 ;
        RECT 67.190000 195.200000 67.390000 195.400000 ;
        RECT 67.190000 195.605000 67.390000 195.805000 ;
        RECT 67.190000 196.010000 67.390000 196.210000 ;
        RECT 67.190000 196.415000 67.390000 196.615000 ;
        RECT 67.190000 196.820000 67.390000 197.020000 ;
        RECT 67.190000 197.225000 67.390000 197.425000 ;
        RECT 67.190000 197.630000 67.390000 197.830000 ;
        RECT 67.190000 198.035000 67.390000 198.235000 ;
        RECT 67.190000 198.440000 67.390000 198.640000 ;
        RECT 67.190000 198.845000 67.390000 199.045000 ;
        RECT 67.190000 199.250000 67.390000 199.450000 ;
        RECT 67.190000 199.655000 67.390000 199.855000 ;
        RECT 67.520000  25.910000 67.720000  26.110000 ;
        RECT 67.520000  26.340000 67.720000  26.540000 ;
        RECT 67.520000  26.770000 67.720000  26.970000 ;
        RECT 67.520000  27.200000 67.720000  27.400000 ;
        RECT 67.520000  27.630000 67.720000  27.830000 ;
        RECT 67.520000  28.060000 67.720000  28.260000 ;
        RECT 67.520000  28.490000 67.720000  28.690000 ;
        RECT 67.520000  28.920000 67.720000  29.120000 ;
        RECT 67.520000  29.350000 67.720000  29.550000 ;
        RECT 67.520000  29.780000 67.720000  29.980000 ;
        RECT 67.520000  30.210000 67.720000  30.410000 ;
        RECT 67.590000 175.995000 67.790000 176.195000 ;
        RECT 67.590000 176.395000 67.790000 176.595000 ;
        RECT 67.590000 176.795000 67.790000 176.995000 ;
        RECT 67.590000 177.195000 67.790000 177.395000 ;
        RECT 67.590000 177.595000 67.790000 177.795000 ;
        RECT 67.590000 177.995000 67.790000 178.195000 ;
        RECT 67.590000 178.395000 67.790000 178.595000 ;
        RECT 67.590000 178.795000 67.790000 178.995000 ;
        RECT 67.590000 179.195000 67.790000 179.395000 ;
        RECT 67.590000 179.595000 67.790000 179.795000 ;
        RECT 67.590000 179.995000 67.790000 180.195000 ;
        RECT 67.590000 180.395000 67.790000 180.595000 ;
        RECT 67.590000 180.795000 67.790000 180.995000 ;
        RECT 67.590000 181.195000 67.790000 181.395000 ;
        RECT 67.590000 181.595000 67.790000 181.795000 ;
        RECT 67.590000 181.995000 67.790000 182.195000 ;
        RECT 67.590000 182.395000 67.790000 182.595000 ;
        RECT 67.590000 182.795000 67.790000 182.995000 ;
        RECT 67.590000 183.195000 67.790000 183.395000 ;
        RECT 67.590000 183.595000 67.790000 183.795000 ;
        RECT 67.590000 183.995000 67.790000 184.195000 ;
        RECT 67.590000 184.395000 67.790000 184.595000 ;
        RECT 67.590000 184.795000 67.790000 184.995000 ;
        RECT 67.590000 185.195000 67.790000 185.395000 ;
        RECT 67.590000 185.595000 67.790000 185.795000 ;
        RECT 67.590000 185.995000 67.790000 186.195000 ;
        RECT 67.590000 186.395000 67.790000 186.595000 ;
        RECT 67.590000 186.795000 67.790000 186.995000 ;
        RECT 67.590000 187.195000 67.790000 187.395000 ;
        RECT 67.590000 187.595000 67.790000 187.795000 ;
        RECT 67.590000 187.995000 67.790000 188.195000 ;
        RECT 67.590000 188.395000 67.790000 188.595000 ;
        RECT 67.590000 188.795000 67.790000 188.995000 ;
        RECT 67.590000 189.195000 67.790000 189.395000 ;
        RECT 67.590000 189.595000 67.790000 189.795000 ;
        RECT 67.590000 189.995000 67.790000 190.195000 ;
        RECT 67.590000 190.395000 67.790000 190.595000 ;
        RECT 67.590000 190.795000 67.790000 190.995000 ;
        RECT 67.590000 191.195000 67.790000 191.395000 ;
        RECT 67.590000 191.595000 67.790000 191.795000 ;
        RECT 67.590000 191.995000 67.790000 192.195000 ;
        RECT 67.590000 192.395000 67.790000 192.595000 ;
        RECT 67.590000 192.795000 67.790000 192.995000 ;
        RECT 67.590000 193.195000 67.790000 193.395000 ;
        RECT 67.590000 193.595000 67.790000 193.795000 ;
        RECT 67.590000 193.995000 67.790000 194.195000 ;
        RECT 67.590000 194.395000 67.790000 194.595000 ;
        RECT 67.590000 194.795000 67.790000 194.995000 ;
        RECT 67.590000 195.200000 67.790000 195.400000 ;
        RECT 67.590000 195.605000 67.790000 195.805000 ;
        RECT 67.590000 196.010000 67.790000 196.210000 ;
        RECT 67.590000 196.415000 67.790000 196.615000 ;
        RECT 67.590000 196.820000 67.790000 197.020000 ;
        RECT 67.590000 197.225000 67.790000 197.425000 ;
        RECT 67.590000 197.630000 67.790000 197.830000 ;
        RECT 67.590000 198.035000 67.790000 198.235000 ;
        RECT 67.590000 198.440000 67.790000 198.640000 ;
        RECT 67.590000 198.845000 67.790000 199.045000 ;
        RECT 67.590000 199.250000 67.790000 199.450000 ;
        RECT 67.590000 199.655000 67.790000 199.855000 ;
        RECT 67.925000  25.910000 68.125000  26.110000 ;
        RECT 67.925000  26.340000 68.125000  26.540000 ;
        RECT 67.925000  26.770000 68.125000  26.970000 ;
        RECT 67.925000  27.200000 68.125000  27.400000 ;
        RECT 67.925000  27.630000 68.125000  27.830000 ;
        RECT 67.925000  28.060000 68.125000  28.260000 ;
        RECT 67.925000  28.490000 68.125000  28.690000 ;
        RECT 67.925000  28.920000 68.125000  29.120000 ;
        RECT 67.925000  29.350000 68.125000  29.550000 ;
        RECT 67.925000  29.780000 68.125000  29.980000 ;
        RECT 67.925000  30.210000 68.125000  30.410000 ;
        RECT 67.990000 175.995000 68.190000 176.195000 ;
        RECT 67.990000 176.395000 68.190000 176.595000 ;
        RECT 67.990000 176.795000 68.190000 176.995000 ;
        RECT 67.990000 177.195000 68.190000 177.395000 ;
        RECT 67.990000 177.595000 68.190000 177.795000 ;
        RECT 67.990000 177.995000 68.190000 178.195000 ;
        RECT 67.990000 178.395000 68.190000 178.595000 ;
        RECT 67.990000 178.795000 68.190000 178.995000 ;
        RECT 67.990000 179.195000 68.190000 179.395000 ;
        RECT 67.990000 179.595000 68.190000 179.795000 ;
        RECT 67.990000 179.995000 68.190000 180.195000 ;
        RECT 67.990000 180.395000 68.190000 180.595000 ;
        RECT 67.990000 180.795000 68.190000 180.995000 ;
        RECT 67.990000 181.195000 68.190000 181.395000 ;
        RECT 67.990000 181.595000 68.190000 181.795000 ;
        RECT 67.990000 181.995000 68.190000 182.195000 ;
        RECT 67.990000 182.395000 68.190000 182.595000 ;
        RECT 67.990000 182.795000 68.190000 182.995000 ;
        RECT 67.990000 183.195000 68.190000 183.395000 ;
        RECT 67.990000 183.595000 68.190000 183.795000 ;
        RECT 67.990000 183.995000 68.190000 184.195000 ;
        RECT 67.990000 184.395000 68.190000 184.595000 ;
        RECT 67.990000 184.795000 68.190000 184.995000 ;
        RECT 67.990000 185.195000 68.190000 185.395000 ;
        RECT 67.990000 185.595000 68.190000 185.795000 ;
        RECT 67.990000 185.995000 68.190000 186.195000 ;
        RECT 67.990000 186.395000 68.190000 186.595000 ;
        RECT 67.990000 186.795000 68.190000 186.995000 ;
        RECT 67.990000 187.195000 68.190000 187.395000 ;
        RECT 67.990000 187.595000 68.190000 187.795000 ;
        RECT 67.990000 187.995000 68.190000 188.195000 ;
        RECT 67.990000 188.395000 68.190000 188.595000 ;
        RECT 67.990000 188.795000 68.190000 188.995000 ;
        RECT 67.990000 189.195000 68.190000 189.395000 ;
        RECT 67.990000 189.595000 68.190000 189.795000 ;
        RECT 67.990000 189.995000 68.190000 190.195000 ;
        RECT 67.990000 190.395000 68.190000 190.595000 ;
        RECT 67.990000 190.795000 68.190000 190.995000 ;
        RECT 67.990000 191.195000 68.190000 191.395000 ;
        RECT 67.990000 191.595000 68.190000 191.795000 ;
        RECT 67.990000 191.995000 68.190000 192.195000 ;
        RECT 67.990000 192.395000 68.190000 192.595000 ;
        RECT 67.990000 192.795000 68.190000 192.995000 ;
        RECT 67.990000 193.195000 68.190000 193.395000 ;
        RECT 67.990000 193.595000 68.190000 193.795000 ;
        RECT 67.990000 193.995000 68.190000 194.195000 ;
        RECT 67.990000 194.395000 68.190000 194.595000 ;
        RECT 67.990000 194.795000 68.190000 194.995000 ;
        RECT 67.990000 195.200000 68.190000 195.400000 ;
        RECT 67.990000 195.605000 68.190000 195.805000 ;
        RECT 67.990000 196.010000 68.190000 196.210000 ;
        RECT 67.990000 196.415000 68.190000 196.615000 ;
        RECT 67.990000 196.820000 68.190000 197.020000 ;
        RECT 67.990000 197.225000 68.190000 197.425000 ;
        RECT 67.990000 197.630000 68.190000 197.830000 ;
        RECT 67.990000 198.035000 68.190000 198.235000 ;
        RECT 67.990000 198.440000 68.190000 198.640000 ;
        RECT 67.990000 198.845000 68.190000 199.045000 ;
        RECT 67.990000 199.250000 68.190000 199.450000 ;
        RECT 67.990000 199.655000 68.190000 199.855000 ;
        RECT 68.330000  25.910000 68.530000  26.110000 ;
        RECT 68.330000  26.340000 68.530000  26.540000 ;
        RECT 68.330000  26.770000 68.530000  26.970000 ;
        RECT 68.330000  27.200000 68.530000  27.400000 ;
        RECT 68.330000  27.630000 68.530000  27.830000 ;
        RECT 68.330000  28.060000 68.530000  28.260000 ;
        RECT 68.330000  28.490000 68.530000  28.690000 ;
        RECT 68.330000  28.920000 68.530000  29.120000 ;
        RECT 68.330000  29.350000 68.530000  29.550000 ;
        RECT 68.330000  29.780000 68.530000  29.980000 ;
        RECT 68.330000  30.210000 68.530000  30.410000 ;
        RECT 68.390000 175.995000 68.590000 176.195000 ;
        RECT 68.390000 176.395000 68.590000 176.595000 ;
        RECT 68.390000 176.795000 68.590000 176.995000 ;
        RECT 68.390000 177.195000 68.590000 177.395000 ;
        RECT 68.390000 177.595000 68.590000 177.795000 ;
        RECT 68.390000 177.995000 68.590000 178.195000 ;
        RECT 68.390000 178.395000 68.590000 178.595000 ;
        RECT 68.390000 178.795000 68.590000 178.995000 ;
        RECT 68.390000 179.195000 68.590000 179.395000 ;
        RECT 68.390000 179.595000 68.590000 179.795000 ;
        RECT 68.390000 179.995000 68.590000 180.195000 ;
        RECT 68.390000 180.395000 68.590000 180.595000 ;
        RECT 68.390000 180.795000 68.590000 180.995000 ;
        RECT 68.390000 181.195000 68.590000 181.395000 ;
        RECT 68.390000 181.595000 68.590000 181.795000 ;
        RECT 68.390000 181.995000 68.590000 182.195000 ;
        RECT 68.390000 182.395000 68.590000 182.595000 ;
        RECT 68.390000 182.795000 68.590000 182.995000 ;
        RECT 68.390000 183.195000 68.590000 183.395000 ;
        RECT 68.390000 183.595000 68.590000 183.795000 ;
        RECT 68.390000 183.995000 68.590000 184.195000 ;
        RECT 68.390000 184.395000 68.590000 184.595000 ;
        RECT 68.390000 184.795000 68.590000 184.995000 ;
        RECT 68.390000 185.195000 68.590000 185.395000 ;
        RECT 68.390000 185.595000 68.590000 185.795000 ;
        RECT 68.390000 185.995000 68.590000 186.195000 ;
        RECT 68.390000 186.395000 68.590000 186.595000 ;
        RECT 68.390000 186.795000 68.590000 186.995000 ;
        RECT 68.390000 187.195000 68.590000 187.395000 ;
        RECT 68.390000 187.595000 68.590000 187.795000 ;
        RECT 68.390000 187.995000 68.590000 188.195000 ;
        RECT 68.390000 188.395000 68.590000 188.595000 ;
        RECT 68.390000 188.795000 68.590000 188.995000 ;
        RECT 68.390000 189.195000 68.590000 189.395000 ;
        RECT 68.390000 189.595000 68.590000 189.795000 ;
        RECT 68.390000 189.995000 68.590000 190.195000 ;
        RECT 68.390000 190.395000 68.590000 190.595000 ;
        RECT 68.390000 190.795000 68.590000 190.995000 ;
        RECT 68.390000 191.195000 68.590000 191.395000 ;
        RECT 68.390000 191.595000 68.590000 191.795000 ;
        RECT 68.390000 191.995000 68.590000 192.195000 ;
        RECT 68.390000 192.395000 68.590000 192.595000 ;
        RECT 68.390000 192.795000 68.590000 192.995000 ;
        RECT 68.390000 193.195000 68.590000 193.395000 ;
        RECT 68.390000 193.595000 68.590000 193.795000 ;
        RECT 68.390000 193.995000 68.590000 194.195000 ;
        RECT 68.390000 194.395000 68.590000 194.595000 ;
        RECT 68.390000 194.795000 68.590000 194.995000 ;
        RECT 68.390000 195.200000 68.590000 195.400000 ;
        RECT 68.390000 195.605000 68.590000 195.805000 ;
        RECT 68.390000 196.010000 68.590000 196.210000 ;
        RECT 68.390000 196.415000 68.590000 196.615000 ;
        RECT 68.390000 196.820000 68.590000 197.020000 ;
        RECT 68.390000 197.225000 68.590000 197.425000 ;
        RECT 68.390000 197.630000 68.590000 197.830000 ;
        RECT 68.390000 198.035000 68.590000 198.235000 ;
        RECT 68.390000 198.440000 68.590000 198.640000 ;
        RECT 68.390000 198.845000 68.590000 199.045000 ;
        RECT 68.390000 199.250000 68.590000 199.450000 ;
        RECT 68.390000 199.655000 68.590000 199.855000 ;
        RECT 68.735000  25.910000 68.935000  26.110000 ;
        RECT 68.735000  26.340000 68.935000  26.540000 ;
        RECT 68.735000  26.770000 68.935000  26.970000 ;
        RECT 68.735000  27.200000 68.935000  27.400000 ;
        RECT 68.735000  27.630000 68.935000  27.830000 ;
        RECT 68.735000  28.060000 68.935000  28.260000 ;
        RECT 68.735000  28.490000 68.935000  28.690000 ;
        RECT 68.735000  28.920000 68.935000  29.120000 ;
        RECT 68.735000  29.350000 68.935000  29.550000 ;
        RECT 68.735000  29.780000 68.935000  29.980000 ;
        RECT 68.735000  30.210000 68.935000  30.410000 ;
        RECT 68.790000 175.995000 68.990000 176.195000 ;
        RECT 68.790000 176.395000 68.990000 176.595000 ;
        RECT 68.790000 176.795000 68.990000 176.995000 ;
        RECT 68.790000 177.195000 68.990000 177.395000 ;
        RECT 68.790000 177.595000 68.990000 177.795000 ;
        RECT 68.790000 177.995000 68.990000 178.195000 ;
        RECT 68.790000 178.395000 68.990000 178.595000 ;
        RECT 68.790000 178.795000 68.990000 178.995000 ;
        RECT 68.790000 179.195000 68.990000 179.395000 ;
        RECT 68.790000 179.595000 68.990000 179.795000 ;
        RECT 68.790000 179.995000 68.990000 180.195000 ;
        RECT 68.790000 180.395000 68.990000 180.595000 ;
        RECT 68.790000 180.795000 68.990000 180.995000 ;
        RECT 68.790000 181.195000 68.990000 181.395000 ;
        RECT 68.790000 181.595000 68.990000 181.795000 ;
        RECT 68.790000 181.995000 68.990000 182.195000 ;
        RECT 68.790000 182.395000 68.990000 182.595000 ;
        RECT 68.790000 182.795000 68.990000 182.995000 ;
        RECT 68.790000 183.195000 68.990000 183.395000 ;
        RECT 68.790000 183.595000 68.990000 183.795000 ;
        RECT 68.790000 183.995000 68.990000 184.195000 ;
        RECT 68.790000 184.395000 68.990000 184.595000 ;
        RECT 68.790000 184.795000 68.990000 184.995000 ;
        RECT 68.790000 185.195000 68.990000 185.395000 ;
        RECT 68.790000 185.595000 68.990000 185.795000 ;
        RECT 68.790000 185.995000 68.990000 186.195000 ;
        RECT 68.790000 186.395000 68.990000 186.595000 ;
        RECT 68.790000 186.795000 68.990000 186.995000 ;
        RECT 68.790000 187.195000 68.990000 187.395000 ;
        RECT 68.790000 187.595000 68.990000 187.795000 ;
        RECT 68.790000 187.995000 68.990000 188.195000 ;
        RECT 68.790000 188.395000 68.990000 188.595000 ;
        RECT 68.790000 188.795000 68.990000 188.995000 ;
        RECT 68.790000 189.195000 68.990000 189.395000 ;
        RECT 68.790000 189.595000 68.990000 189.795000 ;
        RECT 68.790000 189.995000 68.990000 190.195000 ;
        RECT 68.790000 190.395000 68.990000 190.595000 ;
        RECT 68.790000 190.795000 68.990000 190.995000 ;
        RECT 68.790000 191.195000 68.990000 191.395000 ;
        RECT 68.790000 191.595000 68.990000 191.795000 ;
        RECT 68.790000 191.995000 68.990000 192.195000 ;
        RECT 68.790000 192.395000 68.990000 192.595000 ;
        RECT 68.790000 192.795000 68.990000 192.995000 ;
        RECT 68.790000 193.195000 68.990000 193.395000 ;
        RECT 68.790000 193.595000 68.990000 193.795000 ;
        RECT 68.790000 193.995000 68.990000 194.195000 ;
        RECT 68.790000 194.395000 68.990000 194.595000 ;
        RECT 68.790000 194.795000 68.990000 194.995000 ;
        RECT 68.790000 195.200000 68.990000 195.400000 ;
        RECT 68.790000 195.605000 68.990000 195.805000 ;
        RECT 68.790000 196.010000 68.990000 196.210000 ;
        RECT 68.790000 196.415000 68.990000 196.615000 ;
        RECT 68.790000 196.820000 68.990000 197.020000 ;
        RECT 68.790000 197.225000 68.990000 197.425000 ;
        RECT 68.790000 197.630000 68.990000 197.830000 ;
        RECT 68.790000 198.035000 68.990000 198.235000 ;
        RECT 68.790000 198.440000 68.990000 198.640000 ;
        RECT 68.790000 198.845000 68.990000 199.045000 ;
        RECT 68.790000 199.250000 68.990000 199.450000 ;
        RECT 68.790000 199.655000 68.990000 199.855000 ;
        RECT 69.140000  25.910000 69.340000  26.110000 ;
        RECT 69.140000  26.340000 69.340000  26.540000 ;
        RECT 69.140000  26.770000 69.340000  26.970000 ;
        RECT 69.140000  27.200000 69.340000  27.400000 ;
        RECT 69.140000  27.630000 69.340000  27.830000 ;
        RECT 69.140000  28.060000 69.340000  28.260000 ;
        RECT 69.140000  28.490000 69.340000  28.690000 ;
        RECT 69.140000  28.920000 69.340000  29.120000 ;
        RECT 69.140000  29.350000 69.340000  29.550000 ;
        RECT 69.140000  29.780000 69.340000  29.980000 ;
        RECT 69.140000  30.210000 69.340000  30.410000 ;
        RECT 69.190000 175.995000 69.390000 176.195000 ;
        RECT 69.190000 176.395000 69.390000 176.595000 ;
        RECT 69.190000 176.795000 69.390000 176.995000 ;
        RECT 69.190000 177.195000 69.390000 177.395000 ;
        RECT 69.190000 177.595000 69.390000 177.795000 ;
        RECT 69.190000 177.995000 69.390000 178.195000 ;
        RECT 69.190000 178.395000 69.390000 178.595000 ;
        RECT 69.190000 178.795000 69.390000 178.995000 ;
        RECT 69.190000 179.195000 69.390000 179.395000 ;
        RECT 69.190000 179.595000 69.390000 179.795000 ;
        RECT 69.190000 179.995000 69.390000 180.195000 ;
        RECT 69.190000 180.395000 69.390000 180.595000 ;
        RECT 69.190000 180.795000 69.390000 180.995000 ;
        RECT 69.190000 181.195000 69.390000 181.395000 ;
        RECT 69.190000 181.595000 69.390000 181.795000 ;
        RECT 69.190000 181.995000 69.390000 182.195000 ;
        RECT 69.190000 182.395000 69.390000 182.595000 ;
        RECT 69.190000 182.795000 69.390000 182.995000 ;
        RECT 69.190000 183.195000 69.390000 183.395000 ;
        RECT 69.190000 183.595000 69.390000 183.795000 ;
        RECT 69.190000 183.995000 69.390000 184.195000 ;
        RECT 69.190000 184.395000 69.390000 184.595000 ;
        RECT 69.190000 184.795000 69.390000 184.995000 ;
        RECT 69.190000 185.195000 69.390000 185.395000 ;
        RECT 69.190000 185.595000 69.390000 185.795000 ;
        RECT 69.190000 185.995000 69.390000 186.195000 ;
        RECT 69.190000 186.395000 69.390000 186.595000 ;
        RECT 69.190000 186.795000 69.390000 186.995000 ;
        RECT 69.190000 187.195000 69.390000 187.395000 ;
        RECT 69.190000 187.595000 69.390000 187.795000 ;
        RECT 69.190000 187.995000 69.390000 188.195000 ;
        RECT 69.190000 188.395000 69.390000 188.595000 ;
        RECT 69.190000 188.795000 69.390000 188.995000 ;
        RECT 69.190000 189.195000 69.390000 189.395000 ;
        RECT 69.190000 189.595000 69.390000 189.795000 ;
        RECT 69.190000 189.995000 69.390000 190.195000 ;
        RECT 69.190000 190.395000 69.390000 190.595000 ;
        RECT 69.190000 190.795000 69.390000 190.995000 ;
        RECT 69.190000 191.195000 69.390000 191.395000 ;
        RECT 69.190000 191.595000 69.390000 191.795000 ;
        RECT 69.190000 191.995000 69.390000 192.195000 ;
        RECT 69.190000 192.395000 69.390000 192.595000 ;
        RECT 69.190000 192.795000 69.390000 192.995000 ;
        RECT 69.190000 193.195000 69.390000 193.395000 ;
        RECT 69.190000 193.595000 69.390000 193.795000 ;
        RECT 69.190000 193.995000 69.390000 194.195000 ;
        RECT 69.190000 194.395000 69.390000 194.595000 ;
        RECT 69.190000 194.795000 69.390000 194.995000 ;
        RECT 69.190000 195.200000 69.390000 195.400000 ;
        RECT 69.190000 195.605000 69.390000 195.805000 ;
        RECT 69.190000 196.010000 69.390000 196.210000 ;
        RECT 69.190000 196.415000 69.390000 196.615000 ;
        RECT 69.190000 196.820000 69.390000 197.020000 ;
        RECT 69.190000 197.225000 69.390000 197.425000 ;
        RECT 69.190000 197.630000 69.390000 197.830000 ;
        RECT 69.190000 198.035000 69.390000 198.235000 ;
        RECT 69.190000 198.440000 69.390000 198.640000 ;
        RECT 69.190000 198.845000 69.390000 199.045000 ;
        RECT 69.190000 199.250000 69.390000 199.450000 ;
        RECT 69.190000 199.655000 69.390000 199.855000 ;
        RECT 69.545000  25.910000 69.745000  26.110000 ;
        RECT 69.545000  26.340000 69.745000  26.540000 ;
        RECT 69.545000  26.770000 69.745000  26.970000 ;
        RECT 69.545000  27.200000 69.745000  27.400000 ;
        RECT 69.545000  27.630000 69.745000  27.830000 ;
        RECT 69.545000  28.060000 69.745000  28.260000 ;
        RECT 69.545000  28.490000 69.745000  28.690000 ;
        RECT 69.545000  28.920000 69.745000  29.120000 ;
        RECT 69.545000  29.350000 69.745000  29.550000 ;
        RECT 69.545000  29.780000 69.745000  29.980000 ;
        RECT 69.545000  30.210000 69.745000  30.410000 ;
        RECT 69.590000 175.995000 69.790000 176.195000 ;
        RECT 69.590000 176.395000 69.790000 176.595000 ;
        RECT 69.590000 176.795000 69.790000 176.995000 ;
        RECT 69.590000 177.195000 69.790000 177.395000 ;
        RECT 69.590000 177.595000 69.790000 177.795000 ;
        RECT 69.590000 177.995000 69.790000 178.195000 ;
        RECT 69.590000 178.395000 69.790000 178.595000 ;
        RECT 69.590000 178.795000 69.790000 178.995000 ;
        RECT 69.590000 179.195000 69.790000 179.395000 ;
        RECT 69.590000 179.595000 69.790000 179.795000 ;
        RECT 69.590000 179.995000 69.790000 180.195000 ;
        RECT 69.590000 180.395000 69.790000 180.595000 ;
        RECT 69.590000 180.795000 69.790000 180.995000 ;
        RECT 69.590000 181.195000 69.790000 181.395000 ;
        RECT 69.590000 181.595000 69.790000 181.795000 ;
        RECT 69.590000 181.995000 69.790000 182.195000 ;
        RECT 69.590000 182.395000 69.790000 182.595000 ;
        RECT 69.590000 182.795000 69.790000 182.995000 ;
        RECT 69.590000 183.195000 69.790000 183.395000 ;
        RECT 69.590000 183.595000 69.790000 183.795000 ;
        RECT 69.590000 183.995000 69.790000 184.195000 ;
        RECT 69.590000 184.395000 69.790000 184.595000 ;
        RECT 69.590000 184.795000 69.790000 184.995000 ;
        RECT 69.590000 185.195000 69.790000 185.395000 ;
        RECT 69.590000 185.595000 69.790000 185.795000 ;
        RECT 69.590000 185.995000 69.790000 186.195000 ;
        RECT 69.590000 186.395000 69.790000 186.595000 ;
        RECT 69.590000 186.795000 69.790000 186.995000 ;
        RECT 69.590000 187.195000 69.790000 187.395000 ;
        RECT 69.590000 187.595000 69.790000 187.795000 ;
        RECT 69.590000 187.995000 69.790000 188.195000 ;
        RECT 69.590000 188.395000 69.790000 188.595000 ;
        RECT 69.590000 188.795000 69.790000 188.995000 ;
        RECT 69.590000 189.195000 69.790000 189.395000 ;
        RECT 69.590000 189.595000 69.790000 189.795000 ;
        RECT 69.590000 189.995000 69.790000 190.195000 ;
        RECT 69.590000 190.395000 69.790000 190.595000 ;
        RECT 69.590000 190.795000 69.790000 190.995000 ;
        RECT 69.590000 191.195000 69.790000 191.395000 ;
        RECT 69.590000 191.595000 69.790000 191.795000 ;
        RECT 69.590000 191.995000 69.790000 192.195000 ;
        RECT 69.590000 192.395000 69.790000 192.595000 ;
        RECT 69.590000 192.795000 69.790000 192.995000 ;
        RECT 69.590000 193.195000 69.790000 193.395000 ;
        RECT 69.590000 193.595000 69.790000 193.795000 ;
        RECT 69.590000 193.995000 69.790000 194.195000 ;
        RECT 69.590000 194.395000 69.790000 194.595000 ;
        RECT 69.590000 194.795000 69.790000 194.995000 ;
        RECT 69.590000 195.200000 69.790000 195.400000 ;
        RECT 69.590000 195.605000 69.790000 195.805000 ;
        RECT 69.590000 196.010000 69.790000 196.210000 ;
        RECT 69.590000 196.415000 69.790000 196.615000 ;
        RECT 69.590000 196.820000 69.790000 197.020000 ;
        RECT 69.590000 197.225000 69.790000 197.425000 ;
        RECT 69.590000 197.630000 69.790000 197.830000 ;
        RECT 69.590000 198.035000 69.790000 198.235000 ;
        RECT 69.590000 198.440000 69.790000 198.640000 ;
        RECT 69.590000 198.845000 69.790000 199.045000 ;
        RECT 69.590000 199.250000 69.790000 199.450000 ;
        RECT 69.590000 199.655000 69.790000 199.855000 ;
        RECT 69.950000  25.910000 70.150000  26.110000 ;
        RECT 69.950000  26.340000 70.150000  26.540000 ;
        RECT 69.950000  26.770000 70.150000  26.970000 ;
        RECT 69.950000  27.200000 70.150000  27.400000 ;
        RECT 69.950000  27.630000 70.150000  27.830000 ;
        RECT 69.950000  28.060000 70.150000  28.260000 ;
        RECT 69.950000  28.490000 70.150000  28.690000 ;
        RECT 69.950000  28.920000 70.150000  29.120000 ;
        RECT 69.950000  29.350000 70.150000  29.550000 ;
        RECT 69.950000  29.780000 70.150000  29.980000 ;
        RECT 69.950000  30.210000 70.150000  30.410000 ;
        RECT 69.990000 175.995000 70.190000 176.195000 ;
        RECT 69.990000 176.395000 70.190000 176.595000 ;
        RECT 69.990000 176.795000 70.190000 176.995000 ;
        RECT 69.990000 177.195000 70.190000 177.395000 ;
        RECT 69.990000 177.595000 70.190000 177.795000 ;
        RECT 69.990000 177.995000 70.190000 178.195000 ;
        RECT 69.990000 178.395000 70.190000 178.595000 ;
        RECT 69.990000 178.795000 70.190000 178.995000 ;
        RECT 69.990000 179.195000 70.190000 179.395000 ;
        RECT 69.990000 179.595000 70.190000 179.795000 ;
        RECT 69.990000 179.995000 70.190000 180.195000 ;
        RECT 69.990000 180.395000 70.190000 180.595000 ;
        RECT 69.990000 180.795000 70.190000 180.995000 ;
        RECT 69.990000 181.195000 70.190000 181.395000 ;
        RECT 69.990000 181.595000 70.190000 181.795000 ;
        RECT 69.990000 181.995000 70.190000 182.195000 ;
        RECT 69.990000 182.395000 70.190000 182.595000 ;
        RECT 69.990000 182.795000 70.190000 182.995000 ;
        RECT 69.990000 183.195000 70.190000 183.395000 ;
        RECT 69.990000 183.595000 70.190000 183.795000 ;
        RECT 69.990000 183.995000 70.190000 184.195000 ;
        RECT 69.990000 184.395000 70.190000 184.595000 ;
        RECT 69.990000 184.795000 70.190000 184.995000 ;
        RECT 69.990000 185.195000 70.190000 185.395000 ;
        RECT 69.990000 185.595000 70.190000 185.795000 ;
        RECT 69.990000 185.995000 70.190000 186.195000 ;
        RECT 69.990000 186.395000 70.190000 186.595000 ;
        RECT 69.990000 186.795000 70.190000 186.995000 ;
        RECT 69.990000 187.195000 70.190000 187.395000 ;
        RECT 69.990000 187.595000 70.190000 187.795000 ;
        RECT 69.990000 187.995000 70.190000 188.195000 ;
        RECT 69.990000 188.395000 70.190000 188.595000 ;
        RECT 69.990000 188.795000 70.190000 188.995000 ;
        RECT 69.990000 189.195000 70.190000 189.395000 ;
        RECT 69.990000 189.595000 70.190000 189.795000 ;
        RECT 69.990000 189.995000 70.190000 190.195000 ;
        RECT 69.990000 190.395000 70.190000 190.595000 ;
        RECT 69.990000 190.795000 70.190000 190.995000 ;
        RECT 69.990000 191.195000 70.190000 191.395000 ;
        RECT 69.990000 191.595000 70.190000 191.795000 ;
        RECT 69.990000 191.995000 70.190000 192.195000 ;
        RECT 69.990000 192.395000 70.190000 192.595000 ;
        RECT 69.990000 192.795000 70.190000 192.995000 ;
        RECT 69.990000 193.195000 70.190000 193.395000 ;
        RECT 69.990000 193.595000 70.190000 193.795000 ;
        RECT 69.990000 193.995000 70.190000 194.195000 ;
        RECT 69.990000 194.395000 70.190000 194.595000 ;
        RECT 69.990000 194.795000 70.190000 194.995000 ;
        RECT 69.990000 195.200000 70.190000 195.400000 ;
        RECT 69.990000 195.605000 70.190000 195.805000 ;
        RECT 69.990000 196.010000 70.190000 196.210000 ;
        RECT 69.990000 196.415000 70.190000 196.615000 ;
        RECT 69.990000 196.820000 70.190000 197.020000 ;
        RECT 69.990000 197.225000 70.190000 197.425000 ;
        RECT 69.990000 197.630000 70.190000 197.830000 ;
        RECT 69.990000 198.035000 70.190000 198.235000 ;
        RECT 69.990000 198.440000 70.190000 198.640000 ;
        RECT 69.990000 198.845000 70.190000 199.045000 ;
        RECT 69.990000 199.250000 70.190000 199.450000 ;
        RECT 69.990000 199.655000 70.190000 199.855000 ;
        RECT 70.355000  25.910000 70.555000  26.110000 ;
        RECT 70.355000  26.340000 70.555000  26.540000 ;
        RECT 70.355000  26.770000 70.555000  26.970000 ;
        RECT 70.355000  27.200000 70.555000  27.400000 ;
        RECT 70.355000  27.630000 70.555000  27.830000 ;
        RECT 70.355000  28.060000 70.555000  28.260000 ;
        RECT 70.355000  28.490000 70.555000  28.690000 ;
        RECT 70.355000  28.920000 70.555000  29.120000 ;
        RECT 70.355000  29.350000 70.555000  29.550000 ;
        RECT 70.355000  29.780000 70.555000  29.980000 ;
        RECT 70.355000  30.210000 70.555000  30.410000 ;
        RECT 70.390000 175.995000 70.590000 176.195000 ;
        RECT 70.390000 176.395000 70.590000 176.595000 ;
        RECT 70.390000 176.795000 70.590000 176.995000 ;
        RECT 70.390000 177.195000 70.590000 177.395000 ;
        RECT 70.390000 177.595000 70.590000 177.795000 ;
        RECT 70.390000 177.995000 70.590000 178.195000 ;
        RECT 70.390000 178.395000 70.590000 178.595000 ;
        RECT 70.390000 178.795000 70.590000 178.995000 ;
        RECT 70.390000 179.195000 70.590000 179.395000 ;
        RECT 70.390000 179.595000 70.590000 179.795000 ;
        RECT 70.390000 179.995000 70.590000 180.195000 ;
        RECT 70.390000 180.395000 70.590000 180.595000 ;
        RECT 70.390000 180.795000 70.590000 180.995000 ;
        RECT 70.390000 181.195000 70.590000 181.395000 ;
        RECT 70.390000 181.595000 70.590000 181.795000 ;
        RECT 70.390000 181.995000 70.590000 182.195000 ;
        RECT 70.390000 182.395000 70.590000 182.595000 ;
        RECT 70.390000 182.795000 70.590000 182.995000 ;
        RECT 70.390000 183.195000 70.590000 183.395000 ;
        RECT 70.390000 183.595000 70.590000 183.795000 ;
        RECT 70.390000 183.995000 70.590000 184.195000 ;
        RECT 70.390000 184.395000 70.590000 184.595000 ;
        RECT 70.390000 184.795000 70.590000 184.995000 ;
        RECT 70.390000 185.195000 70.590000 185.395000 ;
        RECT 70.390000 185.595000 70.590000 185.795000 ;
        RECT 70.390000 185.995000 70.590000 186.195000 ;
        RECT 70.390000 186.395000 70.590000 186.595000 ;
        RECT 70.390000 186.795000 70.590000 186.995000 ;
        RECT 70.390000 187.195000 70.590000 187.395000 ;
        RECT 70.390000 187.595000 70.590000 187.795000 ;
        RECT 70.390000 187.995000 70.590000 188.195000 ;
        RECT 70.390000 188.395000 70.590000 188.595000 ;
        RECT 70.390000 188.795000 70.590000 188.995000 ;
        RECT 70.390000 189.195000 70.590000 189.395000 ;
        RECT 70.390000 189.595000 70.590000 189.795000 ;
        RECT 70.390000 189.995000 70.590000 190.195000 ;
        RECT 70.390000 190.395000 70.590000 190.595000 ;
        RECT 70.390000 190.795000 70.590000 190.995000 ;
        RECT 70.390000 191.195000 70.590000 191.395000 ;
        RECT 70.390000 191.595000 70.590000 191.795000 ;
        RECT 70.390000 191.995000 70.590000 192.195000 ;
        RECT 70.390000 192.395000 70.590000 192.595000 ;
        RECT 70.390000 192.795000 70.590000 192.995000 ;
        RECT 70.390000 193.195000 70.590000 193.395000 ;
        RECT 70.390000 193.595000 70.590000 193.795000 ;
        RECT 70.390000 193.995000 70.590000 194.195000 ;
        RECT 70.390000 194.395000 70.590000 194.595000 ;
        RECT 70.390000 194.795000 70.590000 194.995000 ;
        RECT 70.390000 195.200000 70.590000 195.400000 ;
        RECT 70.390000 195.605000 70.590000 195.805000 ;
        RECT 70.390000 196.010000 70.590000 196.210000 ;
        RECT 70.390000 196.415000 70.590000 196.615000 ;
        RECT 70.390000 196.820000 70.590000 197.020000 ;
        RECT 70.390000 197.225000 70.590000 197.425000 ;
        RECT 70.390000 197.630000 70.590000 197.830000 ;
        RECT 70.390000 198.035000 70.590000 198.235000 ;
        RECT 70.390000 198.440000 70.590000 198.640000 ;
        RECT 70.390000 198.845000 70.590000 199.045000 ;
        RECT 70.390000 199.250000 70.590000 199.450000 ;
        RECT 70.390000 199.655000 70.590000 199.855000 ;
        RECT 70.760000  25.910000 70.960000  26.110000 ;
        RECT 70.760000  26.340000 70.960000  26.540000 ;
        RECT 70.760000  26.770000 70.960000  26.970000 ;
        RECT 70.760000  27.200000 70.960000  27.400000 ;
        RECT 70.760000  27.630000 70.960000  27.830000 ;
        RECT 70.760000  28.060000 70.960000  28.260000 ;
        RECT 70.760000  28.490000 70.960000  28.690000 ;
        RECT 70.760000  28.920000 70.960000  29.120000 ;
        RECT 70.760000  29.350000 70.960000  29.550000 ;
        RECT 70.760000  29.780000 70.960000  29.980000 ;
        RECT 70.760000  30.210000 70.960000  30.410000 ;
        RECT 70.790000 175.995000 70.990000 176.195000 ;
        RECT 70.790000 176.395000 70.990000 176.595000 ;
        RECT 70.790000 176.795000 70.990000 176.995000 ;
        RECT 70.790000 177.195000 70.990000 177.395000 ;
        RECT 70.790000 177.595000 70.990000 177.795000 ;
        RECT 70.790000 177.995000 70.990000 178.195000 ;
        RECT 70.790000 178.395000 70.990000 178.595000 ;
        RECT 70.790000 178.795000 70.990000 178.995000 ;
        RECT 70.790000 179.195000 70.990000 179.395000 ;
        RECT 70.790000 179.595000 70.990000 179.795000 ;
        RECT 70.790000 179.995000 70.990000 180.195000 ;
        RECT 70.790000 180.395000 70.990000 180.595000 ;
        RECT 70.790000 180.795000 70.990000 180.995000 ;
        RECT 70.790000 181.195000 70.990000 181.395000 ;
        RECT 70.790000 181.595000 70.990000 181.795000 ;
        RECT 70.790000 181.995000 70.990000 182.195000 ;
        RECT 70.790000 182.395000 70.990000 182.595000 ;
        RECT 70.790000 182.795000 70.990000 182.995000 ;
        RECT 70.790000 183.195000 70.990000 183.395000 ;
        RECT 70.790000 183.595000 70.990000 183.795000 ;
        RECT 70.790000 183.995000 70.990000 184.195000 ;
        RECT 70.790000 184.395000 70.990000 184.595000 ;
        RECT 70.790000 184.795000 70.990000 184.995000 ;
        RECT 70.790000 185.195000 70.990000 185.395000 ;
        RECT 70.790000 185.595000 70.990000 185.795000 ;
        RECT 70.790000 185.995000 70.990000 186.195000 ;
        RECT 70.790000 186.395000 70.990000 186.595000 ;
        RECT 70.790000 186.795000 70.990000 186.995000 ;
        RECT 70.790000 187.195000 70.990000 187.395000 ;
        RECT 70.790000 187.595000 70.990000 187.795000 ;
        RECT 70.790000 187.995000 70.990000 188.195000 ;
        RECT 70.790000 188.395000 70.990000 188.595000 ;
        RECT 70.790000 188.795000 70.990000 188.995000 ;
        RECT 70.790000 189.195000 70.990000 189.395000 ;
        RECT 70.790000 189.595000 70.990000 189.795000 ;
        RECT 70.790000 189.995000 70.990000 190.195000 ;
        RECT 70.790000 190.395000 70.990000 190.595000 ;
        RECT 70.790000 190.795000 70.990000 190.995000 ;
        RECT 70.790000 191.195000 70.990000 191.395000 ;
        RECT 70.790000 191.595000 70.990000 191.795000 ;
        RECT 70.790000 191.995000 70.990000 192.195000 ;
        RECT 70.790000 192.395000 70.990000 192.595000 ;
        RECT 70.790000 192.795000 70.990000 192.995000 ;
        RECT 70.790000 193.195000 70.990000 193.395000 ;
        RECT 70.790000 193.595000 70.990000 193.795000 ;
        RECT 70.790000 193.995000 70.990000 194.195000 ;
        RECT 70.790000 194.395000 70.990000 194.595000 ;
        RECT 70.790000 194.795000 70.990000 194.995000 ;
        RECT 70.790000 195.200000 70.990000 195.400000 ;
        RECT 70.790000 195.605000 70.990000 195.805000 ;
        RECT 70.790000 196.010000 70.990000 196.210000 ;
        RECT 70.790000 196.415000 70.990000 196.615000 ;
        RECT 70.790000 196.820000 70.990000 197.020000 ;
        RECT 70.790000 197.225000 70.990000 197.425000 ;
        RECT 70.790000 197.630000 70.990000 197.830000 ;
        RECT 70.790000 198.035000 70.990000 198.235000 ;
        RECT 70.790000 198.440000 70.990000 198.640000 ;
        RECT 70.790000 198.845000 70.990000 199.045000 ;
        RECT 70.790000 199.250000 70.990000 199.450000 ;
        RECT 70.790000 199.655000 70.990000 199.855000 ;
        RECT 71.165000  25.910000 71.365000  26.110000 ;
        RECT 71.165000  26.340000 71.365000  26.540000 ;
        RECT 71.165000  26.770000 71.365000  26.970000 ;
        RECT 71.165000  27.200000 71.365000  27.400000 ;
        RECT 71.165000  27.630000 71.365000  27.830000 ;
        RECT 71.165000  28.060000 71.365000  28.260000 ;
        RECT 71.165000  28.490000 71.365000  28.690000 ;
        RECT 71.165000  28.920000 71.365000  29.120000 ;
        RECT 71.165000  29.350000 71.365000  29.550000 ;
        RECT 71.165000  29.780000 71.365000  29.980000 ;
        RECT 71.165000  30.210000 71.365000  30.410000 ;
        RECT 71.190000 175.995000 71.390000 176.195000 ;
        RECT 71.190000 176.395000 71.390000 176.595000 ;
        RECT 71.190000 176.795000 71.390000 176.995000 ;
        RECT 71.190000 177.195000 71.390000 177.395000 ;
        RECT 71.190000 177.595000 71.390000 177.795000 ;
        RECT 71.190000 177.995000 71.390000 178.195000 ;
        RECT 71.190000 178.395000 71.390000 178.595000 ;
        RECT 71.190000 178.795000 71.390000 178.995000 ;
        RECT 71.190000 179.195000 71.390000 179.395000 ;
        RECT 71.190000 179.595000 71.390000 179.795000 ;
        RECT 71.190000 179.995000 71.390000 180.195000 ;
        RECT 71.190000 180.395000 71.390000 180.595000 ;
        RECT 71.190000 180.795000 71.390000 180.995000 ;
        RECT 71.190000 181.195000 71.390000 181.395000 ;
        RECT 71.190000 181.595000 71.390000 181.795000 ;
        RECT 71.190000 181.995000 71.390000 182.195000 ;
        RECT 71.190000 182.395000 71.390000 182.595000 ;
        RECT 71.190000 182.795000 71.390000 182.995000 ;
        RECT 71.190000 183.195000 71.390000 183.395000 ;
        RECT 71.190000 183.595000 71.390000 183.795000 ;
        RECT 71.190000 183.995000 71.390000 184.195000 ;
        RECT 71.190000 184.395000 71.390000 184.595000 ;
        RECT 71.190000 184.795000 71.390000 184.995000 ;
        RECT 71.190000 185.195000 71.390000 185.395000 ;
        RECT 71.190000 185.595000 71.390000 185.795000 ;
        RECT 71.190000 185.995000 71.390000 186.195000 ;
        RECT 71.190000 186.395000 71.390000 186.595000 ;
        RECT 71.190000 186.795000 71.390000 186.995000 ;
        RECT 71.190000 187.195000 71.390000 187.395000 ;
        RECT 71.190000 187.595000 71.390000 187.795000 ;
        RECT 71.190000 187.995000 71.390000 188.195000 ;
        RECT 71.190000 188.395000 71.390000 188.595000 ;
        RECT 71.190000 188.795000 71.390000 188.995000 ;
        RECT 71.190000 189.195000 71.390000 189.395000 ;
        RECT 71.190000 189.595000 71.390000 189.795000 ;
        RECT 71.190000 189.995000 71.390000 190.195000 ;
        RECT 71.190000 190.395000 71.390000 190.595000 ;
        RECT 71.190000 190.795000 71.390000 190.995000 ;
        RECT 71.190000 191.195000 71.390000 191.395000 ;
        RECT 71.190000 191.595000 71.390000 191.795000 ;
        RECT 71.190000 191.995000 71.390000 192.195000 ;
        RECT 71.190000 192.395000 71.390000 192.595000 ;
        RECT 71.190000 192.795000 71.390000 192.995000 ;
        RECT 71.190000 193.195000 71.390000 193.395000 ;
        RECT 71.190000 193.595000 71.390000 193.795000 ;
        RECT 71.190000 193.995000 71.390000 194.195000 ;
        RECT 71.190000 194.395000 71.390000 194.595000 ;
        RECT 71.190000 194.795000 71.390000 194.995000 ;
        RECT 71.190000 195.200000 71.390000 195.400000 ;
        RECT 71.190000 195.605000 71.390000 195.805000 ;
        RECT 71.190000 196.010000 71.390000 196.210000 ;
        RECT 71.190000 196.415000 71.390000 196.615000 ;
        RECT 71.190000 196.820000 71.390000 197.020000 ;
        RECT 71.190000 197.225000 71.390000 197.425000 ;
        RECT 71.190000 197.630000 71.390000 197.830000 ;
        RECT 71.190000 198.035000 71.390000 198.235000 ;
        RECT 71.190000 198.440000 71.390000 198.640000 ;
        RECT 71.190000 198.845000 71.390000 199.045000 ;
        RECT 71.190000 199.250000 71.390000 199.450000 ;
        RECT 71.190000 199.655000 71.390000 199.855000 ;
        RECT 71.570000  25.910000 71.770000  26.110000 ;
        RECT 71.570000  26.340000 71.770000  26.540000 ;
        RECT 71.570000  26.770000 71.770000  26.970000 ;
        RECT 71.570000  27.200000 71.770000  27.400000 ;
        RECT 71.570000  27.630000 71.770000  27.830000 ;
        RECT 71.570000  28.060000 71.770000  28.260000 ;
        RECT 71.570000  28.490000 71.770000  28.690000 ;
        RECT 71.570000  28.920000 71.770000  29.120000 ;
        RECT 71.570000  29.350000 71.770000  29.550000 ;
        RECT 71.570000  29.780000 71.770000  29.980000 ;
        RECT 71.570000  30.210000 71.770000  30.410000 ;
        RECT 71.590000 175.995000 71.790000 176.195000 ;
        RECT 71.590000 176.395000 71.790000 176.595000 ;
        RECT 71.590000 176.795000 71.790000 176.995000 ;
        RECT 71.590000 177.195000 71.790000 177.395000 ;
        RECT 71.590000 177.595000 71.790000 177.795000 ;
        RECT 71.590000 177.995000 71.790000 178.195000 ;
        RECT 71.590000 178.395000 71.790000 178.595000 ;
        RECT 71.590000 178.795000 71.790000 178.995000 ;
        RECT 71.590000 179.195000 71.790000 179.395000 ;
        RECT 71.590000 179.595000 71.790000 179.795000 ;
        RECT 71.590000 179.995000 71.790000 180.195000 ;
        RECT 71.590000 180.395000 71.790000 180.595000 ;
        RECT 71.590000 180.795000 71.790000 180.995000 ;
        RECT 71.590000 181.195000 71.790000 181.395000 ;
        RECT 71.590000 181.595000 71.790000 181.795000 ;
        RECT 71.590000 181.995000 71.790000 182.195000 ;
        RECT 71.590000 182.395000 71.790000 182.595000 ;
        RECT 71.590000 182.795000 71.790000 182.995000 ;
        RECT 71.590000 183.195000 71.790000 183.395000 ;
        RECT 71.590000 183.595000 71.790000 183.795000 ;
        RECT 71.590000 183.995000 71.790000 184.195000 ;
        RECT 71.590000 184.395000 71.790000 184.595000 ;
        RECT 71.590000 184.795000 71.790000 184.995000 ;
        RECT 71.590000 185.195000 71.790000 185.395000 ;
        RECT 71.590000 185.595000 71.790000 185.795000 ;
        RECT 71.590000 185.995000 71.790000 186.195000 ;
        RECT 71.590000 186.395000 71.790000 186.595000 ;
        RECT 71.590000 186.795000 71.790000 186.995000 ;
        RECT 71.590000 187.195000 71.790000 187.395000 ;
        RECT 71.590000 187.595000 71.790000 187.795000 ;
        RECT 71.590000 187.995000 71.790000 188.195000 ;
        RECT 71.590000 188.395000 71.790000 188.595000 ;
        RECT 71.590000 188.795000 71.790000 188.995000 ;
        RECT 71.590000 189.195000 71.790000 189.395000 ;
        RECT 71.590000 189.595000 71.790000 189.795000 ;
        RECT 71.590000 189.995000 71.790000 190.195000 ;
        RECT 71.590000 190.395000 71.790000 190.595000 ;
        RECT 71.590000 190.795000 71.790000 190.995000 ;
        RECT 71.590000 191.195000 71.790000 191.395000 ;
        RECT 71.590000 191.595000 71.790000 191.795000 ;
        RECT 71.590000 191.995000 71.790000 192.195000 ;
        RECT 71.590000 192.395000 71.790000 192.595000 ;
        RECT 71.590000 192.795000 71.790000 192.995000 ;
        RECT 71.590000 193.195000 71.790000 193.395000 ;
        RECT 71.590000 193.595000 71.790000 193.795000 ;
        RECT 71.590000 193.995000 71.790000 194.195000 ;
        RECT 71.590000 194.395000 71.790000 194.595000 ;
        RECT 71.590000 194.795000 71.790000 194.995000 ;
        RECT 71.590000 195.200000 71.790000 195.400000 ;
        RECT 71.590000 195.605000 71.790000 195.805000 ;
        RECT 71.590000 196.010000 71.790000 196.210000 ;
        RECT 71.590000 196.415000 71.790000 196.615000 ;
        RECT 71.590000 196.820000 71.790000 197.020000 ;
        RECT 71.590000 197.225000 71.790000 197.425000 ;
        RECT 71.590000 197.630000 71.790000 197.830000 ;
        RECT 71.590000 198.035000 71.790000 198.235000 ;
        RECT 71.590000 198.440000 71.790000 198.640000 ;
        RECT 71.590000 198.845000 71.790000 199.045000 ;
        RECT 71.590000 199.250000 71.790000 199.450000 ;
        RECT 71.590000 199.655000 71.790000 199.855000 ;
        RECT 71.975000  25.910000 72.175000  26.110000 ;
        RECT 71.975000  26.340000 72.175000  26.540000 ;
        RECT 71.975000  26.770000 72.175000  26.970000 ;
        RECT 71.975000  27.200000 72.175000  27.400000 ;
        RECT 71.975000  27.630000 72.175000  27.830000 ;
        RECT 71.975000  28.060000 72.175000  28.260000 ;
        RECT 71.975000  28.490000 72.175000  28.690000 ;
        RECT 71.975000  28.920000 72.175000  29.120000 ;
        RECT 71.975000  29.350000 72.175000  29.550000 ;
        RECT 71.975000  29.780000 72.175000  29.980000 ;
        RECT 71.975000  30.210000 72.175000  30.410000 ;
        RECT 71.990000 175.995000 72.190000 176.195000 ;
        RECT 71.990000 176.395000 72.190000 176.595000 ;
        RECT 71.990000 176.795000 72.190000 176.995000 ;
        RECT 71.990000 177.195000 72.190000 177.395000 ;
        RECT 71.990000 177.595000 72.190000 177.795000 ;
        RECT 71.990000 177.995000 72.190000 178.195000 ;
        RECT 71.990000 178.395000 72.190000 178.595000 ;
        RECT 71.990000 178.795000 72.190000 178.995000 ;
        RECT 71.990000 179.195000 72.190000 179.395000 ;
        RECT 71.990000 179.595000 72.190000 179.795000 ;
        RECT 71.990000 179.995000 72.190000 180.195000 ;
        RECT 71.990000 180.395000 72.190000 180.595000 ;
        RECT 71.990000 180.795000 72.190000 180.995000 ;
        RECT 71.990000 181.195000 72.190000 181.395000 ;
        RECT 71.990000 181.595000 72.190000 181.795000 ;
        RECT 71.990000 181.995000 72.190000 182.195000 ;
        RECT 71.990000 182.395000 72.190000 182.595000 ;
        RECT 71.990000 182.795000 72.190000 182.995000 ;
        RECT 71.990000 183.195000 72.190000 183.395000 ;
        RECT 71.990000 183.595000 72.190000 183.795000 ;
        RECT 71.990000 183.995000 72.190000 184.195000 ;
        RECT 71.990000 184.395000 72.190000 184.595000 ;
        RECT 71.990000 184.795000 72.190000 184.995000 ;
        RECT 71.990000 185.195000 72.190000 185.395000 ;
        RECT 71.990000 185.595000 72.190000 185.795000 ;
        RECT 71.990000 185.995000 72.190000 186.195000 ;
        RECT 71.990000 186.395000 72.190000 186.595000 ;
        RECT 71.990000 186.795000 72.190000 186.995000 ;
        RECT 71.990000 187.195000 72.190000 187.395000 ;
        RECT 71.990000 187.595000 72.190000 187.795000 ;
        RECT 71.990000 187.995000 72.190000 188.195000 ;
        RECT 71.990000 188.395000 72.190000 188.595000 ;
        RECT 71.990000 188.795000 72.190000 188.995000 ;
        RECT 71.990000 189.195000 72.190000 189.395000 ;
        RECT 71.990000 189.595000 72.190000 189.795000 ;
        RECT 71.990000 189.995000 72.190000 190.195000 ;
        RECT 71.990000 190.395000 72.190000 190.595000 ;
        RECT 71.990000 190.795000 72.190000 190.995000 ;
        RECT 71.990000 191.195000 72.190000 191.395000 ;
        RECT 71.990000 191.595000 72.190000 191.795000 ;
        RECT 71.990000 191.995000 72.190000 192.195000 ;
        RECT 71.990000 192.395000 72.190000 192.595000 ;
        RECT 71.990000 192.795000 72.190000 192.995000 ;
        RECT 71.990000 193.195000 72.190000 193.395000 ;
        RECT 71.990000 193.595000 72.190000 193.795000 ;
        RECT 71.990000 193.995000 72.190000 194.195000 ;
        RECT 71.990000 194.395000 72.190000 194.595000 ;
        RECT 71.990000 194.795000 72.190000 194.995000 ;
        RECT 71.990000 195.200000 72.190000 195.400000 ;
        RECT 71.990000 195.605000 72.190000 195.805000 ;
        RECT 71.990000 196.010000 72.190000 196.210000 ;
        RECT 71.990000 196.415000 72.190000 196.615000 ;
        RECT 71.990000 196.820000 72.190000 197.020000 ;
        RECT 71.990000 197.225000 72.190000 197.425000 ;
        RECT 71.990000 197.630000 72.190000 197.830000 ;
        RECT 71.990000 198.035000 72.190000 198.235000 ;
        RECT 71.990000 198.440000 72.190000 198.640000 ;
        RECT 71.990000 198.845000 72.190000 199.045000 ;
        RECT 71.990000 199.250000 72.190000 199.450000 ;
        RECT 71.990000 199.655000 72.190000 199.855000 ;
        RECT 72.380000  25.910000 72.580000  26.110000 ;
        RECT 72.380000  26.340000 72.580000  26.540000 ;
        RECT 72.380000  26.770000 72.580000  26.970000 ;
        RECT 72.380000  27.200000 72.580000  27.400000 ;
        RECT 72.380000  27.630000 72.580000  27.830000 ;
        RECT 72.380000  28.060000 72.580000  28.260000 ;
        RECT 72.380000  28.490000 72.580000  28.690000 ;
        RECT 72.380000  28.920000 72.580000  29.120000 ;
        RECT 72.380000  29.350000 72.580000  29.550000 ;
        RECT 72.380000  29.780000 72.580000  29.980000 ;
        RECT 72.380000  30.210000 72.580000  30.410000 ;
        RECT 72.390000 175.995000 72.590000 176.195000 ;
        RECT 72.390000 176.395000 72.590000 176.595000 ;
        RECT 72.390000 176.795000 72.590000 176.995000 ;
        RECT 72.390000 177.195000 72.590000 177.395000 ;
        RECT 72.390000 177.595000 72.590000 177.795000 ;
        RECT 72.390000 177.995000 72.590000 178.195000 ;
        RECT 72.390000 178.395000 72.590000 178.595000 ;
        RECT 72.390000 178.795000 72.590000 178.995000 ;
        RECT 72.390000 179.195000 72.590000 179.395000 ;
        RECT 72.390000 179.595000 72.590000 179.795000 ;
        RECT 72.390000 179.995000 72.590000 180.195000 ;
        RECT 72.390000 180.395000 72.590000 180.595000 ;
        RECT 72.390000 180.795000 72.590000 180.995000 ;
        RECT 72.390000 181.195000 72.590000 181.395000 ;
        RECT 72.390000 181.595000 72.590000 181.795000 ;
        RECT 72.390000 181.995000 72.590000 182.195000 ;
        RECT 72.390000 182.395000 72.590000 182.595000 ;
        RECT 72.390000 182.795000 72.590000 182.995000 ;
        RECT 72.390000 183.195000 72.590000 183.395000 ;
        RECT 72.390000 183.595000 72.590000 183.795000 ;
        RECT 72.390000 183.995000 72.590000 184.195000 ;
        RECT 72.390000 184.395000 72.590000 184.595000 ;
        RECT 72.390000 184.795000 72.590000 184.995000 ;
        RECT 72.390000 185.195000 72.590000 185.395000 ;
        RECT 72.390000 185.595000 72.590000 185.795000 ;
        RECT 72.390000 185.995000 72.590000 186.195000 ;
        RECT 72.390000 186.395000 72.590000 186.595000 ;
        RECT 72.390000 186.795000 72.590000 186.995000 ;
        RECT 72.390000 187.195000 72.590000 187.395000 ;
        RECT 72.390000 187.595000 72.590000 187.795000 ;
        RECT 72.390000 187.995000 72.590000 188.195000 ;
        RECT 72.390000 188.395000 72.590000 188.595000 ;
        RECT 72.390000 188.795000 72.590000 188.995000 ;
        RECT 72.390000 189.195000 72.590000 189.395000 ;
        RECT 72.390000 189.595000 72.590000 189.795000 ;
        RECT 72.390000 189.995000 72.590000 190.195000 ;
        RECT 72.390000 190.395000 72.590000 190.595000 ;
        RECT 72.390000 190.795000 72.590000 190.995000 ;
        RECT 72.390000 191.195000 72.590000 191.395000 ;
        RECT 72.390000 191.595000 72.590000 191.795000 ;
        RECT 72.390000 191.995000 72.590000 192.195000 ;
        RECT 72.390000 192.395000 72.590000 192.595000 ;
        RECT 72.390000 192.795000 72.590000 192.995000 ;
        RECT 72.390000 193.195000 72.590000 193.395000 ;
        RECT 72.390000 193.595000 72.590000 193.795000 ;
        RECT 72.390000 193.995000 72.590000 194.195000 ;
        RECT 72.390000 194.395000 72.590000 194.595000 ;
        RECT 72.390000 194.795000 72.590000 194.995000 ;
        RECT 72.390000 195.200000 72.590000 195.400000 ;
        RECT 72.390000 195.605000 72.590000 195.805000 ;
        RECT 72.390000 196.010000 72.590000 196.210000 ;
        RECT 72.390000 196.415000 72.590000 196.615000 ;
        RECT 72.390000 196.820000 72.590000 197.020000 ;
        RECT 72.390000 197.225000 72.590000 197.425000 ;
        RECT 72.390000 197.630000 72.590000 197.830000 ;
        RECT 72.390000 198.035000 72.590000 198.235000 ;
        RECT 72.390000 198.440000 72.590000 198.640000 ;
        RECT 72.390000 198.845000 72.590000 199.045000 ;
        RECT 72.390000 199.250000 72.590000 199.450000 ;
        RECT 72.390000 199.655000 72.590000 199.855000 ;
        RECT 72.785000  25.910000 72.985000  26.110000 ;
        RECT 72.785000  26.340000 72.985000  26.540000 ;
        RECT 72.785000  26.770000 72.985000  26.970000 ;
        RECT 72.785000  27.200000 72.985000  27.400000 ;
        RECT 72.785000  27.630000 72.985000  27.830000 ;
        RECT 72.785000  28.060000 72.985000  28.260000 ;
        RECT 72.785000  28.490000 72.985000  28.690000 ;
        RECT 72.785000  28.920000 72.985000  29.120000 ;
        RECT 72.785000  29.350000 72.985000  29.550000 ;
        RECT 72.785000  29.780000 72.985000  29.980000 ;
        RECT 72.785000  30.210000 72.985000  30.410000 ;
        RECT 72.790000 175.995000 72.990000 176.195000 ;
        RECT 72.790000 176.395000 72.990000 176.595000 ;
        RECT 72.790000 176.795000 72.990000 176.995000 ;
        RECT 72.790000 177.195000 72.990000 177.395000 ;
        RECT 72.790000 177.595000 72.990000 177.795000 ;
        RECT 72.790000 177.995000 72.990000 178.195000 ;
        RECT 72.790000 178.395000 72.990000 178.595000 ;
        RECT 72.790000 178.795000 72.990000 178.995000 ;
        RECT 72.790000 179.195000 72.990000 179.395000 ;
        RECT 72.790000 179.595000 72.990000 179.795000 ;
        RECT 72.790000 179.995000 72.990000 180.195000 ;
        RECT 72.790000 180.395000 72.990000 180.595000 ;
        RECT 72.790000 180.795000 72.990000 180.995000 ;
        RECT 72.790000 181.195000 72.990000 181.395000 ;
        RECT 72.790000 181.595000 72.990000 181.795000 ;
        RECT 72.790000 181.995000 72.990000 182.195000 ;
        RECT 72.790000 182.395000 72.990000 182.595000 ;
        RECT 72.790000 182.795000 72.990000 182.995000 ;
        RECT 72.790000 183.195000 72.990000 183.395000 ;
        RECT 72.790000 183.595000 72.990000 183.795000 ;
        RECT 72.790000 183.995000 72.990000 184.195000 ;
        RECT 72.790000 184.395000 72.990000 184.595000 ;
        RECT 72.790000 184.795000 72.990000 184.995000 ;
        RECT 72.790000 185.195000 72.990000 185.395000 ;
        RECT 72.790000 185.595000 72.990000 185.795000 ;
        RECT 72.790000 185.995000 72.990000 186.195000 ;
        RECT 72.790000 186.395000 72.990000 186.595000 ;
        RECT 72.790000 186.795000 72.990000 186.995000 ;
        RECT 72.790000 187.195000 72.990000 187.395000 ;
        RECT 72.790000 187.595000 72.990000 187.795000 ;
        RECT 72.790000 187.995000 72.990000 188.195000 ;
        RECT 72.790000 188.395000 72.990000 188.595000 ;
        RECT 72.790000 188.795000 72.990000 188.995000 ;
        RECT 72.790000 189.195000 72.990000 189.395000 ;
        RECT 72.790000 189.595000 72.990000 189.795000 ;
        RECT 72.790000 189.995000 72.990000 190.195000 ;
        RECT 72.790000 190.395000 72.990000 190.595000 ;
        RECT 72.790000 190.795000 72.990000 190.995000 ;
        RECT 72.790000 191.195000 72.990000 191.395000 ;
        RECT 72.790000 191.595000 72.990000 191.795000 ;
        RECT 72.790000 191.995000 72.990000 192.195000 ;
        RECT 72.790000 192.395000 72.990000 192.595000 ;
        RECT 72.790000 192.795000 72.990000 192.995000 ;
        RECT 72.790000 193.195000 72.990000 193.395000 ;
        RECT 72.790000 193.595000 72.990000 193.795000 ;
        RECT 72.790000 193.995000 72.990000 194.195000 ;
        RECT 72.790000 194.395000 72.990000 194.595000 ;
        RECT 72.790000 194.795000 72.990000 194.995000 ;
        RECT 72.790000 195.200000 72.990000 195.400000 ;
        RECT 72.790000 195.605000 72.990000 195.805000 ;
        RECT 72.790000 196.010000 72.990000 196.210000 ;
        RECT 72.790000 196.415000 72.990000 196.615000 ;
        RECT 72.790000 196.820000 72.990000 197.020000 ;
        RECT 72.790000 197.225000 72.990000 197.425000 ;
        RECT 72.790000 197.630000 72.990000 197.830000 ;
        RECT 72.790000 198.035000 72.990000 198.235000 ;
        RECT 72.790000 198.440000 72.990000 198.640000 ;
        RECT 72.790000 198.845000 72.990000 199.045000 ;
        RECT 72.790000 199.250000 72.990000 199.450000 ;
        RECT 72.790000 199.655000 72.990000 199.855000 ;
        RECT 73.190000  25.910000 73.390000  26.110000 ;
        RECT 73.190000  26.340000 73.390000  26.540000 ;
        RECT 73.190000  26.770000 73.390000  26.970000 ;
        RECT 73.190000  27.200000 73.390000  27.400000 ;
        RECT 73.190000  27.630000 73.390000  27.830000 ;
        RECT 73.190000  28.060000 73.390000  28.260000 ;
        RECT 73.190000  28.490000 73.390000  28.690000 ;
        RECT 73.190000  28.920000 73.390000  29.120000 ;
        RECT 73.190000  29.350000 73.390000  29.550000 ;
        RECT 73.190000  29.780000 73.390000  29.980000 ;
        RECT 73.190000  30.210000 73.390000  30.410000 ;
        RECT 73.190000 175.995000 73.390000 176.195000 ;
        RECT 73.190000 176.395000 73.390000 176.595000 ;
        RECT 73.190000 176.795000 73.390000 176.995000 ;
        RECT 73.190000 177.195000 73.390000 177.395000 ;
        RECT 73.190000 177.595000 73.390000 177.795000 ;
        RECT 73.190000 177.995000 73.390000 178.195000 ;
        RECT 73.190000 178.395000 73.390000 178.595000 ;
        RECT 73.190000 178.795000 73.390000 178.995000 ;
        RECT 73.190000 179.195000 73.390000 179.395000 ;
        RECT 73.190000 179.595000 73.390000 179.795000 ;
        RECT 73.190000 179.995000 73.390000 180.195000 ;
        RECT 73.190000 180.395000 73.390000 180.595000 ;
        RECT 73.190000 180.795000 73.390000 180.995000 ;
        RECT 73.190000 181.195000 73.390000 181.395000 ;
        RECT 73.190000 181.595000 73.390000 181.795000 ;
        RECT 73.190000 181.995000 73.390000 182.195000 ;
        RECT 73.190000 182.395000 73.390000 182.595000 ;
        RECT 73.190000 182.795000 73.390000 182.995000 ;
        RECT 73.190000 183.195000 73.390000 183.395000 ;
        RECT 73.190000 183.595000 73.390000 183.795000 ;
        RECT 73.190000 183.995000 73.390000 184.195000 ;
        RECT 73.190000 184.395000 73.390000 184.595000 ;
        RECT 73.190000 184.795000 73.390000 184.995000 ;
        RECT 73.190000 185.195000 73.390000 185.395000 ;
        RECT 73.190000 185.595000 73.390000 185.795000 ;
        RECT 73.190000 185.995000 73.390000 186.195000 ;
        RECT 73.190000 186.395000 73.390000 186.595000 ;
        RECT 73.190000 186.795000 73.390000 186.995000 ;
        RECT 73.190000 187.195000 73.390000 187.395000 ;
        RECT 73.190000 187.595000 73.390000 187.795000 ;
        RECT 73.190000 187.995000 73.390000 188.195000 ;
        RECT 73.190000 188.395000 73.390000 188.595000 ;
        RECT 73.190000 188.795000 73.390000 188.995000 ;
        RECT 73.190000 189.195000 73.390000 189.395000 ;
        RECT 73.190000 189.595000 73.390000 189.795000 ;
        RECT 73.190000 189.995000 73.390000 190.195000 ;
        RECT 73.190000 190.395000 73.390000 190.595000 ;
        RECT 73.190000 190.795000 73.390000 190.995000 ;
        RECT 73.190000 191.195000 73.390000 191.395000 ;
        RECT 73.190000 191.595000 73.390000 191.795000 ;
        RECT 73.190000 191.995000 73.390000 192.195000 ;
        RECT 73.190000 192.395000 73.390000 192.595000 ;
        RECT 73.190000 192.795000 73.390000 192.995000 ;
        RECT 73.190000 193.195000 73.390000 193.395000 ;
        RECT 73.190000 193.595000 73.390000 193.795000 ;
        RECT 73.190000 193.995000 73.390000 194.195000 ;
        RECT 73.190000 194.395000 73.390000 194.595000 ;
        RECT 73.190000 194.795000 73.390000 194.995000 ;
        RECT 73.190000 195.200000 73.390000 195.400000 ;
        RECT 73.190000 195.605000 73.390000 195.805000 ;
        RECT 73.190000 196.010000 73.390000 196.210000 ;
        RECT 73.190000 196.415000 73.390000 196.615000 ;
        RECT 73.190000 196.820000 73.390000 197.020000 ;
        RECT 73.190000 197.225000 73.390000 197.425000 ;
        RECT 73.190000 197.630000 73.390000 197.830000 ;
        RECT 73.190000 198.035000 73.390000 198.235000 ;
        RECT 73.190000 198.440000 73.390000 198.640000 ;
        RECT 73.190000 198.845000 73.390000 199.045000 ;
        RECT 73.190000 199.250000 73.390000 199.450000 ;
        RECT 73.190000 199.655000 73.390000 199.855000 ;
        RECT 73.590000 175.995000 73.790000 176.195000 ;
        RECT 73.590000 176.395000 73.790000 176.595000 ;
        RECT 73.590000 176.795000 73.790000 176.995000 ;
        RECT 73.590000 177.195000 73.790000 177.395000 ;
        RECT 73.590000 177.595000 73.790000 177.795000 ;
        RECT 73.590000 177.995000 73.790000 178.195000 ;
        RECT 73.590000 178.395000 73.790000 178.595000 ;
        RECT 73.590000 178.795000 73.790000 178.995000 ;
        RECT 73.590000 179.195000 73.790000 179.395000 ;
        RECT 73.590000 179.595000 73.790000 179.795000 ;
        RECT 73.590000 179.995000 73.790000 180.195000 ;
        RECT 73.590000 180.395000 73.790000 180.595000 ;
        RECT 73.590000 180.795000 73.790000 180.995000 ;
        RECT 73.590000 181.195000 73.790000 181.395000 ;
        RECT 73.590000 181.595000 73.790000 181.795000 ;
        RECT 73.590000 181.995000 73.790000 182.195000 ;
        RECT 73.590000 182.395000 73.790000 182.595000 ;
        RECT 73.590000 182.795000 73.790000 182.995000 ;
        RECT 73.590000 183.195000 73.790000 183.395000 ;
        RECT 73.590000 183.595000 73.790000 183.795000 ;
        RECT 73.590000 183.995000 73.790000 184.195000 ;
        RECT 73.590000 184.395000 73.790000 184.595000 ;
        RECT 73.590000 184.795000 73.790000 184.995000 ;
        RECT 73.590000 185.195000 73.790000 185.395000 ;
        RECT 73.590000 185.595000 73.790000 185.795000 ;
        RECT 73.590000 185.995000 73.790000 186.195000 ;
        RECT 73.590000 186.395000 73.790000 186.595000 ;
        RECT 73.590000 186.795000 73.790000 186.995000 ;
        RECT 73.590000 187.195000 73.790000 187.395000 ;
        RECT 73.590000 187.595000 73.790000 187.795000 ;
        RECT 73.590000 187.995000 73.790000 188.195000 ;
        RECT 73.590000 188.395000 73.790000 188.595000 ;
        RECT 73.590000 188.795000 73.790000 188.995000 ;
        RECT 73.590000 189.195000 73.790000 189.395000 ;
        RECT 73.590000 189.595000 73.790000 189.795000 ;
        RECT 73.590000 189.995000 73.790000 190.195000 ;
        RECT 73.590000 190.395000 73.790000 190.595000 ;
        RECT 73.590000 190.795000 73.790000 190.995000 ;
        RECT 73.590000 191.195000 73.790000 191.395000 ;
        RECT 73.590000 191.595000 73.790000 191.795000 ;
        RECT 73.590000 191.995000 73.790000 192.195000 ;
        RECT 73.590000 192.395000 73.790000 192.595000 ;
        RECT 73.590000 192.795000 73.790000 192.995000 ;
        RECT 73.590000 193.195000 73.790000 193.395000 ;
        RECT 73.590000 193.595000 73.790000 193.795000 ;
        RECT 73.590000 193.995000 73.790000 194.195000 ;
        RECT 73.590000 194.395000 73.790000 194.595000 ;
        RECT 73.590000 194.795000 73.790000 194.995000 ;
        RECT 73.590000 195.200000 73.790000 195.400000 ;
        RECT 73.590000 195.605000 73.790000 195.805000 ;
        RECT 73.590000 196.010000 73.790000 196.210000 ;
        RECT 73.590000 196.415000 73.790000 196.615000 ;
        RECT 73.590000 196.820000 73.790000 197.020000 ;
        RECT 73.590000 197.225000 73.790000 197.425000 ;
        RECT 73.590000 197.630000 73.790000 197.830000 ;
        RECT 73.590000 198.035000 73.790000 198.235000 ;
        RECT 73.590000 198.440000 73.790000 198.640000 ;
        RECT 73.590000 198.845000 73.790000 199.045000 ;
        RECT 73.590000 199.250000 73.790000 199.450000 ;
        RECT 73.590000 199.655000 73.790000 199.855000 ;
        RECT 73.595000  25.910000 73.795000  26.110000 ;
        RECT 73.595000  26.340000 73.795000  26.540000 ;
        RECT 73.595000  26.770000 73.795000  26.970000 ;
        RECT 73.595000  27.200000 73.795000  27.400000 ;
        RECT 73.595000  27.630000 73.795000  27.830000 ;
        RECT 73.595000  28.060000 73.795000  28.260000 ;
        RECT 73.595000  28.490000 73.795000  28.690000 ;
        RECT 73.595000  28.920000 73.795000  29.120000 ;
        RECT 73.595000  29.350000 73.795000  29.550000 ;
        RECT 73.595000  29.780000 73.795000  29.980000 ;
        RECT 73.595000  30.210000 73.795000  30.410000 ;
        RECT 73.990000 175.995000 74.190000 176.195000 ;
        RECT 73.990000 176.395000 74.190000 176.595000 ;
        RECT 73.990000 176.795000 74.190000 176.995000 ;
        RECT 73.990000 177.195000 74.190000 177.395000 ;
        RECT 73.990000 177.595000 74.190000 177.795000 ;
        RECT 73.990000 177.995000 74.190000 178.195000 ;
        RECT 73.990000 178.395000 74.190000 178.595000 ;
        RECT 73.990000 178.795000 74.190000 178.995000 ;
        RECT 73.990000 179.195000 74.190000 179.395000 ;
        RECT 73.990000 179.595000 74.190000 179.795000 ;
        RECT 73.990000 179.995000 74.190000 180.195000 ;
        RECT 73.990000 180.395000 74.190000 180.595000 ;
        RECT 73.990000 180.795000 74.190000 180.995000 ;
        RECT 73.990000 181.195000 74.190000 181.395000 ;
        RECT 73.990000 181.595000 74.190000 181.795000 ;
        RECT 73.990000 181.995000 74.190000 182.195000 ;
        RECT 73.990000 182.395000 74.190000 182.595000 ;
        RECT 73.990000 182.795000 74.190000 182.995000 ;
        RECT 73.990000 183.195000 74.190000 183.395000 ;
        RECT 73.990000 183.595000 74.190000 183.795000 ;
        RECT 73.990000 183.995000 74.190000 184.195000 ;
        RECT 73.990000 184.395000 74.190000 184.595000 ;
        RECT 73.990000 184.795000 74.190000 184.995000 ;
        RECT 73.990000 185.195000 74.190000 185.395000 ;
        RECT 73.990000 185.595000 74.190000 185.795000 ;
        RECT 73.990000 185.995000 74.190000 186.195000 ;
        RECT 73.990000 186.395000 74.190000 186.595000 ;
        RECT 73.990000 186.795000 74.190000 186.995000 ;
        RECT 73.990000 187.195000 74.190000 187.395000 ;
        RECT 73.990000 187.595000 74.190000 187.795000 ;
        RECT 73.990000 187.995000 74.190000 188.195000 ;
        RECT 73.990000 188.395000 74.190000 188.595000 ;
        RECT 73.990000 188.795000 74.190000 188.995000 ;
        RECT 73.990000 189.195000 74.190000 189.395000 ;
        RECT 73.990000 189.595000 74.190000 189.795000 ;
        RECT 73.990000 189.995000 74.190000 190.195000 ;
        RECT 73.990000 190.395000 74.190000 190.595000 ;
        RECT 73.990000 190.795000 74.190000 190.995000 ;
        RECT 73.990000 191.195000 74.190000 191.395000 ;
        RECT 73.990000 191.595000 74.190000 191.795000 ;
        RECT 73.990000 191.995000 74.190000 192.195000 ;
        RECT 73.990000 192.395000 74.190000 192.595000 ;
        RECT 73.990000 192.795000 74.190000 192.995000 ;
        RECT 73.990000 193.195000 74.190000 193.395000 ;
        RECT 73.990000 193.595000 74.190000 193.795000 ;
        RECT 73.990000 193.995000 74.190000 194.195000 ;
        RECT 73.990000 194.395000 74.190000 194.595000 ;
        RECT 73.990000 194.795000 74.190000 194.995000 ;
        RECT 73.990000 195.200000 74.190000 195.400000 ;
        RECT 73.990000 195.605000 74.190000 195.805000 ;
        RECT 73.990000 196.010000 74.190000 196.210000 ;
        RECT 73.990000 196.415000 74.190000 196.615000 ;
        RECT 73.990000 196.820000 74.190000 197.020000 ;
        RECT 73.990000 197.225000 74.190000 197.425000 ;
        RECT 73.990000 197.630000 74.190000 197.830000 ;
        RECT 73.990000 198.035000 74.190000 198.235000 ;
        RECT 73.990000 198.440000 74.190000 198.640000 ;
        RECT 73.990000 198.845000 74.190000 199.045000 ;
        RECT 73.990000 199.250000 74.190000 199.450000 ;
        RECT 73.990000 199.655000 74.190000 199.855000 ;
        RECT 74.000000  25.910000 74.200000  26.110000 ;
        RECT 74.000000  26.340000 74.200000  26.540000 ;
        RECT 74.000000  26.770000 74.200000  26.970000 ;
        RECT 74.000000  27.200000 74.200000  27.400000 ;
        RECT 74.000000  27.630000 74.200000  27.830000 ;
        RECT 74.000000  28.060000 74.200000  28.260000 ;
        RECT 74.000000  28.490000 74.200000  28.690000 ;
        RECT 74.000000  28.920000 74.200000  29.120000 ;
        RECT 74.000000  29.350000 74.200000  29.550000 ;
        RECT 74.000000  29.780000 74.200000  29.980000 ;
        RECT 74.000000  30.210000 74.200000  30.410000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.495000 58.240000 24.395000 62.680000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 58.240000 74.290000 62.680000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 24.370000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.585000 58.310000  0.785000 58.510000 ;
        RECT  0.585000 58.720000  0.785000 58.920000 ;
        RECT  0.585000 59.130000  0.785000 59.330000 ;
        RECT  0.585000 59.540000  0.785000 59.740000 ;
        RECT  0.585000 59.950000  0.785000 60.150000 ;
        RECT  0.585000 60.360000  0.785000 60.560000 ;
        RECT  0.585000 60.770000  0.785000 60.970000 ;
        RECT  0.585000 61.180000  0.785000 61.380000 ;
        RECT  0.585000 61.590000  0.785000 61.790000 ;
        RECT  0.585000 62.000000  0.785000 62.200000 ;
        RECT  0.585000 62.410000  0.785000 62.610000 ;
        RECT  0.995000 58.310000  1.195000 58.510000 ;
        RECT  0.995000 58.720000  1.195000 58.920000 ;
        RECT  0.995000 59.130000  1.195000 59.330000 ;
        RECT  0.995000 59.540000  1.195000 59.740000 ;
        RECT  0.995000 59.950000  1.195000 60.150000 ;
        RECT  0.995000 60.360000  1.195000 60.560000 ;
        RECT  0.995000 60.770000  1.195000 60.970000 ;
        RECT  0.995000 61.180000  1.195000 61.380000 ;
        RECT  0.995000 61.590000  1.195000 61.790000 ;
        RECT  0.995000 62.000000  1.195000 62.200000 ;
        RECT  0.995000 62.410000  1.195000 62.610000 ;
        RECT  1.405000 58.310000  1.605000 58.510000 ;
        RECT  1.405000 58.720000  1.605000 58.920000 ;
        RECT  1.405000 59.130000  1.605000 59.330000 ;
        RECT  1.405000 59.540000  1.605000 59.740000 ;
        RECT  1.405000 59.950000  1.605000 60.150000 ;
        RECT  1.405000 60.360000  1.605000 60.560000 ;
        RECT  1.405000 60.770000  1.605000 60.970000 ;
        RECT  1.405000 61.180000  1.605000 61.380000 ;
        RECT  1.405000 61.590000  1.605000 61.790000 ;
        RECT  1.405000 62.000000  1.605000 62.200000 ;
        RECT  1.405000 62.410000  1.605000 62.610000 ;
        RECT  1.815000 58.310000  2.015000 58.510000 ;
        RECT  1.815000 58.720000  2.015000 58.920000 ;
        RECT  1.815000 59.130000  2.015000 59.330000 ;
        RECT  1.815000 59.540000  2.015000 59.740000 ;
        RECT  1.815000 59.950000  2.015000 60.150000 ;
        RECT  1.815000 60.360000  2.015000 60.560000 ;
        RECT  1.815000 60.770000  2.015000 60.970000 ;
        RECT  1.815000 61.180000  2.015000 61.380000 ;
        RECT  1.815000 61.590000  2.015000 61.790000 ;
        RECT  1.815000 62.000000  2.015000 62.200000 ;
        RECT  1.815000 62.410000  2.015000 62.610000 ;
        RECT  2.225000 58.310000  2.425000 58.510000 ;
        RECT  2.225000 58.720000  2.425000 58.920000 ;
        RECT  2.225000 59.130000  2.425000 59.330000 ;
        RECT  2.225000 59.540000  2.425000 59.740000 ;
        RECT  2.225000 59.950000  2.425000 60.150000 ;
        RECT  2.225000 60.360000  2.425000 60.560000 ;
        RECT  2.225000 60.770000  2.425000 60.970000 ;
        RECT  2.225000 61.180000  2.425000 61.380000 ;
        RECT  2.225000 61.590000  2.425000 61.790000 ;
        RECT  2.225000 62.000000  2.425000 62.200000 ;
        RECT  2.225000 62.410000  2.425000 62.610000 ;
        RECT  2.635000 58.310000  2.835000 58.510000 ;
        RECT  2.635000 58.720000  2.835000 58.920000 ;
        RECT  2.635000 59.130000  2.835000 59.330000 ;
        RECT  2.635000 59.540000  2.835000 59.740000 ;
        RECT  2.635000 59.950000  2.835000 60.150000 ;
        RECT  2.635000 60.360000  2.835000 60.560000 ;
        RECT  2.635000 60.770000  2.835000 60.970000 ;
        RECT  2.635000 61.180000  2.835000 61.380000 ;
        RECT  2.635000 61.590000  2.835000 61.790000 ;
        RECT  2.635000 62.000000  2.835000 62.200000 ;
        RECT  2.635000 62.410000  2.835000 62.610000 ;
        RECT  3.045000 58.310000  3.245000 58.510000 ;
        RECT  3.045000 58.720000  3.245000 58.920000 ;
        RECT  3.045000 59.130000  3.245000 59.330000 ;
        RECT  3.045000 59.540000  3.245000 59.740000 ;
        RECT  3.045000 59.950000  3.245000 60.150000 ;
        RECT  3.045000 60.360000  3.245000 60.560000 ;
        RECT  3.045000 60.770000  3.245000 60.970000 ;
        RECT  3.045000 61.180000  3.245000 61.380000 ;
        RECT  3.045000 61.590000  3.245000 61.790000 ;
        RECT  3.045000 62.000000  3.245000 62.200000 ;
        RECT  3.045000 62.410000  3.245000 62.610000 ;
        RECT  3.450000 58.310000  3.650000 58.510000 ;
        RECT  3.450000 58.720000  3.650000 58.920000 ;
        RECT  3.450000 59.130000  3.650000 59.330000 ;
        RECT  3.450000 59.540000  3.650000 59.740000 ;
        RECT  3.450000 59.950000  3.650000 60.150000 ;
        RECT  3.450000 60.360000  3.650000 60.560000 ;
        RECT  3.450000 60.770000  3.650000 60.970000 ;
        RECT  3.450000 61.180000  3.650000 61.380000 ;
        RECT  3.450000 61.590000  3.650000 61.790000 ;
        RECT  3.450000 62.000000  3.650000 62.200000 ;
        RECT  3.450000 62.410000  3.650000 62.610000 ;
        RECT  3.855000 58.310000  4.055000 58.510000 ;
        RECT  3.855000 58.720000  4.055000 58.920000 ;
        RECT  3.855000 59.130000  4.055000 59.330000 ;
        RECT  3.855000 59.540000  4.055000 59.740000 ;
        RECT  3.855000 59.950000  4.055000 60.150000 ;
        RECT  3.855000 60.360000  4.055000 60.560000 ;
        RECT  3.855000 60.770000  4.055000 60.970000 ;
        RECT  3.855000 61.180000  4.055000 61.380000 ;
        RECT  3.855000 61.590000  4.055000 61.790000 ;
        RECT  3.855000 62.000000  4.055000 62.200000 ;
        RECT  3.855000 62.410000  4.055000 62.610000 ;
        RECT  4.260000 58.310000  4.460000 58.510000 ;
        RECT  4.260000 58.720000  4.460000 58.920000 ;
        RECT  4.260000 59.130000  4.460000 59.330000 ;
        RECT  4.260000 59.540000  4.460000 59.740000 ;
        RECT  4.260000 59.950000  4.460000 60.150000 ;
        RECT  4.260000 60.360000  4.460000 60.560000 ;
        RECT  4.260000 60.770000  4.460000 60.970000 ;
        RECT  4.260000 61.180000  4.460000 61.380000 ;
        RECT  4.260000 61.590000  4.460000 61.790000 ;
        RECT  4.260000 62.000000  4.460000 62.200000 ;
        RECT  4.260000 62.410000  4.460000 62.610000 ;
        RECT  4.665000 58.310000  4.865000 58.510000 ;
        RECT  4.665000 58.720000  4.865000 58.920000 ;
        RECT  4.665000 59.130000  4.865000 59.330000 ;
        RECT  4.665000 59.540000  4.865000 59.740000 ;
        RECT  4.665000 59.950000  4.865000 60.150000 ;
        RECT  4.665000 60.360000  4.865000 60.560000 ;
        RECT  4.665000 60.770000  4.865000 60.970000 ;
        RECT  4.665000 61.180000  4.865000 61.380000 ;
        RECT  4.665000 61.590000  4.865000 61.790000 ;
        RECT  4.665000 62.000000  4.865000 62.200000 ;
        RECT  4.665000 62.410000  4.865000 62.610000 ;
        RECT  5.070000 58.310000  5.270000 58.510000 ;
        RECT  5.070000 58.720000  5.270000 58.920000 ;
        RECT  5.070000 59.130000  5.270000 59.330000 ;
        RECT  5.070000 59.540000  5.270000 59.740000 ;
        RECT  5.070000 59.950000  5.270000 60.150000 ;
        RECT  5.070000 60.360000  5.270000 60.560000 ;
        RECT  5.070000 60.770000  5.270000 60.970000 ;
        RECT  5.070000 61.180000  5.270000 61.380000 ;
        RECT  5.070000 61.590000  5.270000 61.790000 ;
        RECT  5.070000 62.000000  5.270000 62.200000 ;
        RECT  5.070000 62.410000  5.270000 62.610000 ;
        RECT  5.475000 58.310000  5.675000 58.510000 ;
        RECT  5.475000 58.720000  5.675000 58.920000 ;
        RECT  5.475000 59.130000  5.675000 59.330000 ;
        RECT  5.475000 59.540000  5.675000 59.740000 ;
        RECT  5.475000 59.950000  5.675000 60.150000 ;
        RECT  5.475000 60.360000  5.675000 60.560000 ;
        RECT  5.475000 60.770000  5.675000 60.970000 ;
        RECT  5.475000 61.180000  5.675000 61.380000 ;
        RECT  5.475000 61.590000  5.675000 61.790000 ;
        RECT  5.475000 62.000000  5.675000 62.200000 ;
        RECT  5.475000 62.410000  5.675000 62.610000 ;
        RECT  5.880000 58.310000  6.080000 58.510000 ;
        RECT  5.880000 58.720000  6.080000 58.920000 ;
        RECT  5.880000 59.130000  6.080000 59.330000 ;
        RECT  5.880000 59.540000  6.080000 59.740000 ;
        RECT  5.880000 59.950000  6.080000 60.150000 ;
        RECT  5.880000 60.360000  6.080000 60.560000 ;
        RECT  5.880000 60.770000  6.080000 60.970000 ;
        RECT  5.880000 61.180000  6.080000 61.380000 ;
        RECT  5.880000 61.590000  6.080000 61.790000 ;
        RECT  5.880000 62.000000  6.080000 62.200000 ;
        RECT  5.880000 62.410000  6.080000 62.610000 ;
        RECT  6.285000 58.310000  6.485000 58.510000 ;
        RECT  6.285000 58.720000  6.485000 58.920000 ;
        RECT  6.285000 59.130000  6.485000 59.330000 ;
        RECT  6.285000 59.540000  6.485000 59.740000 ;
        RECT  6.285000 59.950000  6.485000 60.150000 ;
        RECT  6.285000 60.360000  6.485000 60.560000 ;
        RECT  6.285000 60.770000  6.485000 60.970000 ;
        RECT  6.285000 61.180000  6.485000 61.380000 ;
        RECT  6.285000 61.590000  6.485000 61.790000 ;
        RECT  6.285000 62.000000  6.485000 62.200000 ;
        RECT  6.285000 62.410000  6.485000 62.610000 ;
        RECT  6.690000 58.310000  6.890000 58.510000 ;
        RECT  6.690000 58.720000  6.890000 58.920000 ;
        RECT  6.690000 59.130000  6.890000 59.330000 ;
        RECT  6.690000 59.540000  6.890000 59.740000 ;
        RECT  6.690000 59.950000  6.890000 60.150000 ;
        RECT  6.690000 60.360000  6.890000 60.560000 ;
        RECT  6.690000 60.770000  6.890000 60.970000 ;
        RECT  6.690000 61.180000  6.890000 61.380000 ;
        RECT  6.690000 61.590000  6.890000 61.790000 ;
        RECT  6.690000 62.000000  6.890000 62.200000 ;
        RECT  6.690000 62.410000  6.890000 62.610000 ;
        RECT  7.095000 58.310000  7.295000 58.510000 ;
        RECT  7.095000 58.720000  7.295000 58.920000 ;
        RECT  7.095000 59.130000  7.295000 59.330000 ;
        RECT  7.095000 59.540000  7.295000 59.740000 ;
        RECT  7.095000 59.950000  7.295000 60.150000 ;
        RECT  7.095000 60.360000  7.295000 60.560000 ;
        RECT  7.095000 60.770000  7.295000 60.970000 ;
        RECT  7.095000 61.180000  7.295000 61.380000 ;
        RECT  7.095000 61.590000  7.295000 61.790000 ;
        RECT  7.095000 62.000000  7.295000 62.200000 ;
        RECT  7.095000 62.410000  7.295000 62.610000 ;
        RECT  7.500000 58.310000  7.700000 58.510000 ;
        RECT  7.500000 58.720000  7.700000 58.920000 ;
        RECT  7.500000 59.130000  7.700000 59.330000 ;
        RECT  7.500000 59.540000  7.700000 59.740000 ;
        RECT  7.500000 59.950000  7.700000 60.150000 ;
        RECT  7.500000 60.360000  7.700000 60.560000 ;
        RECT  7.500000 60.770000  7.700000 60.970000 ;
        RECT  7.500000 61.180000  7.700000 61.380000 ;
        RECT  7.500000 61.590000  7.700000 61.790000 ;
        RECT  7.500000 62.000000  7.700000 62.200000 ;
        RECT  7.500000 62.410000  7.700000 62.610000 ;
        RECT  7.905000 58.310000  8.105000 58.510000 ;
        RECT  7.905000 58.720000  8.105000 58.920000 ;
        RECT  7.905000 59.130000  8.105000 59.330000 ;
        RECT  7.905000 59.540000  8.105000 59.740000 ;
        RECT  7.905000 59.950000  8.105000 60.150000 ;
        RECT  7.905000 60.360000  8.105000 60.560000 ;
        RECT  7.905000 60.770000  8.105000 60.970000 ;
        RECT  7.905000 61.180000  8.105000 61.380000 ;
        RECT  7.905000 61.590000  8.105000 61.790000 ;
        RECT  7.905000 62.000000  8.105000 62.200000 ;
        RECT  7.905000 62.410000  8.105000 62.610000 ;
        RECT  8.310000 58.310000  8.510000 58.510000 ;
        RECT  8.310000 58.720000  8.510000 58.920000 ;
        RECT  8.310000 59.130000  8.510000 59.330000 ;
        RECT  8.310000 59.540000  8.510000 59.740000 ;
        RECT  8.310000 59.950000  8.510000 60.150000 ;
        RECT  8.310000 60.360000  8.510000 60.560000 ;
        RECT  8.310000 60.770000  8.510000 60.970000 ;
        RECT  8.310000 61.180000  8.510000 61.380000 ;
        RECT  8.310000 61.590000  8.510000 61.790000 ;
        RECT  8.310000 62.000000  8.510000 62.200000 ;
        RECT  8.310000 62.410000  8.510000 62.610000 ;
        RECT  8.715000 58.310000  8.915000 58.510000 ;
        RECT  8.715000 58.720000  8.915000 58.920000 ;
        RECT  8.715000 59.130000  8.915000 59.330000 ;
        RECT  8.715000 59.540000  8.915000 59.740000 ;
        RECT  8.715000 59.950000  8.915000 60.150000 ;
        RECT  8.715000 60.360000  8.915000 60.560000 ;
        RECT  8.715000 60.770000  8.915000 60.970000 ;
        RECT  8.715000 61.180000  8.915000 61.380000 ;
        RECT  8.715000 61.590000  8.915000 61.790000 ;
        RECT  8.715000 62.000000  8.915000 62.200000 ;
        RECT  8.715000 62.410000  8.915000 62.610000 ;
        RECT  9.120000 58.310000  9.320000 58.510000 ;
        RECT  9.120000 58.720000  9.320000 58.920000 ;
        RECT  9.120000 59.130000  9.320000 59.330000 ;
        RECT  9.120000 59.540000  9.320000 59.740000 ;
        RECT  9.120000 59.950000  9.320000 60.150000 ;
        RECT  9.120000 60.360000  9.320000 60.560000 ;
        RECT  9.120000 60.770000  9.320000 60.970000 ;
        RECT  9.120000 61.180000  9.320000 61.380000 ;
        RECT  9.120000 61.590000  9.320000 61.790000 ;
        RECT  9.120000 62.000000  9.320000 62.200000 ;
        RECT  9.120000 62.410000  9.320000 62.610000 ;
        RECT  9.525000 58.310000  9.725000 58.510000 ;
        RECT  9.525000 58.720000  9.725000 58.920000 ;
        RECT  9.525000 59.130000  9.725000 59.330000 ;
        RECT  9.525000 59.540000  9.725000 59.740000 ;
        RECT  9.525000 59.950000  9.725000 60.150000 ;
        RECT  9.525000 60.360000  9.725000 60.560000 ;
        RECT  9.525000 60.770000  9.725000 60.970000 ;
        RECT  9.525000 61.180000  9.725000 61.380000 ;
        RECT  9.525000 61.590000  9.725000 61.790000 ;
        RECT  9.525000 62.000000  9.725000 62.200000 ;
        RECT  9.525000 62.410000  9.725000 62.610000 ;
        RECT  9.930000 58.310000 10.130000 58.510000 ;
        RECT  9.930000 58.720000 10.130000 58.920000 ;
        RECT  9.930000 59.130000 10.130000 59.330000 ;
        RECT  9.930000 59.540000 10.130000 59.740000 ;
        RECT  9.930000 59.950000 10.130000 60.150000 ;
        RECT  9.930000 60.360000 10.130000 60.560000 ;
        RECT  9.930000 60.770000 10.130000 60.970000 ;
        RECT  9.930000 61.180000 10.130000 61.380000 ;
        RECT  9.930000 61.590000 10.130000 61.790000 ;
        RECT  9.930000 62.000000 10.130000 62.200000 ;
        RECT  9.930000 62.410000 10.130000 62.610000 ;
        RECT 10.335000 58.310000 10.535000 58.510000 ;
        RECT 10.335000 58.720000 10.535000 58.920000 ;
        RECT 10.335000 59.130000 10.535000 59.330000 ;
        RECT 10.335000 59.540000 10.535000 59.740000 ;
        RECT 10.335000 59.950000 10.535000 60.150000 ;
        RECT 10.335000 60.360000 10.535000 60.560000 ;
        RECT 10.335000 60.770000 10.535000 60.970000 ;
        RECT 10.335000 61.180000 10.535000 61.380000 ;
        RECT 10.335000 61.590000 10.535000 61.790000 ;
        RECT 10.335000 62.000000 10.535000 62.200000 ;
        RECT 10.335000 62.410000 10.535000 62.610000 ;
        RECT 10.740000 58.310000 10.940000 58.510000 ;
        RECT 10.740000 58.720000 10.940000 58.920000 ;
        RECT 10.740000 59.130000 10.940000 59.330000 ;
        RECT 10.740000 59.540000 10.940000 59.740000 ;
        RECT 10.740000 59.950000 10.940000 60.150000 ;
        RECT 10.740000 60.360000 10.940000 60.560000 ;
        RECT 10.740000 60.770000 10.940000 60.970000 ;
        RECT 10.740000 61.180000 10.940000 61.380000 ;
        RECT 10.740000 61.590000 10.940000 61.790000 ;
        RECT 10.740000 62.000000 10.940000 62.200000 ;
        RECT 10.740000 62.410000 10.940000 62.610000 ;
        RECT 11.145000 58.310000 11.345000 58.510000 ;
        RECT 11.145000 58.720000 11.345000 58.920000 ;
        RECT 11.145000 59.130000 11.345000 59.330000 ;
        RECT 11.145000 59.540000 11.345000 59.740000 ;
        RECT 11.145000 59.950000 11.345000 60.150000 ;
        RECT 11.145000 60.360000 11.345000 60.560000 ;
        RECT 11.145000 60.770000 11.345000 60.970000 ;
        RECT 11.145000 61.180000 11.345000 61.380000 ;
        RECT 11.145000 61.590000 11.345000 61.790000 ;
        RECT 11.145000 62.000000 11.345000 62.200000 ;
        RECT 11.145000 62.410000 11.345000 62.610000 ;
        RECT 11.550000 58.310000 11.750000 58.510000 ;
        RECT 11.550000 58.720000 11.750000 58.920000 ;
        RECT 11.550000 59.130000 11.750000 59.330000 ;
        RECT 11.550000 59.540000 11.750000 59.740000 ;
        RECT 11.550000 59.950000 11.750000 60.150000 ;
        RECT 11.550000 60.360000 11.750000 60.560000 ;
        RECT 11.550000 60.770000 11.750000 60.970000 ;
        RECT 11.550000 61.180000 11.750000 61.380000 ;
        RECT 11.550000 61.590000 11.750000 61.790000 ;
        RECT 11.550000 62.000000 11.750000 62.200000 ;
        RECT 11.550000 62.410000 11.750000 62.610000 ;
        RECT 11.955000 58.310000 12.155000 58.510000 ;
        RECT 11.955000 58.720000 12.155000 58.920000 ;
        RECT 11.955000 59.130000 12.155000 59.330000 ;
        RECT 11.955000 59.540000 12.155000 59.740000 ;
        RECT 11.955000 59.950000 12.155000 60.150000 ;
        RECT 11.955000 60.360000 12.155000 60.560000 ;
        RECT 11.955000 60.770000 12.155000 60.970000 ;
        RECT 11.955000 61.180000 12.155000 61.380000 ;
        RECT 11.955000 61.590000 12.155000 61.790000 ;
        RECT 11.955000 62.000000 12.155000 62.200000 ;
        RECT 11.955000 62.410000 12.155000 62.610000 ;
        RECT 12.360000 58.310000 12.560000 58.510000 ;
        RECT 12.360000 58.720000 12.560000 58.920000 ;
        RECT 12.360000 59.130000 12.560000 59.330000 ;
        RECT 12.360000 59.540000 12.560000 59.740000 ;
        RECT 12.360000 59.950000 12.560000 60.150000 ;
        RECT 12.360000 60.360000 12.560000 60.560000 ;
        RECT 12.360000 60.770000 12.560000 60.970000 ;
        RECT 12.360000 61.180000 12.560000 61.380000 ;
        RECT 12.360000 61.590000 12.560000 61.790000 ;
        RECT 12.360000 62.000000 12.560000 62.200000 ;
        RECT 12.360000 62.410000 12.560000 62.610000 ;
        RECT 12.765000 58.310000 12.965000 58.510000 ;
        RECT 12.765000 58.720000 12.965000 58.920000 ;
        RECT 12.765000 59.130000 12.965000 59.330000 ;
        RECT 12.765000 59.540000 12.965000 59.740000 ;
        RECT 12.765000 59.950000 12.965000 60.150000 ;
        RECT 12.765000 60.360000 12.965000 60.560000 ;
        RECT 12.765000 60.770000 12.965000 60.970000 ;
        RECT 12.765000 61.180000 12.965000 61.380000 ;
        RECT 12.765000 61.590000 12.965000 61.790000 ;
        RECT 12.765000 62.000000 12.965000 62.200000 ;
        RECT 12.765000 62.410000 12.965000 62.610000 ;
        RECT 13.170000 58.310000 13.370000 58.510000 ;
        RECT 13.170000 58.720000 13.370000 58.920000 ;
        RECT 13.170000 59.130000 13.370000 59.330000 ;
        RECT 13.170000 59.540000 13.370000 59.740000 ;
        RECT 13.170000 59.950000 13.370000 60.150000 ;
        RECT 13.170000 60.360000 13.370000 60.560000 ;
        RECT 13.170000 60.770000 13.370000 60.970000 ;
        RECT 13.170000 61.180000 13.370000 61.380000 ;
        RECT 13.170000 61.590000 13.370000 61.790000 ;
        RECT 13.170000 62.000000 13.370000 62.200000 ;
        RECT 13.170000 62.410000 13.370000 62.610000 ;
        RECT 13.575000 58.310000 13.775000 58.510000 ;
        RECT 13.575000 58.720000 13.775000 58.920000 ;
        RECT 13.575000 59.130000 13.775000 59.330000 ;
        RECT 13.575000 59.540000 13.775000 59.740000 ;
        RECT 13.575000 59.950000 13.775000 60.150000 ;
        RECT 13.575000 60.360000 13.775000 60.560000 ;
        RECT 13.575000 60.770000 13.775000 60.970000 ;
        RECT 13.575000 61.180000 13.775000 61.380000 ;
        RECT 13.575000 61.590000 13.775000 61.790000 ;
        RECT 13.575000 62.000000 13.775000 62.200000 ;
        RECT 13.575000 62.410000 13.775000 62.610000 ;
        RECT 13.980000 58.310000 14.180000 58.510000 ;
        RECT 13.980000 58.720000 14.180000 58.920000 ;
        RECT 13.980000 59.130000 14.180000 59.330000 ;
        RECT 13.980000 59.540000 14.180000 59.740000 ;
        RECT 13.980000 59.950000 14.180000 60.150000 ;
        RECT 13.980000 60.360000 14.180000 60.560000 ;
        RECT 13.980000 60.770000 14.180000 60.970000 ;
        RECT 13.980000 61.180000 14.180000 61.380000 ;
        RECT 13.980000 61.590000 14.180000 61.790000 ;
        RECT 13.980000 62.000000 14.180000 62.200000 ;
        RECT 13.980000 62.410000 14.180000 62.610000 ;
        RECT 14.385000 58.310000 14.585000 58.510000 ;
        RECT 14.385000 58.720000 14.585000 58.920000 ;
        RECT 14.385000 59.130000 14.585000 59.330000 ;
        RECT 14.385000 59.540000 14.585000 59.740000 ;
        RECT 14.385000 59.950000 14.585000 60.150000 ;
        RECT 14.385000 60.360000 14.585000 60.560000 ;
        RECT 14.385000 60.770000 14.585000 60.970000 ;
        RECT 14.385000 61.180000 14.585000 61.380000 ;
        RECT 14.385000 61.590000 14.585000 61.790000 ;
        RECT 14.385000 62.000000 14.585000 62.200000 ;
        RECT 14.385000 62.410000 14.585000 62.610000 ;
        RECT 14.790000 58.310000 14.990000 58.510000 ;
        RECT 14.790000 58.720000 14.990000 58.920000 ;
        RECT 14.790000 59.130000 14.990000 59.330000 ;
        RECT 14.790000 59.540000 14.990000 59.740000 ;
        RECT 14.790000 59.950000 14.990000 60.150000 ;
        RECT 14.790000 60.360000 14.990000 60.560000 ;
        RECT 14.790000 60.770000 14.990000 60.970000 ;
        RECT 14.790000 61.180000 14.990000 61.380000 ;
        RECT 14.790000 61.590000 14.990000 61.790000 ;
        RECT 14.790000 62.000000 14.990000 62.200000 ;
        RECT 14.790000 62.410000 14.990000 62.610000 ;
        RECT 15.195000 58.310000 15.395000 58.510000 ;
        RECT 15.195000 58.720000 15.395000 58.920000 ;
        RECT 15.195000 59.130000 15.395000 59.330000 ;
        RECT 15.195000 59.540000 15.395000 59.740000 ;
        RECT 15.195000 59.950000 15.395000 60.150000 ;
        RECT 15.195000 60.360000 15.395000 60.560000 ;
        RECT 15.195000 60.770000 15.395000 60.970000 ;
        RECT 15.195000 61.180000 15.395000 61.380000 ;
        RECT 15.195000 61.590000 15.395000 61.790000 ;
        RECT 15.195000 62.000000 15.395000 62.200000 ;
        RECT 15.195000 62.410000 15.395000 62.610000 ;
        RECT 15.600000 58.310000 15.800000 58.510000 ;
        RECT 15.600000 58.720000 15.800000 58.920000 ;
        RECT 15.600000 59.130000 15.800000 59.330000 ;
        RECT 15.600000 59.540000 15.800000 59.740000 ;
        RECT 15.600000 59.950000 15.800000 60.150000 ;
        RECT 15.600000 60.360000 15.800000 60.560000 ;
        RECT 15.600000 60.770000 15.800000 60.970000 ;
        RECT 15.600000 61.180000 15.800000 61.380000 ;
        RECT 15.600000 61.590000 15.800000 61.790000 ;
        RECT 15.600000 62.000000 15.800000 62.200000 ;
        RECT 15.600000 62.410000 15.800000 62.610000 ;
        RECT 16.005000 58.310000 16.205000 58.510000 ;
        RECT 16.005000 58.720000 16.205000 58.920000 ;
        RECT 16.005000 59.130000 16.205000 59.330000 ;
        RECT 16.005000 59.540000 16.205000 59.740000 ;
        RECT 16.005000 59.950000 16.205000 60.150000 ;
        RECT 16.005000 60.360000 16.205000 60.560000 ;
        RECT 16.005000 60.770000 16.205000 60.970000 ;
        RECT 16.005000 61.180000 16.205000 61.380000 ;
        RECT 16.005000 61.590000 16.205000 61.790000 ;
        RECT 16.005000 62.000000 16.205000 62.200000 ;
        RECT 16.005000 62.410000 16.205000 62.610000 ;
        RECT 16.410000 58.310000 16.610000 58.510000 ;
        RECT 16.410000 58.720000 16.610000 58.920000 ;
        RECT 16.410000 59.130000 16.610000 59.330000 ;
        RECT 16.410000 59.540000 16.610000 59.740000 ;
        RECT 16.410000 59.950000 16.610000 60.150000 ;
        RECT 16.410000 60.360000 16.610000 60.560000 ;
        RECT 16.410000 60.770000 16.610000 60.970000 ;
        RECT 16.410000 61.180000 16.610000 61.380000 ;
        RECT 16.410000 61.590000 16.610000 61.790000 ;
        RECT 16.410000 62.000000 16.610000 62.200000 ;
        RECT 16.410000 62.410000 16.610000 62.610000 ;
        RECT 16.815000 58.310000 17.015000 58.510000 ;
        RECT 16.815000 58.720000 17.015000 58.920000 ;
        RECT 16.815000 59.130000 17.015000 59.330000 ;
        RECT 16.815000 59.540000 17.015000 59.740000 ;
        RECT 16.815000 59.950000 17.015000 60.150000 ;
        RECT 16.815000 60.360000 17.015000 60.560000 ;
        RECT 16.815000 60.770000 17.015000 60.970000 ;
        RECT 16.815000 61.180000 17.015000 61.380000 ;
        RECT 16.815000 61.590000 17.015000 61.790000 ;
        RECT 16.815000 62.000000 17.015000 62.200000 ;
        RECT 16.815000 62.410000 17.015000 62.610000 ;
        RECT 17.220000 58.310000 17.420000 58.510000 ;
        RECT 17.220000 58.720000 17.420000 58.920000 ;
        RECT 17.220000 59.130000 17.420000 59.330000 ;
        RECT 17.220000 59.540000 17.420000 59.740000 ;
        RECT 17.220000 59.950000 17.420000 60.150000 ;
        RECT 17.220000 60.360000 17.420000 60.560000 ;
        RECT 17.220000 60.770000 17.420000 60.970000 ;
        RECT 17.220000 61.180000 17.420000 61.380000 ;
        RECT 17.220000 61.590000 17.420000 61.790000 ;
        RECT 17.220000 62.000000 17.420000 62.200000 ;
        RECT 17.220000 62.410000 17.420000 62.610000 ;
        RECT 17.625000 58.310000 17.825000 58.510000 ;
        RECT 17.625000 58.720000 17.825000 58.920000 ;
        RECT 17.625000 59.130000 17.825000 59.330000 ;
        RECT 17.625000 59.540000 17.825000 59.740000 ;
        RECT 17.625000 59.950000 17.825000 60.150000 ;
        RECT 17.625000 60.360000 17.825000 60.560000 ;
        RECT 17.625000 60.770000 17.825000 60.970000 ;
        RECT 17.625000 61.180000 17.825000 61.380000 ;
        RECT 17.625000 61.590000 17.825000 61.790000 ;
        RECT 17.625000 62.000000 17.825000 62.200000 ;
        RECT 17.625000 62.410000 17.825000 62.610000 ;
        RECT 18.030000 58.310000 18.230000 58.510000 ;
        RECT 18.030000 58.720000 18.230000 58.920000 ;
        RECT 18.030000 59.130000 18.230000 59.330000 ;
        RECT 18.030000 59.540000 18.230000 59.740000 ;
        RECT 18.030000 59.950000 18.230000 60.150000 ;
        RECT 18.030000 60.360000 18.230000 60.560000 ;
        RECT 18.030000 60.770000 18.230000 60.970000 ;
        RECT 18.030000 61.180000 18.230000 61.380000 ;
        RECT 18.030000 61.590000 18.230000 61.790000 ;
        RECT 18.030000 62.000000 18.230000 62.200000 ;
        RECT 18.030000 62.410000 18.230000 62.610000 ;
        RECT 18.435000 58.310000 18.635000 58.510000 ;
        RECT 18.435000 58.720000 18.635000 58.920000 ;
        RECT 18.435000 59.130000 18.635000 59.330000 ;
        RECT 18.435000 59.540000 18.635000 59.740000 ;
        RECT 18.435000 59.950000 18.635000 60.150000 ;
        RECT 18.435000 60.360000 18.635000 60.560000 ;
        RECT 18.435000 60.770000 18.635000 60.970000 ;
        RECT 18.435000 61.180000 18.635000 61.380000 ;
        RECT 18.435000 61.590000 18.635000 61.790000 ;
        RECT 18.435000 62.000000 18.635000 62.200000 ;
        RECT 18.435000 62.410000 18.635000 62.610000 ;
        RECT 18.840000 58.310000 19.040000 58.510000 ;
        RECT 18.840000 58.720000 19.040000 58.920000 ;
        RECT 18.840000 59.130000 19.040000 59.330000 ;
        RECT 18.840000 59.540000 19.040000 59.740000 ;
        RECT 18.840000 59.950000 19.040000 60.150000 ;
        RECT 18.840000 60.360000 19.040000 60.560000 ;
        RECT 18.840000 60.770000 19.040000 60.970000 ;
        RECT 18.840000 61.180000 19.040000 61.380000 ;
        RECT 18.840000 61.590000 19.040000 61.790000 ;
        RECT 18.840000 62.000000 19.040000 62.200000 ;
        RECT 18.840000 62.410000 19.040000 62.610000 ;
        RECT 19.245000 58.310000 19.445000 58.510000 ;
        RECT 19.245000 58.720000 19.445000 58.920000 ;
        RECT 19.245000 59.130000 19.445000 59.330000 ;
        RECT 19.245000 59.540000 19.445000 59.740000 ;
        RECT 19.245000 59.950000 19.445000 60.150000 ;
        RECT 19.245000 60.360000 19.445000 60.560000 ;
        RECT 19.245000 60.770000 19.445000 60.970000 ;
        RECT 19.245000 61.180000 19.445000 61.380000 ;
        RECT 19.245000 61.590000 19.445000 61.790000 ;
        RECT 19.245000 62.000000 19.445000 62.200000 ;
        RECT 19.245000 62.410000 19.445000 62.610000 ;
        RECT 19.650000 58.310000 19.850000 58.510000 ;
        RECT 19.650000 58.720000 19.850000 58.920000 ;
        RECT 19.650000 59.130000 19.850000 59.330000 ;
        RECT 19.650000 59.540000 19.850000 59.740000 ;
        RECT 19.650000 59.950000 19.850000 60.150000 ;
        RECT 19.650000 60.360000 19.850000 60.560000 ;
        RECT 19.650000 60.770000 19.850000 60.970000 ;
        RECT 19.650000 61.180000 19.850000 61.380000 ;
        RECT 19.650000 61.590000 19.850000 61.790000 ;
        RECT 19.650000 62.000000 19.850000 62.200000 ;
        RECT 19.650000 62.410000 19.850000 62.610000 ;
        RECT 20.055000 58.310000 20.255000 58.510000 ;
        RECT 20.055000 58.720000 20.255000 58.920000 ;
        RECT 20.055000 59.130000 20.255000 59.330000 ;
        RECT 20.055000 59.540000 20.255000 59.740000 ;
        RECT 20.055000 59.950000 20.255000 60.150000 ;
        RECT 20.055000 60.360000 20.255000 60.560000 ;
        RECT 20.055000 60.770000 20.255000 60.970000 ;
        RECT 20.055000 61.180000 20.255000 61.380000 ;
        RECT 20.055000 61.590000 20.255000 61.790000 ;
        RECT 20.055000 62.000000 20.255000 62.200000 ;
        RECT 20.055000 62.410000 20.255000 62.610000 ;
        RECT 20.460000 58.310000 20.660000 58.510000 ;
        RECT 20.460000 58.720000 20.660000 58.920000 ;
        RECT 20.460000 59.130000 20.660000 59.330000 ;
        RECT 20.460000 59.540000 20.660000 59.740000 ;
        RECT 20.460000 59.950000 20.660000 60.150000 ;
        RECT 20.460000 60.360000 20.660000 60.560000 ;
        RECT 20.460000 60.770000 20.660000 60.970000 ;
        RECT 20.460000 61.180000 20.660000 61.380000 ;
        RECT 20.460000 61.590000 20.660000 61.790000 ;
        RECT 20.460000 62.000000 20.660000 62.200000 ;
        RECT 20.460000 62.410000 20.660000 62.610000 ;
        RECT 20.865000 58.310000 21.065000 58.510000 ;
        RECT 20.865000 58.720000 21.065000 58.920000 ;
        RECT 20.865000 59.130000 21.065000 59.330000 ;
        RECT 20.865000 59.540000 21.065000 59.740000 ;
        RECT 20.865000 59.950000 21.065000 60.150000 ;
        RECT 20.865000 60.360000 21.065000 60.560000 ;
        RECT 20.865000 60.770000 21.065000 60.970000 ;
        RECT 20.865000 61.180000 21.065000 61.380000 ;
        RECT 20.865000 61.590000 21.065000 61.790000 ;
        RECT 20.865000 62.000000 21.065000 62.200000 ;
        RECT 20.865000 62.410000 21.065000 62.610000 ;
        RECT 21.270000 58.310000 21.470000 58.510000 ;
        RECT 21.270000 58.720000 21.470000 58.920000 ;
        RECT 21.270000 59.130000 21.470000 59.330000 ;
        RECT 21.270000 59.540000 21.470000 59.740000 ;
        RECT 21.270000 59.950000 21.470000 60.150000 ;
        RECT 21.270000 60.360000 21.470000 60.560000 ;
        RECT 21.270000 60.770000 21.470000 60.970000 ;
        RECT 21.270000 61.180000 21.470000 61.380000 ;
        RECT 21.270000 61.590000 21.470000 61.790000 ;
        RECT 21.270000 62.000000 21.470000 62.200000 ;
        RECT 21.270000 62.410000 21.470000 62.610000 ;
        RECT 21.675000 58.310000 21.875000 58.510000 ;
        RECT 21.675000 58.720000 21.875000 58.920000 ;
        RECT 21.675000 59.130000 21.875000 59.330000 ;
        RECT 21.675000 59.540000 21.875000 59.740000 ;
        RECT 21.675000 59.950000 21.875000 60.150000 ;
        RECT 21.675000 60.360000 21.875000 60.560000 ;
        RECT 21.675000 60.770000 21.875000 60.970000 ;
        RECT 21.675000 61.180000 21.875000 61.380000 ;
        RECT 21.675000 61.590000 21.875000 61.790000 ;
        RECT 21.675000 62.000000 21.875000 62.200000 ;
        RECT 21.675000 62.410000 21.875000 62.610000 ;
        RECT 22.080000 58.310000 22.280000 58.510000 ;
        RECT 22.080000 58.720000 22.280000 58.920000 ;
        RECT 22.080000 59.130000 22.280000 59.330000 ;
        RECT 22.080000 59.540000 22.280000 59.740000 ;
        RECT 22.080000 59.950000 22.280000 60.150000 ;
        RECT 22.080000 60.360000 22.280000 60.560000 ;
        RECT 22.080000 60.770000 22.280000 60.970000 ;
        RECT 22.080000 61.180000 22.280000 61.380000 ;
        RECT 22.080000 61.590000 22.280000 61.790000 ;
        RECT 22.080000 62.000000 22.280000 62.200000 ;
        RECT 22.080000 62.410000 22.280000 62.610000 ;
        RECT 22.485000 58.310000 22.685000 58.510000 ;
        RECT 22.485000 58.720000 22.685000 58.920000 ;
        RECT 22.485000 59.130000 22.685000 59.330000 ;
        RECT 22.485000 59.540000 22.685000 59.740000 ;
        RECT 22.485000 59.950000 22.685000 60.150000 ;
        RECT 22.485000 60.360000 22.685000 60.560000 ;
        RECT 22.485000 60.770000 22.685000 60.970000 ;
        RECT 22.485000 61.180000 22.685000 61.380000 ;
        RECT 22.485000 61.590000 22.685000 61.790000 ;
        RECT 22.485000 62.000000 22.685000 62.200000 ;
        RECT 22.485000 62.410000 22.685000 62.610000 ;
        RECT 22.890000 58.310000 23.090000 58.510000 ;
        RECT 22.890000 58.720000 23.090000 58.920000 ;
        RECT 22.890000 59.130000 23.090000 59.330000 ;
        RECT 22.890000 59.540000 23.090000 59.740000 ;
        RECT 22.890000 59.950000 23.090000 60.150000 ;
        RECT 22.890000 60.360000 23.090000 60.560000 ;
        RECT 22.890000 60.770000 23.090000 60.970000 ;
        RECT 22.890000 61.180000 23.090000 61.380000 ;
        RECT 22.890000 61.590000 23.090000 61.790000 ;
        RECT 22.890000 62.000000 23.090000 62.200000 ;
        RECT 22.890000 62.410000 23.090000 62.610000 ;
        RECT 23.295000 58.310000 23.495000 58.510000 ;
        RECT 23.295000 58.720000 23.495000 58.920000 ;
        RECT 23.295000 59.130000 23.495000 59.330000 ;
        RECT 23.295000 59.540000 23.495000 59.740000 ;
        RECT 23.295000 59.950000 23.495000 60.150000 ;
        RECT 23.295000 60.360000 23.495000 60.560000 ;
        RECT 23.295000 60.770000 23.495000 60.970000 ;
        RECT 23.295000 61.180000 23.495000 61.380000 ;
        RECT 23.295000 61.590000 23.495000 61.790000 ;
        RECT 23.295000 62.000000 23.495000 62.200000 ;
        RECT 23.295000 62.410000 23.495000 62.610000 ;
        RECT 23.700000 58.310000 23.900000 58.510000 ;
        RECT 23.700000 58.720000 23.900000 58.920000 ;
        RECT 23.700000 59.130000 23.900000 59.330000 ;
        RECT 23.700000 59.540000 23.900000 59.740000 ;
        RECT 23.700000 59.950000 23.900000 60.150000 ;
        RECT 23.700000 60.360000 23.900000 60.560000 ;
        RECT 23.700000 60.770000 23.900000 60.970000 ;
        RECT 23.700000 61.180000 23.900000 61.380000 ;
        RECT 23.700000 61.590000 23.900000 61.790000 ;
        RECT 23.700000 62.000000 23.900000 62.200000 ;
        RECT 23.700000 62.410000 23.900000 62.610000 ;
        RECT 24.105000 58.310000 24.305000 58.510000 ;
        RECT 24.105000 58.720000 24.305000 58.920000 ;
        RECT 24.105000 59.130000 24.305000 59.330000 ;
        RECT 24.105000 59.540000 24.305000 59.740000 ;
        RECT 24.105000 59.950000 24.305000 60.150000 ;
        RECT 24.105000 60.360000 24.305000 60.560000 ;
        RECT 24.105000 60.770000 24.305000 60.970000 ;
        RECT 24.105000 61.180000 24.305000 61.380000 ;
        RECT 24.105000 61.590000 24.305000 61.790000 ;
        RECT 24.105000 62.000000 24.305000 62.200000 ;
        RECT 24.105000 62.410000 24.305000 62.610000 ;
        RECT 50.480000 58.310000 50.680000 58.510000 ;
        RECT 50.480000 58.720000 50.680000 58.920000 ;
        RECT 50.480000 59.130000 50.680000 59.330000 ;
        RECT 50.480000 59.540000 50.680000 59.740000 ;
        RECT 50.480000 59.950000 50.680000 60.150000 ;
        RECT 50.480000 60.360000 50.680000 60.560000 ;
        RECT 50.480000 60.770000 50.680000 60.970000 ;
        RECT 50.480000 61.180000 50.680000 61.380000 ;
        RECT 50.480000 61.590000 50.680000 61.790000 ;
        RECT 50.480000 62.000000 50.680000 62.200000 ;
        RECT 50.480000 62.410000 50.680000 62.610000 ;
        RECT 50.890000 58.310000 51.090000 58.510000 ;
        RECT 50.890000 58.720000 51.090000 58.920000 ;
        RECT 50.890000 59.130000 51.090000 59.330000 ;
        RECT 50.890000 59.540000 51.090000 59.740000 ;
        RECT 50.890000 59.950000 51.090000 60.150000 ;
        RECT 50.890000 60.360000 51.090000 60.560000 ;
        RECT 50.890000 60.770000 51.090000 60.970000 ;
        RECT 50.890000 61.180000 51.090000 61.380000 ;
        RECT 50.890000 61.590000 51.090000 61.790000 ;
        RECT 50.890000 62.000000 51.090000 62.200000 ;
        RECT 50.890000 62.410000 51.090000 62.610000 ;
        RECT 51.300000 58.310000 51.500000 58.510000 ;
        RECT 51.300000 58.720000 51.500000 58.920000 ;
        RECT 51.300000 59.130000 51.500000 59.330000 ;
        RECT 51.300000 59.540000 51.500000 59.740000 ;
        RECT 51.300000 59.950000 51.500000 60.150000 ;
        RECT 51.300000 60.360000 51.500000 60.560000 ;
        RECT 51.300000 60.770000 51.500000 60.970000 ;
        RECT 51.300000 61.180000 51.500000 61.380000 ;
        RECT 51.300000 61.590000 51.500000 61.790000 ;
        RECT 51.300000 62.000000 51.500000 62.200000 ;
        RECT 51.300000 62.410000 51.500000 62.610000 ;
        RECT 51.710000 58.310000 51.910000 58.510000 ;
        RECT 51.710000 58.720000 51.910000 58.920000 ;
        RECT 51.710000 59.130000 51.910000 59.330000 ;
        RECT 51.710000 59.540000 51.910000 59.740000 ;
        RECT 51.710000 59.950000 51.910000 60.150000 ;
        RECT 51.710000 60.360000 51.910000 60.560000 ;
        RECT 51.710000 60.770000 51.910000 60.970000 ;
        RECT 51.710000 61.180000 51.910000 61.380000 ;
        RECT 51.710000 61.590000 51.910000 61.790000 ;
        RECT 51.710000 62.000000 51.910000 62.200000 ;
        RECT 51.710000 62.410000 51.910000 62.610000 ;
        RECT 52.120000 58.310000 52.320000 58.510000 ;
        RECT 52.120000 58.720000 52.320000 58.920000 ;
        RECT 52.120000 59.130000 52.320000 59.330000 ;
        RECT 52.120000 59.540000 52.320000 59.740000 ;
        RECT 52.120000 59.950000 52.320000 60.150000 ;
        RECT 52.120000 60.360000 52.320000 60.560000 ;
        RECT 52.120000 60.770000 52.320000 60.970000 ;
        RECT 52.120000 61.180000 52.320000 61.380000 ;
        RECT 52.120000 61.590000 52.320000 61.790000 ;
        RECT 52.120000 62.000000 52.320000 62.200000 ;
        RECT 52.120000 62.410000 52.320000 62.610000 ;
        RECT 52.530000 58.310000 52.730000 58.510000 ;
        RECT 52.530000 58.720000 52.730000 58.920000 ;
        RECT 52.530000 59.130000 52.730000 59.330000 ;
        RECT 52.530000 59.540000 52.730000 59.740000 ;
        RECT 52.530000 59.950000 52.730000 60.150000 ;
        RECT 52.530000 60.360000 52.730000 60.560000 ;
        RECT 52.530000 60.770000 52.730000 60.970000 ;
        RECT 52.530000 61.180000 52.730000 61.380000 ;
        RECT 52.530000 61.590000 52.730000 61.790000 ;
        RECT 52.530000 62.000000 52.730000 62.200000 ;
        RECT 52.530000 62.410000 52.730000 62.610000 ;
        RECT 52.940000 58.310000 53.140000 58.510000 ;
        RECT 52.940000 58.720000 53.140000 58.920000 ;
        RECT 52.940000 59.130000 53.140000 59.330000 ;
        RECT 52.940000 59.540000 53.140000 59.740000 ;
        RECT 52.940000 59.950000 53.140000 60.150000 ;
        RECT 52.940000 60.360000 53.140000 60.560000 ;
        RECT 52.940000 60.770000 53.140000 60.970000 ;
        RECT 52.940000 61.180000 53.140000 61.380000 ;
        RECT 52.940000 61.590000 53.140000 61.790000 ;
        RECT 52.940000 62.000000 53.140000 62.200000 ;
        RECT 52.940000 62.410000 53.140000 62.610000 ;
        RECT 53.345000 58.310000 53.545000 58.510000 ;
        RECT 53.345000 58.720000 53.545000 58.920000 ;
        RECT 53.345000 59.130000 53.545000 59.330000 ;
        RECT 53.345000 59.540000 53.545000 59.740000 ;
        RECT 53.345000 59.950000 53.545000 60.150000 ;
        RECT 53.345000 60.360000 53.545000 60.560000 ;
        RECT 53.345000 60.770000 53.545000 60.970000 ;
        RECT 53.345000 61.180000 53.545000 61.380000 ;
        RECT 53.345000 61.590000 53.545000 61.790000 ;
        RECT 53.345000 62.000000 53.545000 62.200000 ;
        RECT 53.345000 62.410000 53.545000 62.610000 ;
        RECT 53.750000 58.310000 53.950000 58.510000 ;
        RECT 53.750000 58.720000 53.950000 58.920000 ;
        RECT 53.750000 59.130000 53.950000 59.330000 ;
        RECT 53.750000 59.540000 53.950000 59.740000 ;
        RECT 53.750000 59.950000 53.950000 60.150000 ;
        RECT 53.750000 60.360000 53.950000 60.560000 ;
        RECT 53.750000 60.770000 53.950000 60.970000 ;
        RECT 53.750000 61.180000 53.950000 61.380000 ;
        RECT 53.750000 61.590000 53.950000 61.790000 ;
        RECT 53.750000 62.000000 53.950000 62.200000 ;
        RECT 53.750000 62.410000 53.950000 62.610000 ;
        RECT 54.155000 58.310000 54.355000 58.510000 ;
        RECT 54.155000 58.720000 54.355000 58.920000 ;
        RECT 54.155000 59.130000 54.355000 59.330000 ;
        RECT 54.155000 59.540000 54.355000 59.740000 ;
        RECT 54.155000 59.950000 54.355000 60.150000 ;
        RECT 54.155000 60.360000 54.355000 60.560000 ;
        RECT 54.155000 60.770000 54.355000 60.970000 ;
        RECT 54.155000 61.180000 54.355000 61.380000 ;
        RECT 54.155000 61.590000 54.355000 61.790000 ;
        RECT 54.155000 62.000000 54.355000 62.200000 ;
        RECT 54.155000 62.410000 54.355000 62.610000 ;
        RECT 54.560000 58.310000 54.760000 58.510000 ;
        RECT 54.560000 58.720000 54.760000 58.920000 ;
        RECT 54.560000 59.130000 54.760000 59.330000 ;
        RECT 54.560000 59.540000 54.760000 59.740000 ;
        RECT 54.560000 59.950000 54.760000 60.150000 ;
        RECT 54.560000 60.360000 54.760000 60.560000 ;
        RECT 54.560000 60.770000 54.760000 60.970000 ;
        RECT 54.560000 61.180000 54.760000 61.380000 ;
        RECT 54.560000 61.590000 54.760000 61.790000 ;
        RECT 54.560000 62.000000 54.760000 62.200000 ;
        RECT 54.560000 62.410000 54.760000 62.610000 ;
        RECT 54.965000 58.310000 55.165000 58.510000 ;
        RECT 54.965000 58.720000 55.165000 58.920000 ;
        RECT 54.965000 59.130000 55.165000 59.330000 ;
        RECT 54.965000 59.540000 55.165000 59.740000 ;
        RECT 54.965000 59.950000 55.165000 60.150000 ;
        RECT 54.965000 60.360000 55.165000 60.560000 ;
        RECT 54.965000 60.770000 55.165000 60.970000 ;
        RECT 54.965000 61.180000 55.165000 61.380000 ;
        RECT 54.965000 61.590000 55.165000 61.790000 ;
        RECT 54.965000 62.000000 55.165000 62.200000 ;
        RECT 54.965000 62.410000 55.165000 62.610000 ;
        RECT 55.370000 58.310000 55.570000 58.510000 ;
        RECT 55.370000 58.720000 55.570000 58.920000 ;
        RECT 55.370000 59.130000 55.570000 59.330000 ;
        RECT 55.370000 59.540000 55.570000 59.740000 ;
        RECT 55.370000 59.950000 55.570000 60.150000 ;
        RECT 55.370000 60.360000 55.570000 60.560000 ;
        RECT 55.370000 60.770000 55.570000 60.970000 ;
        RECT 55.370000 61.180000 55.570000 61.380000 ;
        RECT 55.370000 61.590000 55.570000 61.790000 ;
        RECT 55.370000 62.000000 55.570000 62.200000 ;
        RECT 55.370000 62.410000 55.570000 62.610000 ;
        RECT 55.775000 58.310000 55.975000 58.510000 ;
        RECT 55.775000 58.720000 55.975000 58.920000 ;
        RECT 55.775000 59.130000 55.975000 59.330000 ;
        RECT 55.775000 59.540000 55.975000 59.740000 ;
        RECT 55.775000 59.950000 55.975000 60.150000 ;
        RECT 55.775000 60.360000 55.975000 60.560000 ;
        RECT 55.775000 60.770000 55.975000 60.970000 ;
        RECT 55.775000 61.180000 55.975000 61.380000 ;
        RECT 55.775000 61.590000 55.975000 61.790000 ;
        RECT 55.775000 62.000000 55.975000 62.200000 ;
        RECT 55.775000 62.410000 55.975000 62.610000 ;
        RECT 56.180000 58.310000 56.380000 58.510000 ;
        RECT 56.180000 58.720000 56.380000 58.920000 ;
        RECT 56.180000 59.130000 56.380000 59.330000 ;
        RECT 56.180000 59.540000 56.380000 59.740000 ;
        RECT 56.180000 59.950000 56.380000 60.150000 ;
        RECT 56.180000 60.360000 56.380000 60.560000 ;
        RECT 56.180000 60.770000 56.380000 60.970000 ;
        RECT 56.180000 61.180000 56.380000 61.380000 ;
        RECT 56.180000 61.590000 56.380000 61.790000 ;
        RECT 56.180000 62.000000 56.380000 62.200000 ;
        RECT 56.180000 62.410000 56.380000 62.610000 ;
        RECT 56.585000 58.310000 56.785000 58.510000 ;
        RECT 56.585000 58.720000 56.785000 58.920000 ;
        RECT 56.585000 59.130000 56.785000 59.330000 ;
        RECT 56.585000 59.540000 56.785000 59.740000 ;
        RECT 56.585000 59.950000 56.785000 60.150000 ;
        RECT 56.585000 60.360000 56.785000 60.560000 ;
        RECT 56.585000 60.770000 56.785000 60.970000 ;
        RECT 56.585000 61.180000 56.785000 61.380000 ;
        RECT 56.585000 61.590000 56.785000 61.790000 ;
        RECT 56.585000 62.000000 56.785000 62.200000 ;
        RECT 56.585000 62.410000 56.785000 62.610000 ;
        RECT 56.990000 58.310000 57.190000 58.510000 ;
        RECT 56.990000 58.720000 57.190000 58.920000 ;
        RECT 56.990000 59.130000 57.190000 59.330000 ;
        RECT 56.990000 59.540000 57.190000 59.740000 ;
        RECT 56.990000 59.950000 57.190000 60.150000 ;
        RECT 56.990000 60.360000 57.190000 60.560000 ;
        RECT 56.990000 60.770000 57.190000 60.970000 ;
        RECT 56.990000 61.180000 57.190000 61.380000 ;
        RECT 56.990000 61.590000 57.190000 61.790000 ;
        RECT 56.990000 62.000000 57.190000 62.200000 ;
        RECT 56.990000 62.410000 57.190000 62.610000 ;
        RECT 57.395000 58.310000 57.595000 58.510000 ;
        RECT 57.395000 58.720000 57.595000 58.920000 ;
        RECT 57.395000 59.130000 57.595000 59.330000 ;
        RECT 57.395000 59.540000 57.595000 59.740000 ;
        RECT 57.395000 59.950000 57.595000 60.150000 ;
        RECT 57.395000 60.360000 57.595000 60.560000 ;
        RECT 57.395000 60.770000 57.595000 60.970000 ;
        RECT 57.395000 61.180000 57.595000 61.380000 ;
        RECT 57.395000 61.590000 57.595000 61.790000 ;
        RECT 57.395000 62.000000 57.595000 62.200000 ;
        RECT 57.395000 62.410000 57.595000 62.610000 ;
        RECT 57.800000 58.310000 58.000000 58.510000 ;
        RECT 57.800000 58.720000 58.000000 58.920000 ;
        RECT 57.800000 59.130000 58.000000 59.330000 ;
        RECT 57.800000 59.540000 58.000000 59.740000 ;
        RECT 57.800000 59.950000 58.000000 60.150000 ;
        RECT 57.800000 60.360000 58.000000 60.560000 ;
        RECT 57.800000 60.770000 58.000000 60.970000 ;
        RECT 57.800000 61.180000 58.000000 61.380000 ;
        RECT 57.800000 61.590000 58.000000 61.790000 ;
        RECT 57.800000 62.000000 58.000000 62.200000 ;
        RECT 57.800000 62.410000 58.000000 62.610000 ;
        RECT 58.205000 58.310000 58.405000 58.510000 ;
        RECT 58.205000 58.720000 58.405000 58.920000 ;
        RECT 58.205000 59.130000 58.405000 59.330000 ;
        RECT 58.205000 59.540000 58.405000 59.740000 ;
        RECT 58.205000 59.950000 58.405000 60.150000 ;
        RECT 58.205000 60.360000 58.405000 60.560000 ;
        RECT 58.205000 60.770000 58.405000 60.970000 ;
        RECT 58.205000 61.180000 58.405000 61.380000 ;
        RECT 58.205000 61.590000 58.405000 61.790000 ;
        RECT 58.205000 62.000000 58.405000 62.200000 ;
        RECT 58.205000 62.410000 58.405000 62.610000 ;
        RECT 58.610000 58.310000 58.810000 58.510000 ;
        RECT 58.610000 58.720000 58.810000 58.920000 ;
        RECT 58.610000 59.130000 58.810000 59.330000 ;
        RECT 58.610000 59.540000 58.810000 59.740000 ;
        RECT 58.610000 59.950000 58.810000 60.150000 ;
        RECT 58.610000 60.360000 58.810000 60.560000 ;
        RECT 58.610000 60.770000 58.810000 60.970000 ;
        RECT 58.610000 61.180000 58.810000 61.380000 ;
        RECT 58.610000 61.590000 58.810000 61.790000 ;
        RECT 58.610000 62.000000 58.810000 62.200000 ;
        RECT 58.610000 62.410000 58.810000 62.610000 ;
        RECT 59.015000 58.310000 59.215000 58.510000 ;
        RECT 59.015000 58.720000 59.215000 58.920000 ;
        RECT 59.015000 59.130000 59.215000 59.330000 ;
        RECT 59.015000 59.540000 59.215000 59.740000 ;
        RECT 59.015000 59.950000 59.215000 60.150000 ;
        RECT 59.015000 60.360000 59.215000 60.560000 ;
        RECT 59.015000 60.770000 59.215000 60.970000 ;
        RECT 59.015000 61.180000 59.215000 61.380000 ;
        RECT 59.015000 61.590000 59.215000 61.790000 ;
        RECT 59.015000 62.000000 59.215000 62.200000 ;
        RECT 59.015000 62.410000 59.215000 62.610000 ;
        RECT 59.420000 58.310000 59.620000 58.510000 ;
        RECT 59.420000 58.720000 59.620000 58.920000 ;
        RECT 59.420000 59.130000 59.620000 59.330000 ;
        RECT 59.420000 59.540000 59.620000 59.740000 ;
        RECT 59.420000 59.950000 59.620000 60.150000 ;
        RECT 59.420000 60.360000 59.620000 60.560000 ;
        RECT 59.420000 60.770000 59.620000 60.970000 ;
        RECT 59.420000 61.180000 59.620000 61.380000 ;
        RECT 59.420000 61.590000 59.620000 61.790000 ;
        RECT 59.420000 62.000000 59.620000 62.200000 ;
        RECT 59.420000 62.410000 59.620000 62.610000 ;
        RECT 59.825000 58.310000 60.025000 58.510000 ;
        RECT 59.825000 58.720000 60.025000 58.920000 ;
        RECT 59.825000 59.130000 60.025000 59.330000 ;
        RECT 59.825000 59.540000 60.025000 59.740000 ;
        RECT 59.825000 59.950000 60.025000 60.150000 ;
        RECT 59.825000 60.360000 60.025000 60.560000 ;
        RECT 59.825000 60.770000 60.025000 60.970000 ;
        RECT 59.825000 61.180000 60.025000 61.380000 ;
        RECT 59.825000 61.590000 60.025000 61.790000 ;
        RECT 59.825000 62.000000 60.025000 62.200000 ;
        RECT 59.825000 62.410000 60.025000 62.610000 ;
        RECT 60.230000 58.310000 60.430000 58.510000 ;
        RECT 60.230000 58.720000 60.430000 58.920000 ;
        RECT 60.230000 59.130000 60.430000 59.330000 ;
        RECT 60.230000 59.540000 60.430000 59.740000 ;
        RECT 60.230000 59.950000 60.430000 60.150000 ;
        RECT 60.230000 60.360000 60.430000 60.560000 ;
        RECT 60.230000 60.770000 60.430000 60.970000 ;
        RECT 60.230000 61.180000 60.430000 61.380000 ;
        RECT 60.230000 61.590000 60.430000 61.790000 ;
        RECT 60.230000 62.000000 60.430000 62.200000 ;
        RECT 60.230000 62.410000 60.430000 62.610000 ;
        RECT 60.635000 58.310000 60.835000 58.510000 ;
        RECT 60.635000 58.720000 60.835000 58.920000 ;
        RECT 60.635000 59.130000 60.835000 59.330000 ;
        RECT 60.635000 59.540000 60.835000 59.740000 ;
        RECT 60.635000 59.950000 60.835000 60.150000 ;
        RECT 60.635000 60.360000 60.835000 60.560000 ;
        RECT 60.635000 60.770000 60.835000 60.970000 ;
        RECT 60.635000 61.180000 60.835000 61.380000 ;
        RECT 60.635000 61.590000 60.835000 61.790000 ;
        RECT 60.635000 62.000000 60.835000 62.200000 ;
        RECT 60.635000 62.410000 60.835000 62.610000 ;
        RECT 61.040000 58.310000 61.240000 58.510000 ;
        RECT 61.040000 58.720000 61.240000 58.920000 ;
        RECT 61.040000 59.130000 61.240000 59.330000 ;
        RECT 61.040000 59.540000 61.240000 59.740000 ;
        RECT 61.040000 59.950000 61.240000 60.150000 ;
        RECT 61.040000 60.360000 61.240000 60.560000 ;
        RECT 61.040000 60.770000 61.240000 60.970000 ;
        RECT 61.040000 61.180000 61.240000 61.380000 ;
        RECT 61.040000 61.590000 61.240000 61.790000 ;
        RECT 61.040000 62.000000 61.240000 62.200000 ;
        RECT 61.040000 62.410000 61.240000 62.610000 ;
        RECT 61.445000 58.310000 61.645000 58.510000 ;
        RECT 61.445000 58.720000 61.645000 58.920000 ;
        RECT 61.445000 59.130000 61.645000 59.330000 ;
        RECT 61.445000 59.540000 61.645000 59.740000 ;
        RECT 61.445000 59.950000 61.645000 60.150000 ;
        RECT 61.445000 60.360000 61.645000 60.560000 ;
        RECT 61.445000 60.770000 61.645000 60.970000 ;
        RECT 61.445000 61.180000 61.645000 61.380000 ;
        RECT 61.445000 61.590000 61.645000 61.790000 ;
        RECT 61.445000 62.000000 61.645000 62.200000 ;
        RECT 61.445000 62.410000 61.645000 62.610000 ;
        RECT 61.850000 58.310000 62.050000 58.510000 ;
        RECT 61.850000 58.720000 62.050000 58.920000 ;
        RECT 61.850000 59.130000 62.050000 59.330000 ;
        RECT 61.850000 59.540000 62.050000 59.740000 ;
        RECT 61.850000 59.950000 62.050000 60.150000 ;
        RECT 61.850000 60.360000 62.050000 60.560000 ;
        RECT 61.850000 60.770000 62.050000 60.970000 ;
        RECT 61.850000 61.180000 62.050000 61.380000 ;
        RECT 61.850000 61.590000 62.050000 61.790000 ;
        RECT 61.850000 62.000000 62.050000 62.200000 ;
        RECT 61.850000 62.410000 62.050000 62.610000 ;
        RECT 62.255000 58.310000 62.455000 58.510000 ;
        RECT 62.255000 58.720000 62.455000 58.920000 ;
        RECT 62.255000 59.130000 62.455000 59.330000 ;
        RECT 62.255000 59.540000 62.455000 59.740000 ;
        RECT 62.255000 59.950000 62.455000 60.150000 ;
        RECT 62.255000 60.360000 62.455000 60.560000 ;
        RECT 62.255000 60.770000 62.455000 60.970000 ;
        RECT 62.255000 61.180000 62.455000 61.380000 ;
        RECT 62.255000 61.590000 62.455000 61.790000 ;
        RECT 62.255000 62.000000 62.455000 62.200000 ;
        RECT 62.255000 62.410000 62.455000 62.610000 ;
        RECT 62.660000 58.310000 62.860000 58.510000 ;
        RECT 62.660000 58.720000 62.860000 58.920000 ;
        RECT 62.660000 59.130000 62.860000 59.330000 ;
        RECT 62.660000 59.540000 62.860000 59.740000 ;
        RECT 62.660000 59.950000 62.860000 60.150000 ;
        RECT 62.660000 60.360000 62.860000 60.560000 ;
        RECT 62.660000 60.770000 62.860000 60.970000 ;
        RECT 62.660000 61.180000 62.860000 61.380000 ;
        RECT 62.660000 61.590000 62.860000 61.790000 ;
        RECT 62.660000 62.000000 62.860000 62.200000 ;
        RECT 62.660000 62.410000 62.860000 62.610000 ;
        RECT 63.065000 58.310000 63.265000 58.510000 ;
        RECT 63.065000 58.720000 63.265000 58.920000 ;
        RECT 63.065000 59.130000 63.265000 59.330000 ;
        RECT 63.065000 59.540000 63.265000 59.740000 ;
        RECT 63.065000 59.950000 63.265000 60.150000 ;
        RECT 63.065000 60.360000 63.265000 60.560000 ;
        RECT 63.065000 60.770000 63.265000 60.970000 ;
        RECT 63.065000 61.180000 63.265000 61.380000 ;
        RECT 63.065000 61.590000 63.265000 61.790000 ;
        RECT 63.065000 62.000000 63.265000 62.200000 ;
        RECT 63.065000 62.410000 63.265000 62.610000 ;
        RECT 63.470000 58.310000 63.670000 58.510000 ;
        RECT 63.470000 58.720000 63.670000 58.920000 ;
        RECT 63.470000 59.130000 63.670000 59.330000 ;
        RECT 63.470000 59.540000 63.670000 59.740000 ;
        RECT 63.470000 59.950000 63.670000 60.150000 ;
        RECT 63.470000 60.360000 63.670000 60.560000 ;
        RECT 63.470000 60.770000 63.670000 60.970000 ;
        RECT 63.470000 61.180000 63.670000 61.380000 ;
        RECT 63.470000 61.590000 63.670000 61.790000 ;
        RECT 63.470000 62.000000 63.670000 62.200000 ;
        RECT 63.470000 62.410000 63.670000 62.610000 ;
        RECT 63.875000 58.310000 64.075000 58.510000 ;
        RECT 63.875000 58.720000 64.075000 58.920000 ;
        RECT 63.875000 59.130000 64.075000 59.330000 ;
        RECT 63.875000 59.540000 64.075000 59.740000 ;
        RECT 63.875000 59.950000 64.075000 60.150000 ;
        RECT 63.875000 60.360000 64.075000 60.560000 ;
        RECT 63.875000 60.770000 64.075000 60.970000 ;
        RECT 63.875000 61.180000 64.075000 61.380000 ;
        RECT 63.875000 61.590000 64.075000 61.790000 ;
        RECT 63.875000 62.000000 64.075000 62.200000 ;
        RECT 63.875000 62.410000 64.075000 62.610000 ;
        RECT 64.280000 58.310000 64.480000 58.510000 ;
        RECT 64.280000 58.720000 64.480000 58.920000 ;
        RECT 64.280000 59.130000 64.480000 59.330000 ;
        RECT 64.280000 59.540000 64.480000 59.740000 ;
        RECT 64.280000 59.950000 64.480000 60.150000 ;
        RECT 64.280000 60.360000 64.480000 60.560000 ;
        RECT 64.280000 60.770000 64.480000 60.970000 ;
        RECT 64.280000 61.180000 64.480000 61.380000 ;
        RECT 64.280000 61.590000 64.480000 61.790000 ;
        RECT 64.280000 62.000000 64.480000 62.200000 ;
        RECT 64.280000 62.410000 64.480000 62.610000 ;
        RECT 64.685000 58.310000 64.885000 58.510000 ;
        RECT 64.685000 58.720000 64.885000 58.920000 ;
        RECT 64.685000 59.130000 64.885000 59.330000 ;
        RECT 64.685000 59.540000 64.885000 59.740000 ;
        RECT 64.685000 59.950000 64.885000 60.150000 ;
        RECT 64.685000 60.360000 64.885000 60.560000 ;
        RECT 64.685000 60.770000 64.885000 60.970000 ;
        RECT 64.685000 61.180000 64.885000 61.380000 ;
        RECT 64.685000 61.590000 64.885000 61.790000 ;
        RECT 64.685000 62.000000 64.885000 62.200000 ;
        RECT 64.685000 62.410000 64.885000 62.610000 ;
        RECT 65.090000 58.310000 65.290000 58.510000 ;
        RECT 65.090000 58.720000 65.290000 58.920000 ;
        RECT 65.090000 59.130000 65.290000 59.330000 ;
        RECT 65.090000 59.540000 65.290000 59.740000 ;
        RECT 65.090000 59.950000 65.290000 60.150000 ;
        RECT 65.090000 60.360000 65.290000 60.560000 ;
        RECT 65.090000 60.770000 65.290000 60.970000 ;
        RECT 65.090000 61.180000 65.290000 61.380000 ;
        RECT 65.090000 61.590000 65.290000 61.790000 ;
        RECT 65.090000 62.000000 65.290000 62.200000 ;
        RECT 65.090000 62.410000 65.290000 62.610000 ;
        RECT 65.495000 58.310000 65.695000 58.510000 ;
        RECT 65.495000 58.720000 65.695000 58.920000 ;
        RECT 65.495000 59.130000 65.695000 59.330000 ;
        RECT 65.495000 59.540000 65.695000 59.740000 ;
        RECT 65.495000 59.950000 65.695000 60.150000 ;
        RECT 65.495000 60.360000 65.695000 60.560000 ;
        RECT 65.495000 60.770000 65.695000 60.970000 ;
        RECT 65.495000 61.180000 65.695000 61.380000 ;
        RECT 65.495000 61.590000 65.695000 61.790000 ;
        RECT 65.495000 62.000000 65.695000 62.200000 ;
        RECT 65.495000 62.410000 65.695000 62.610000 ;
        RECT 65.900000 58.310000 66.100000 58.510000 ;
        RECT 65.900000 58.720000 66.100000 58.920000 ;
        RECT 65.900000 59.130000 66.100000 59.330000 ;
        RECT 65.900000 59.540000 66.100000 59.740000 ;
        RECT 65.900000 59.950000 66.100000 60.150000 ;
        RECT 65.900000 60.360000 66.100000 60.560000 ;
        RECT 65.900000 60.770000 66.100000 60.970000 ;
        RECT 65.900000 61.180000 66.100000 61.380000 ;
        RECT 65.900000 61.590000 66.100000 61.790000 ;
        RECT 65.900000 62.000000 66.100000 62.200000 ;
        RECT 65.900000 62.410000 66.100000 62.610000 ;
        RECT 66.305000 58.310000 66.505000 58.510000 ;
        RECT 66.305000 58.720000 66.505000 58.920000 ;
        RECT 66.305000 59.130000 66.505000 59.330000 ;
        RECT 66.305000 59.540000 66.505000 59.740000 ;
        RECT 66.305000 59.950000 66.505000 60.150000 ;
        RECT 66.305000 60.360000 66.505000 60.560000 ;
        RECT 66.305000 60.770000 66.505000 60.970000 ;
        RECT 66.305000 61.180000 66.505000 61.380000 ;
        RECT 66.305000 61.590000 66.505000 61.790000 ;
        RECT 66.305000 62.000000 66.505000 62.200000 ;
        RECT 66.305000 62.410000 66.505000 62.610000 ;
        RECT 66.710000 58.310000 66.910000 58.510000 ;
        RECT 66.710000 58.720000 66.910000 58.920000 ;
        RECT 66.710000 59.130000 66.910000 59.330000 ;
        RECT 66.710000 59.540000 66.910000 59.740000 ;
        RECT 66.710000 59.950000 66.910000 60.150000 ;
        RECT 66.710000 60.360000 66.910000 60.560000 ;
        RECT 66.710000 60.770000 66.910000 60.970000 ;
        RECT 66.710000 61.180000 66.910000 61.380000 ;
        RECT 66.710000 61.590000 66.910000 61.790000 ;
        RECT 66.710000 62.000000 66.910000 62.200000 ;
        RECT 66.710000 62.410000 66.910000 62.610000 ;
        RECT 67.115000 58.310000 67.315000 58.510000 ;
        RECT 67.115000 58.720000 67.315000 58.920000 ;
        RECT 67.115000 59.130000 67.315000 59.330000 ;
        RECT 67.115000 59.540000 67.315000 59.740000 ;
        RECT 67.115000 59.950000 67.315000 60.150000 ;
        RECT 67.115000 60.360000 67.315000 60.560000 ;
        RECT 67.115000 60.770000 67.315000 60.970000 ;
        RECT 67.115000 61.180000 67.315000 61.380000 ;
        RECT 67.115000 61.590000 67.315000 61.790000 ;
        RECT 67.115000 62.000000 67.315000 62.200000 ;
        RECT 67.115000 62.410000 67.315000 62.610000 ;
        RECT 67.520000 58.310000 67.720000 58.510000 ;
        RECT 67.520000 58.720000 67.720000 58.920000 ;
        RECT 67.520000 59.130000 67.720000 59.330000 ;
        RECT 67.520000 59.540000 67.720000 59.740000 ;
        RECT 67.520000 59.950000 67.720000 60.150000 ;
        RECT 67.520000 60.360000 67.720000 60.560000 ;
        RECT 67.520000 60.770000 67.720000 60.970000 ;
        RECT 67.520000 61.180000 67.720000 61.380000 ;
        RECT 67.520000 61.590000 67.720000 61.790000 ;
        RECT 67.520000 62.000000 67.720000 62.200000 ;
        RECT 67.520000 62.410000 67.720000 62.610000 ;
        RECT 67.925000 58.310000 68.125000 58.510000 ;
        RECT 67.925000 58.720000 68.125000 58.920000 ;
        RECT 67.925000 59.130000 68.125000 59.330000 ;
        RECT 67.925000 59.540000 68.125000 59.740000 ;
        RECT 67.925000 59.950000 68.125000 60.150000 ;
        RECT 67.925000 60.360000 68.125000 60.560000 ;
        RECT 67.925000 60.770000 68.125000 60.970000 ;
        RECT 67.925000 61.180000 68.125000 61.380000 ;
        RECT 67.925000 61.590000 68.125000 61.790000 ;
        RECT 67.925000 62.000000 68.125000 62.200000 ;
        RECT 67.925000 62.410000 68.125000 62.610000 ;
        RECT 68.330000 58.310000 68.530000 58.510000 ;
        RECT 68.330000 58.720000 68.530000 58.920000 ;
        RECT 68.330000 59.130000 68.530000 59.330000 ;
        RECT 68.330000 59.540000 68.530000 59.740000 ;
        RECT 68.330000 59.950000 68.530000 60.150000 ;
        RECT 68.330000 60.360000 68.530000 60.560000 ;
        RECT 68.330000 60.770000 68.530000 60.970000 ;
        RECT 68.330000 61.180000 68.530000 61.380000 ;
        RECT 68.330000 61.590000 68.530000 61.790000 ;
        RECT 68.330000 62.000000 68.530000 62.200000 ;
        RECT 68.330000 62.410000 68.530000 62.610000 ;
        RECT 68.735000 58.310000 68.935000 58.510000 ;
        RECT 68.735000 58.720000 68.935000 58.920000 ;
        RECT 68.735000 59.130000 68.935000 59.330000 ;
        RECT 68.735000 59.540000 68.935000 59.740000 ;
        RECT 68.735000 59.950000 68.935000 60.150000 ;
        RECT 68.735000 60.360000 68.935000 60.560000 ;
        RECT 68.735000 60.770000 68.935000 60.970000 ;
        RECT 68.735000 61.180000 68.935000 61.380000 ;
        RECT 68.735000 61.590000 68.935000 61.790000 ;
        RECT 68.735000 62.000000 68.935000 62.200000 ;
        RECT 68.735000 62.410000 68.935000 62.610000 ;
        RECT 69.140000 58.310000 69.340000 58.510000 ;
        RECT 69.140000 58.720000 69.340000 58.920000 ;
        RECT 69.140000 59.130000 69.340000 59.330000 ;
        RECT 69.140000 59.540000 69.340000 59.740000 ;
        RECT 69.140000 59.950000 69.340000 60.150000 ;
        RECT 69.140000 60.360000 69.340000 60.560000 ;
        RECT 69.140000 60.770000 69.340000 60.970000 ;
        RECT 69.140000 61.180000 69.340000 61.380000 ;
        RECT 69.140000 61.590000 69.340000 61.790000 ;
        RECT 69.140000 62.000000 69.340000 62.200000 ;
        RECT 69.140000 62.410000 69.340000 62.610000 ;
        RECT 69.545000 58.310000 69.745000 58.510000 ;
        RECT 69.545000 58.720000 69.745000 58.920000 ;
        RECT 69.545000 59.130000 69.745000 59.330000 ;
        RECT 69.545000 59.540000 69.745000 59.740000 ;
        RECT 69.545000 59.950000 69.745000 60.150000 ;
        RECT 69.545000 60.360000 69.745000 60.560000 ;
        RECT 69.545000 60.770000 69.745000 60.970000 ;
        RECT 69.545000 61.180000 69.745000 61.380000 ;
        RECT 69.545000 61.590000 69.745000 61.790000 ;
        RECT 69.545000 62.000000 69.745000 62.200000 ;
        RECT 69.545000 62.410000 69.745000 62.610000 ;
        RECT 69.950000 58.310000 70.150000 58.510000 ;
        RECT 69.950000 58.720000 70.150000 58.920000 ;
        RECT 69.950000 59.130000 70.150000 59.330000 ;
        RECT 69.950000 59.540000 70.150000 59.740000 ;
        RECT 69.950000 59.950000 70.150000 60.150000 ;
        RECT 69.950000 60.360000 70.150000 60.560000 ;
        RECT 69.950000 60.770000 70.150000 60.970000 ;
        RECT 69.950000 61.180000 70.150000 61.380000 ;
        RECT 69.950000 61.590000 70.150000 61.790000 ;
        RECT 69.950000 62.000000 70.150000 62.200000 ;
        RECT 69.950000 62.410000 70.150000 62.610000 ;
        RECT 70.355000 58.310000 70.555000 58.510000 ;
        RECT 70.355000 58.720000 70.555000 58.920000 ;
        RECT 70.355000 59.130000 70.555000 59.330000 ;
        RECT 70.355000 59.540000 70.555000 59.740000 ;
        RECT 70.355000 59.950000 70.555000 60.150000 ;
        RECT 70.355000 60.360000 70.555000 60.560000 ;
        RECT 70.355000 60.770000 70.555000 60.970000 ;
        RECT 70.355000 61.180000 70.555000 61.380000 ;
        RECT 70.355000 61.590000 70.555000 61.790000 ;
        RECT 70.355000 62.000000 70.555000 62.200000 ;
        RECT 70.355000 62.410000 70.555000 62.610000 ;
        RECT 70.760000 58.310000 70.960000 58.510000 ;
        RECT 70.760000 58.720000 70.960000 58.920000 ;
        RECT 70.760000 59.130000 70.960000 59.330000 ;
        RECT 70.760000 59.540000 70.960000 59.740000 ;
        RECT 70.760000 59.950000 70.960000 60.150000 ;
        RECT 70.760000 60.360000 70.960000 60.560000 ;
        RECT 70.760000 60.770000 70.960000 60.970000 ;
        RECT 70.760000 61.180000 70.960000 61.380000 ;
        RECT 70.760000 61.590000 70.960000 61.790000 ;
        RECT 70.760000 62.000000 70.960000 62.200000 ;
        RECT 70.760000 62.410000 70.960000 62.610000 ;
        RECT 71.165000 58.310000 71.365000 58.510000 ;
        RECT 71.165000 58.720000 71.365000 58.920000 ;
        RECT 71.165000 59.130000 71.365000 59.330000 ;
        RECT 71.165000 59.540000 71.365000 59.740000 ;
        RECT 71.165000 59.950000 71.365000 60.150000 ;
        RECT 71.165000 60.360000 71.365000 60.560000 ;
        RECT 71.165000 60.770000 71.365000 60.970000 ;
        RECT 71.165000 61.180000 71.365000 61.380000 ;
        RECT 71.165000 61.590000 71.365000 61.790000 ;
        RECT 71.165000 62.000000 71.365000 62.200000 ;
        RECT 71.165000 62.410000 71.365000 62.610000 ;
        RECT 71.570000 58.310000 71.770000 58.510000 ;
        RECT 71.570000 58.720000 71.770000 58.920000 ;
        RECT 71.570000 59.130000 71.770000 59.330000 ;
        RECT 71.570000 59.540000 71.770000 59.740000 ;
        RECT 71.570000 59.950000 71.770000 60.150000 ;
        RECT 71.570000 60.360000 71.770000 60.560000 ;
        RECT 71.570000 60.770000 71.770000 60.970000 ;
        RECT 71.570000 61.180000 71.770000 61.380000 ;
        RECT 71.570000 61.590000 71.770000 61.790000 ;
        RECT 71.570000 62.000000 71.770000 62.200000 ;
        RECT 71.570000 62.410000 71.770000 62.610000 ;
        RECT 71.975000 58.310000 72.175000 58.510000 ;
        RECT 71.975000 58.720000 72.175000 58.920000 ;
        RECT 71.975000 59.130000 72.175000 59.330000 ;
        RECT 71.975000 59.540000 72.175000 59.740000 ;
        RECT 71.975000 59.950000 72.175000 60.150000 ;
        RECT 71.975000 60.360000 72.175000 60.560000 ;
        RECT 71.975000 60.770000 72.175000 60.970000 ;
        RECT 71.975000 61.180000 72.175000 61.380000 ;
        RECT 71.975000 61.590000 72.175000 61.790000 ;
        RECT 71.975000 62.000000 72.175000 62.200000 ;
        RECT 71.975000 62.410000 72.175000 62.610000 ;
        RECT 72.380000 58.310000 72.580000 58.510000 ;
        RECT 72.380000 58.720000 72.580000 58.920000 ;
        RECT 72.380000 59.130000 72.580000 59.330000 ;
        RECT 72.380000 59.540000 72.580000 59.740000 ;
        RECT 72.380000 59.950000 72.580000 60.150000 ;
        RECT 72.380000 60.360000 72.580000 60.560000 ;
        RECT 72.380000 60.770000 72.580000 60.970000 ;
        RECT 72.380000 61.180000 72.580000 61.380000 ;
        RECT 72.380000 61.590000 72.580000 61.790000 ;
        RECT 72.380000 62.000000 72.580000 62.200000 ;
        RECT 72.380000 62.410000 72.580000 62.610000 ;
        RECT 72.785000 58.310000 72.985000 58.510000 ;
        RECT 72.785000 58.720000 72.985000 58.920000 ;
        RECT 72.785000 59.130000 72.985000 59.330000 ;
        RECT 72.785000 59.540000 72.985000 59.740000 ;
        RECT 72.785000 59.950000 72.985000 60.150000 ;
        RECT 72.785000 60.360000 72.985000 60.560000 ;
        RECT 72.785000 60.770000 72.985000 60.970000 ;
        RECT 72.785000 61.180000 72.985000 61.380000 ;
        RECT 72.785000 61.590000 72.985000 61.790000 ;
        RECT 72.785000 62.000000 72.985000 62.200000 ;
        RECT 72.785000 62.410000 72.985000 62.610000 ;
        RECT 73.190000 58.310000 73.390000 58.510000 ;
        RECT 73.190000 58.720000 73.390000 58.920000 ;
        RECT 73.190000 59.130000 73.390000 59.330000 ;
        RECT 73.190000 59.540000 73.390000 59.740000 ;
        RECT 73.190000 59.950000 73.390000 60.150000 ;
        RECT 73.190000 60.360000 73.390000 60.560000 ;
        RECT 73.190000 60.770000 73.390000 60.970000 ;
        RECT 73.190000 61.180000 73.390000 61.380000 ;
        RECT 73.190000 61.590000 73.390000 61.790000 ;
        RECT 73.190000 62.000000 73.390000 62.200000 ;
        RECT 73.190000 62.410000 73.390000 62.610000 ;
        RECT 73.595000 58.310000 73.795000 58.510000 ;
        RECT 73.595000 58.720000 73.795000 58.920000 ;
        RECT 73.595000 59.130000 73.795000 59.330000 ;
        RECT 73.595000 59.540000 73.795000 59.740000 ;
        RECT 73.595000 59.950000 73.795000 60.150000 ;
        RECT 73.595000 60.360000 73.795000 60.560000 ;
        RECT 73.595000 60.770000 73.795000 60.970000 ;
        RECT 73.595000 61.180000 73.795000 61.380000 ;
        RECT 73.595000 61.590000 73.795000 61.790000 ;
        RECT 73.595000 62.000000 73.795000 62.200000 ;
        RECT 73.595000 62.410000 73.795000 62.610000 ;
        RECT 74.000000 58.310000 74.200000 58.510000 ;
        RECT 74.000000 58.720000 74.200000 58.920000 ;
        RECT 74.000000 59.130000 74.200000 59.330000 ;
        RECT 74.000000 59.540000 74.200000 59.740000 ;
        RECT 74.000000 59.950000 74.200000 60.150000 ;
        RECT 74.000000 60.360000 74.200000 60.560000 ;
        RECT 74.000000 60.770000 74.200000 60.970000 ;
        RECT 74.000000 61.180000 74.200000 61.380000 ;
        RECT 74.000000 61.590000 74.200000 61.790000 ;
        RECT 74.000000 62.000000 74.200000 62.200000 ;
        RECT 74.000000 62.410000 74.200000 62.610000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000 75.000000  25.440000 ;
      RECT  0.000000  30.880000 75.000000  57.840000 ;
      RECT  0.000000  63.080000 75.000000 172.755000 ;
      RECT 13.900000  63.080000 61.100000 195.175000 ;
      RECT 13.900000  63.080000 75.000000 172.920000 ;
      RECT 13.900000 172.755000 75.000000 172.920000 ;
      RECT 13.900000 172.920000 61.100000 195.145000 ;
      RECT 13.900000 195.145000 61.085000 195.160000 ;
      RECT 13.900000 195.145000 61.085000 195.160000 ;
      RECT 13.900000 195.160000 61.070000 195.175000 ;
      RECT 13.900000 195.160000 61.070000 195.175000 ;
      RECT 14.050000 195.175000 60.920000 195.325000 ;
      RECT 14.050000 195.175000 60.920000 195.325000 ;
      RECT 14.200000 195.325000 60.770000 195.475000 ;
      RECT 14.200000 195.325000 60.770000 195.475000 ;
      RECT 14.350000 195.475000 60.620000 195.625000 ;
      RECT 14.350000 195.475000 60.620000 195.625000 ;
      RECT 14.500000 195.625000 60.470000 195.775000 ;
      RECT 14.500000 195.625000 60.470000 195.775000 ;
      RECT 14.650000 195.775000 60.320000 195.925000 ;
      RECT 14.650000 195.775000 60.320000 195.925000 ;
      RECT 14.800000 195.925000 60.170000 196.075000 ;
      RECT 14.800000 195.925000 60.170000 196.075000 ;
      RECT 14.950000 196.075000 60.020000 196.225000 ;
      RECT 14.950000 196.075000 60.020000 196.225000 ;
      RECT 15.100000 196.225000 59.870000 196.375000 ;
      RECT 15.100000 196.225000 59.870000 196.375000 ;
      RECT 15.250000 196.375000 59.720000 196.525000 ;
      RECT 15.250000 196.375000 59.720000 196.525000 ;
      RECT 15.400000 196.525000 59.570000 196.675000 ;
      RECT 15.400000 196.525000 59.570000 196.675000 ;
      RECT 15.500000 196.675000 59.470000 196.775000 ;
      RECT 15.500000 196.675000 59.470000 196.775000 ;
      RECT 24.795000   0.000000 49.990000  63.080000 ;
      RECT 24.795000   0.000000 49.990000 172.920000 ;
      RECT 24.795000  25.440000 49.990000  30.880000 ;
      RECT 24.795000  57.840000 49.990000  63.080000 ;
      RECT 74.690000  25.440000 75.000000  30.880000 ;
      RECT 74.690000  57.840000 75.000000  63.080000 ;
      RECT 74.690000 172.920000 75.000000 200.000000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000   0.000000 73.330000  25.435000 ;
      RECT  1.670000   0.000000 73.330000  25.435000 ;
      RECT  1.670000   0.000000 73.330000  25.435000 ;
      RECT  1.670000  19.385000 73.330000  25.435000 ;
      RECT  1.670000  30.885000 73.330000  57.835000 ;
      RECT  1.670000  30.885000 73.330000  57.835000 ;
      RECT  1.670000  30.885000 73.330000  57.835000 ;
      RECT  1.670000  30.885000 73.330000  57.835000 ;
      RECT  1.670000  30.885000 73.330000  57.835000 ;
      RECT  1.670000  63.085000 73.330000  95.400000 ;
      RECT  1.670000  63.085000 73.330000 175.530000 ;
      RECT  1.670000  63.085000 73.330000 175.530000 ;
      RECT  1.670000  63.085000 73.330000 175.530000 ;
      RECT  1.670000 175.385000 73.330000 175.530000 ;
      RECT 13.875000  63.085000 61.105000 195.830000 ;
      RECT 13.875000 175.530000 61.105000 195.830000 ;
      RECT 14.655000  63.085000 60.280000 196.770000 ;
      RECT 14.655000 195.830000 60.280000 196.770000 ;
      RECT 24.770000   0.000000 50.015000  63.085000 ;
      RECT 24.770000   0.000000 50.015000 196.770000 ;
      RECT 24.770000  25.435000 50.015000  30.885000 ;
      RECT 24.770000  57.835000 50.015000  63.085000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT 0.000000   0.000000 75.000000   1.335000 ;
      RECT 0.000000  95.785000 75.000000 174.985000 ;
      RECT 1.765000  14.235000 73.235000  19.085000 ;
      RECT 2.070000   1.335000 72.930000  14.235000 ;
      RECT 2.070000  19.085000 72.930000  95.785000 ;
      RECT 2.070000 174.985000 72.930000 200.000000 ;
  END
END sky130_fd_io__overlay_vssio_hvc


MACRO sky130_fd_io__top_power_hvc_wpad
  CLASS PAD ;
  ORIGIN  0.000000  0.000000 ;
  FOREIGN sky130_fd_io__top_power_hvc_wpad  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN P_PAD
    ANTENNAPARTIALMETALSIDEAREA  284.1730 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT  4.800000 104.230000 70.200000 166.570000 ;
        RECT  4.930000 104.100000 70.070000 104.230000 ;
        RECT  5.200000 166.570000 69.800000 166.970000 ;
        RECT  5.330000 103.700000 69.670000 104.100000 ;
        RECT  5.600000 166.970000 69.400000 167.370000 ;
        RECT  5.730000 103.300000 69.270000 103.700000 ;
        RECT  6.000000 167.370000 69.000000 167.770000 ;
        RECT  6.130000 102.900000 68.870000 103.300000 ;
        RECT  6.400000 167.770000 68.600000 168.170000 ;
        RECT  6.530000 102.500000 68.470000 102.900000 ;
        RECT  6.800000 168.170000 68.200000 168.570000 ;
        RECT  6.930000 102.100000 68.070000 102.500000 ;
        RECT  7.200000 168.570000 67.800000 168.970000 ;
        RECT  7.330000 101.700000 67.670000 102.100000 ;
        RECT  7.600000 168.970000 67.400000 169.370000 ;
        RECT  7.730000 101.300000 67.270000 101.700000 ;
        RECT  8.000000 169.370000 67.000000 169.770000 ;
        RECT  8.130000 100.900000 66.870000 101.300000 ;
        RECT  8.400000 169.770000 66.600000 170.170000 ;
        RECT  8.530000 100.500000 66.470000 100.900000 ;
        RECT  8.800000 170.170000 66.200000 170.570000 ;
        RECT  8.930000 100.100000 66.070000 100.500000 ;
        RECT  9.200000 170.570000 65.800000 170.970000 ;
        RECT  9.330000  99.700000 65.670000 100.100000 ;
        RECT  9.600000 170.970000 65.400000 171.370000 ;
        RECT  9.730000  99.300000 65.270000  99.700000 ;
        RECT 10.000000 171.370000 65.000000 171.770000 ;
        RECT 10.130000  98.900000 64.870000  99.300000 ;
        RECT 10.400000 171.770000 64.600000 172.170000 ;
        RECT 10.530000  98.500000 64.470000  98.900000 ;
        RECT 10.800000 172.170000 64.200000 172.570000 ;
        RECT 10.930000  98.100000 64.070000  98.500000 ;
        RECT 11.200000 172.570000 63.800000 172.970000 ;
        RECT 11.330000  97.700000 63.670000  98.100000 ;
        RECT 11.330000 172.970000 63.670000 173.100000 ;
    END
  END P_PAD
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 15.620000 185.295000 74.290000 190.015000 ;
        RECT 16.805000  47.455000 74.290000  54.765000 ;
        RECT 16.805000 139.455000 74.290000 146.710000 ;
        RECT 16.805000 162.455000 74.290000 171.155000 ;
        RECT 16.875000 146.710000 74.290000 146.780000 ;
        RECT 16.945000 146.780000 74.290000 146.850000 ;
        RECT 17.015000 146.850000 74.290000 146.920000 ;
        RECT 17.085000 146.920000 74.290000 146.990000 ;
        RECT 17.155000 146.990000 74.290000 147.060000 ;
        RECT 17.225000 147.060000 74.290000 147.130000 ;
        RECT 17.295000 147.130000 74.290000 147.200000 ;
        RECT 17.365000 147.200000 74.290000 147.270000 ;
        RECT 17.435000 147.270000 74.290000 147.340000 ;
        RECT 17.505000 147.340000 74.290000 147.410000 ;
        RECT 17.530000  54.765000 74.290000  54.835000 ;
        RECT 17.575000 147.410000 74.290000 147.480000 ;
        RECT 17.600000  54.835000 74.290000  54.905000 ;
        RECT 17.645000 147.480000 74.290000 147.550000 ;
        RECT 17.670000  54.905000 74.290000  54.975000 ;
        RECT 17.715000 147.550000 74.290000 147.620000 ;
        RECT 17.740000  54.975000 74.290000  55.045000 ;
        RECT 17.785000 147.620000 74.290000 147.690000 ;
        RECT 17.810000  55.045000 74.290000  55.115000 ;
        RECT 17.855000 147.690000 74.290000 147.760000 ;
        RECT 17.880000  55.115000 74.290000  55.185000 ;
        RECT 17.925000 147.760000 74.290000 147.830000 ;
        RECT 17.950000  55.185000 74.290000  55.255000 ;
        RECT 17.995000 147.830000 74.290000 147.900000 ;
        RECT 18.020000  55.255000 74.290000  55.325000 ;
        RECT 18.065000 147.900000 74.290000 147.970000 ;
        RECT 18.090000  55.325000 74.290000  55.395000 ;
        RECT 18.135000 147.970000 74.290000 148.040000 ;
        RECT 18.160000  55.395000 74.290000  55.465000 ;
        RECT 18.205000 148.040000 74.290000 148.110000 ;
        RECT 18.230000  55.465000 74.290000  55.535000 ;
        RECT 18.250000 148.110000 74.290000 148.155000 ;
        RECT 18.300000  55.535000 74.290000  55.605000 ;
        RECT 18.370000  55.605000 74.290000  55.675000 ;
        RECT 18.410000  74.155000 74.290000  74.415000 ;
        RECT 18.440000  55.675000 74.290000  55.745000 ;
        RECT 18.510000  55.745000 74.290000  55.815000 ;
        RECT 18.580000  55.815000 74.290000  55.885000 ;
        RECT 18.650000  55.885000 74.290000  55.955000 ;
        RECT 18.720000  55.955000 74.290000  56.025000 ;
        RECT 18.790000  56.025000 74.290000  56.095000 ;
        RECT 18.850000  56.095000 74.290000  56.155000 ;
        RECT 23.690000  74.415000 74.290000  74.485000 ;
        RECT 23.700000  74.105000 74.290000  74.155000 ;
        RECT 23.760000  74.485000 74.290000  74.555000 ;
        RECT 23.770000  74.035000 74.290000  74.105000 ;
        RECT 23.830000  74.555000 74.290000  74.625000 ;
        RECT 23.840000  73.965000 74.290000  74.035000 ;
        RECT 23.900000  74.625000 74.290000  74.695000 ;
        RECT 23.910000  73.895000 74.290000  73.965000 ;
        RECT 23.970000  74.695000 74.290000  74.765000 ;
        RECT 23.980000  73.825000 74.290000  73.895000 ;
        RECT 24.040000  74.765000 74.290000  74.835000 ;
        RECT 24.050000  73.755000 74.290000  73.825000 ;
        RECT 24.110000  74.835000 74.290000  74.905000 ;
        RECT 24.120000  73.685000 74.290000  73.755000 ;
        RECT 24.180000  74.905000 74.290000  74.975000 ;
        RECT 24.190000  73.615000 74.290000  73.685000 ;
        RECT 24.250000  74.975000 74.290000  75.045000 ;
        RECT 24.260000  73.545000 74.290000  73.615000 ;
        RECT 24.320000  75.045000 74.290000  75.115000 ;
        RECT 24.330000  73.475000 74.290000  73.545000 ;
        RECT 24.390000  75.115000 74.290000  75.185000 ;
        RECT 24.400000  73.405000 74.290000  73.475000 ;
        RECT 24.460000  75.185000 74.290000  75.255000 ;
        RECT 24.470000  73.335000 74.290000  73.405000 ;
        RECT 24.530000  75.255000 74.290000  75.325000 ;
        RECT 24.540000  73.265000 74.290000  73.335000 ;
        RECT 24.600000  75.325000 74.290000  75.395000 ;
        RECT 24.610000  73.195000 74.290000  73.265000 ;
        RECT 24.670000  75.395000 74.290000  75.465000 ;
        RECT 24.680000  73.125000 74.290000  73.195000 ;
        RECT 24.740000  75.465000 74.290000  75.535000 ;
        RECT 24.750000  73.055000 74.290000  73.125000 ;
        RECT 24.810000  75.535000 74.290000  75.605000 ;
        RECT 24.820000  70.455000 74.290000  72.985000 ;
        RECT 24.820000  72.985000 74.290000  73.055000 ;
        RECT 24.820000  75.605000 74.290000  75.615000 ;
        RECT 24.820000  75.615000 74.290000  79.155000 ;
        RECT 24.820000  93.455000 74.290000 102.155000 ;
        RECT 24.820000 116.455000 74.290000 125.155000 ;
        RECT 37.890000  12.295000 74.290000  25.660000 ;
        RECT 46.750000  12.265000 74.290000  12.295000 ;
        RECT 46.820000  12.195000 74.290000  12.265000 ;
        RECT 46.890000  12.125000 74.290000  12.195000 ;
        RECT 46.960000  12.055000 74.290000  12.125000 ;
        RECT 47.030000  11.985000 74.290000  12.055000 ;
        RECT 47.100000  11.915000 74.290000  11.985000 ;
        RECT 47.170000  11.845000 74.290000  11.915000 ;
        RECT 47.240000  11.775000 74.290000  11.845000 ;
        RECT 47.310000  11.705000 74.290000  11.775000 ;
        RECT 47.380000  11.635000 74.290000  11.705000 ;
        RECT 47.450000  11.565000 74.290000  11.635000 ;
        RECT 47.520000  11.495000 74.290000  11.565000 ;
        RECT 47.590000  11.425000 74.290000  11.495000 ;
        RECT 47.660000  11.355000 74.290000  11.425000 ;
        RECT 47.730000  11.285000 74.290000  11.355000 ;
        RECT 47.800000  11.215000 74.290000  11.285000 ;
        RECT 47.870000  11.145000 74.290000  11.215000 ;
        RECT 47.940000  11.075000 74.290000  11.145000 ;
        RECT 48.010000  11.005000 74.290000  11.075000 ;
        RECT 48.080000  10.935000 74.290000  11.005000 ;
        RECT 48.150000  10.865000 74.290000  10.935000 ;
        RECT 48.220000  10.795000 74.290000  10.865000 ;
        RECT 48.290000  10.725000 74.290000  10.795000 ;
        RECT 48.360000  10.655000 74.290000  10.725000 ;
        RECT 48.430000  10.585000 74.290000  10.655000 ;
        RECT 48.500000  10.515000 74.290000  10.585000 ;
        RECT 48.570000  10.445000 74.290000  10.515000 ;
        RECT 48.640000  10.375000 74.290000  10.445000 ;
        RECT 48.710000  10.305000 74.290000  10.375000 ;
        RECT 48.780000  10.235000 74.290000  10.305000 ;
        RECT 48.850000  10.165000 74.290000  10.235000 ;
        RECT 48.920000  10.095000 74.290000  10.165000 ;
        RECT 48.990000  10.025000 74.290000  10.095000 ;
        RECT 49.060000   9.955000 74.290000  10.025000 ;
        RECT 49.130000   9.885000 74.290000   9.955000 ;
        RECT 49.200000   9.815000 74.290000   9.885000 ;
        RECT 49.270000   9.745000 74.290000   9.815000 ;
        RECT 49.340000   9.675000 74.290000   9.745000 ;
        RECT 49.410000   9.605000 74.290000   9.675000 ;
        RECT 49.480000   9.535000 74.290000   9.605000 ;
        RECT 49.550000   9.465000 74.290000   9.535000 ;
        RECT 49.620000   9.395000 74.290000   9.465000 ;
        RECT 49.690000   9.325000 74.290000   9.395000 ;
        RECT 49.760000   9.255000 74.290000   9.325000 ;
        RECT 49.830000   9.185000 74.290000   9.255000 ;
        RECT 49.900000   9.115000 74.290000   9.185000 ;
        RECT 49.970000   9.045000 74.290000   9.115000 ;
        RECT 50.040000   8.975000 74.290000   9.045000 ;
        RECT 50.110000   8.905000 74.290000   8.975000 ;
        RECT 50.180000   8.835000 74.290000   8.905000 ;
        RECT 50.250000   8.765000 74.290000   8.835000 ;
        RECT 50.320000   8.695000 74.290000   8.765000 ;
        RECT 50.390000   0.000000 74.290000   8.625000 ;
        RECT 50.390000   8.625000 74.290000   8.695000 ;
        RECT 55.885000  25.660000 74.290000  25.730000 ;
        RECT 55.955000  25.730000 74.290000  25.800000 ;
        RECT 56.025000  25.800000 74.290000  25.870000 ;
        RECT 56.095000  25.870000 74.290000  25.940000 ;
        RECT 56.165000  25.940000 74.290000  26.010000 ;
        RECT 56.235000  26.010000 74.290000  26.080000 ;
        RECT 56.305000  26.080000 74.290000  26.150000 ;
        RECT 56.375000  26.150000 74.290000  26.220000 ;
        RECT 56.445000  26.220000 74.290000  26.290000 ;
        RECT 56.515000  26.290000 74.290000  26.360000 ;
        RECT 56.585000  26.360000 74.290000  26.430000 ;
        RECT 56.655000  26.430000 74.290000  26.500000 ;
        RECT 56.725000  26.500000 74.290000  26.570000 ;
        RECT 56.795000  26.570000 74.290000  26.640000 ;
        RECT 56.865000  26.640000 74.290000  26.710000 ;
        RECT 56.935000  26.710000 74.290000  26.780000 ;
        RECT 57.005000  26.780000 74.290000  26.850000 ;
        RECT 57.075000  26.850000 74.290000  26.920000 ;
        RECT 57.145000  26.920000 74.290000  26.990000 ;
        RECT 57.215000  26.990000 74.290000  27.060000 ;
        RECT 57.285000  27.060000 74.290000  27.130000 ;
        RECT 57.355000  27.130000 74.290000  27.200000 ;
        RECT 57.425000  27.200000 74.290000  27.270000 ;
        RECT 57.495000  27.270000 74.290000  27.340000 ;
        RECT 57.540000  47.390000 74.290000  47.455000 ;
        RECT 57.540000  70.420000 74.290000  70.455000 ;
        RECT 57.540000 116.390000 74.290000 116.455000 ;
        RECT 57.540000 139.425000 74.290000 139.455000 ;
        RECT 57.540000 162.440000 74.290000 162.455000 ;
        RECT 57.555000 148.155000 74.290000 148.225000 ;
        RECT 57.565000  27.340000 74.290000  27.410000 ;
        RECT 57.595000  56.155000 74.290000  56.225000 ;
        RECT 57.610000  47.320000 74.290000  47.390000 ;
        RECT 57.610000  70.350000 74.290000  70.420000 ;
        RECT 57.610000  93.410000 74.290000  93.455000 ;
        RECT 57.610000 116.320000 74.290000 116.390000 ;
        RECT 57.610000 139.355000 74.290000 139.425000 ;
        RECT 57.610000 162.370000 74.290000 162.440000 ;
        RECT 57.625000  79.155000 74.290000  79.225000 ;
        RECT 57.625000 102.155000 74.290000 102.225000 ;
        RECT 57.625000 125.155000 74.290000 125.225000 ;
        RECT 57.625000 148.225000 74.290000 148.295000 ;
        RECT 57.635000  27.410000 74.290000  27.480000 ;
        RECT 57.635000 171.155000 74.290000 171.225000 ;
        RECT 57.665000  56.225000 74.290000  56.295000 ;
        RECT 57.680000  47.250000 74.290000  47.320000 ;
        RECT 57.680000  70.280000 74.290000  70.350000 ;
        RECT 57.680000  93.340000 74.290000  93.410000 ;
        RECT 57.680000 116.250000 74.290000 116.320000 ;
        RECT 57.680000 139.285000 74.290000 139.355000 ;
        RECT 57.680000 162.300000 74.290000 162.370000 ;
        RECT 57.695000  79.225000 74.290000  79.295000 ;
        RECT 57.695000 102.225000 74.290000 102.295000 ;
        RECT 57.695000 125.225000 74.290000 125.295000 ;
        RECT 57.695000 148.295000 74.290000 148.365000 ;
        RECT 57.705000  27.480000 74.290000  27.550000 ;
        RECT 57.705000 171.225000 74.290000 171.295000 ;
        RECT 57.735000  56.295000 74.290000  56.365000 ;
        RECT 57.750000  47.180000 74.290000  47.250000 ;
        RECT 57.750000  70.210000 74.290000  70.280000 ;
        RECT 57.750000  93.270000 74.290000  93.340000 ;
        RECT 57.750000 116.180000 74.290000 116.250000 ;
        RECT 57.750000 139.215000 74.290000 139.285000 ;
        RECT 57.750000 162.230000 74.290000 162.300000 ;
        RECT 57.765000  79.295000 74.290000  79.365000 ;
        RECT 57.765000 102.295000 74.290000 102.365000 ;
        RECT 57.765000 125.295000 74.290000 125.365000 ;
        RECT 57.765000 148.365000 74.290000 148.435000 ;
        RECT 57.775000  27.550000 74.290000  27.620000 ;
        RECT 57.775000 171.295000 74.290000 171.365000 ;
        RECT 57.805000  56.365000 74.290000  56.435000 ;
        RECT 57.820000  47.110000 74.290000  47.180000 ;
        RECT 57.820000  70.140000 74.290000  70.210000 ;
        RECT 57.820000  93.200000 74.290000  93.270000 ;
        RECT 57.820000 116.110000 74.290000 116.180000 ;
        RECT 57.820000 139.145000 74.290000 139.215000 ;
        RECT 57.820000 162.160000 74.290000 162.230000 ;
        RECT 57.835000  79.365000 74.290000  79.435000 ;
        RECT 57.835000 102.365000 74.290000 102.435000 ;
        RECT 57.835000 125.365000 74.290000 125.435000 ;
        RECT 57.835000 148.435000 74.290000 148.505000 ;
        RECT 57.845000  27.620000 74.290000  27.690000 ;
        RECT 57.845000 171.365000 74.290000 171.435000 ;
        RECT 57.875000  56.435000 74.290000  56.505000 ;
        RECT 57.890000  47.040000 74.290000  47.110000 ;
        RECT 57.890000  70.070000 74.290000  70.140000 ;
        RECT 57.890000  93.130000 74.290000  93.200000 ;
        RECT 57.890000 116.040000 74.290000 116.110000 ;
        RECT 57.890000 139.075000 74.290000 139.145000 ;
        RECT 57.890000 162.090000 74.290000 162.160000 ;
        RECT 57.905000  79.435000 74.290000  79.505000 ;
        RECT 57.905000 102.435000 74.290000 102.505000 ;
        RECT 57.905000 125.435000 74.290000 125.505000 ;
        RECT 57.905000 148.505000 74.290000 148.575000 ;
        RECT 57.915000  27.690000 74.290000  27.760000 ;
        RECT 57.915000 171.435000 74.290000 171.505000 ;
        RECT 57.945000  56.505000 74.290000  56.575000 ;
        RECT 57.960000  46.970000 74.290000  47.040000 ;
        RECT 57.960000  70.000000 74.290000  70.070000 ;
        RECT 57.960000  93.060000 74.290000  93.130000 ;
        RECT 57.960000 115.970000 74.290000 116.040000 ;
        RECT 57.960000 139.005000 74.290000 139.075000 ;
        RECT 57.960000 162.020000 74.290000 162.090000 ;
        RECT 57.975000  79.505000 74.290000  79.575000 ;
        RECT 57.975000 102.505000 74.290000 102.575000 ;
        RECT 57.975000 125.505000 74.290000 125.575000 ;
        RECT 57.975000 148.575000 74.290000 148.645000 ;
        RECT 57.985000  27.760000 74.290000  27.830000 ;
        RECT 57.985000 171.505000 74.290000 171.575000 ;
        RECT 58.015000  56.575000 74.290000  56.645000 ;
        RECT 58.030000  46.900000 74.290000  46.970000 ;
        RECT 58.030000  69.930000 74.290000  70.000000 ;
        RECT 58.030000  92.990000 74.290000  93.060000 ;
        RECT 58.030000 115.900000 74.290000 115.970000 ;
        RECT 58.030000 138.935000 74.290000 139.005000 ;
        RECT 58.030000 161.950000 74.290000 162.020000 ;
        RECT 58.045000  79.575000 74.290000  79.645000 ;
        RECT 58.045000 102.575000 74.290000 102.645000 ;
        RECT 58.045000 125.575000 74.290000 125.645000 ;
        RECT 58.045000 148.645000 74.290000 148.715000 ;
        RECT 58.055000  27.830000 74.290000  27.900000 ;
        RECT 58.055000 171.575000 74.290000 171.645000 ;
        RECT 58.085000  56.645000 74.290000  56.715000 ;
        RECT 58.100000  46.830000 74.290000  46.900000 ;
        RECT 58.100000  69.860000 74.290000  69.930000 ;
        RECT 58.100000  92.920000 74.290000  92.990000 ;
        RECT 58.100000 115.830000 74.290000 115.900000 ;
        RECT 58.100000 138.865000 74.290000 138.935000 ;
        RECT 58.100000 161.880000 74.290000 161.950000 ;
        RECT 58.115000  79.645000 74.290000  79.715000 ;
        RECT 58.115000 102.645000 74.290000 102.715000 ;
        RECT 58.115000 125.645000 74.290000 125.715000 ;
        RECT 58.115000 148.715000 74.290000 148.785000 ;
        RECT 58.125000  27.900000 74.290000  27.970000 ;
        RECT 58.125000 171.645000 74.290000 171.715000 ;
        RECT 58.155000  56.715000 74.290000  56.785000 ;
        RECT 58.170000  46.760000 74.290000  46.830000 ;
        RECT 58.170000  69.790000 74.290000  69.860000 ;
        RECT 58.170000  92.850000 74.290000  92.920000 ;
        RECT 58.170000 115.760000 74.290000 115.830000 ;
        RECT 58.170000 138.795000 74.290000 138.865000 ;
        RECT 58.170000 161.810000 74.290000 161.880000 ;
        RECT 58.185000  79.715000 74.290000  79.785000 ;
        RECT 58.185000 102.715000 74.290000 102.785000 ;
        RECT 58.185000 125.715000 74.290000 125.785000 ;
        RECT 58.185000 148.785000 74.290000 148.855000 ;
        RECT 58.195000  27.970000 74.290000  28.040000 ;
        RECT 58.195000 171.715000 74.290000 171.785000 ;
        RECT 58.225000  56.785000 74.290000  56.855000 ;
        RECT 58.240000  46.690000 74.290000  46.760000 ;
        RECT 58.240000  69.720000 74.290000  69.790000 ;
        RECT 58.240000  92.780000 74.290000  92.850000 ;
        RECT 58.240000 115.690000 74.290000 115.760000 ;
        RECT 58.240000 138.725000 74.290000 138.795000 ;
        RECT 58.240000 161.740000 74.290000 161.810000 ;
        RECT 58.255000  79.785000 74.290000  79.855000 ;
        RECT 58.255000 102.785000 74.290000 102.855000 ;
        RECT 58.255000 125.785000 74.290000 125.855000 ;
        RECT 58.255000 148.855000 74.290000 148.925000 ;
        RECT 58.265000  28.040000 74.290000  28.110000 ;
        RECT 58.265000 171.785000 74.290000 171.855000 ;
        RECT 58.295000  56.855000 74.290000  56.925000 ;
        RECT 58.310000  46.620000 74.290000  46.690000 ;
        RECT 58.310000  69.650000 74.290000  69.720000 ;
        RECT 58.310000  92.710000 74.290000  92.780000 ;
        RECT 58.310000 115.620000 74.290000 115.690000 ;
        RECT 58.310000 138.655000 74.290000 138.725000 ;
        RECT 58.310000 161.670000 74.290000 161.740000 ;
        RECT 58.325000  79.855000 74.290000  79.925000 ;
        RECT 58.325000 102.855000 74.290000 102.925000 ;
        RECT 58.325000 125.855000 74.290000 125.925000 ;
        RECT 58.325000 148.925000 74.290000 148.995000 ;
        RECT 58.335000  28.110000 74.290000  28.180000 ;
        RECT 58.335000 171.855000 74.290000 171.925000 ;
        RECT 58.365000  56.925000 74.290000  56.995000 ;
        RECT 58.380000  46.550000 74.290000  46.620000 ;
        RECT 58.380000  69.580000 74.290000  69.650000 ;
        RECT 58.380000  92.640000 74.290000  92.710000 ;
        RECT 58.380000 115.550000 74.290000 115.620000 ;
        RECT 58.380000 138.585000 74.290000 138.655000 ;
        RECT 58.380000 161.600000 74.290000 161.670000 ;
        RECT 58.395000  79.925000 74.290000  79.995000 ;
        RECT 58.395000 102.925000 74.290000 102.995000 ;
        RECT 58.395000 125.925000 74.290000 125.995000 ;
        RECT 58.395000 148.995000 74.290000 149.065000 ;
        RECT 58.405000  28.180000 74.290000  28.250000 ;
        RECT 58.405000 171.925000 74.290000 171.995000 ;
        RECT 58.435000  56.995000 74.290000  57.065000 ;
        RECT 58.450000  46.480000 74.290000  46.550000 ;
        RECT 58.450000  69.510000 74.290000  69.580000 ;
        RECT 58.450000  92.570000 74.290000  92.640000 ;
        RECT 58.450000 115.480000 74.290000 115.550000 ;
        RECT 58.450000 138.515000 74.290000 138.585000 ;
        RECT 58.450000 161.530000 74.290000 161.600000 ;
        RECT 58.465000  79.995000 74.290000  80.065000 ;
        RECT 58.465000 102.995000 74.290000 103.065000 ;
        RECT 58.465000 125.995000 74.290000 126.065000 ;
        RECT 58.465000 149.065000 74.290000 149.135000 ;
        RECT 58.475000  28.250000 74.290000  28.320000 ;
        RECT 58.475000 171.995000 74.290000 172.065000 ;
        RECT 58.505000  57.065000 74.290000  57.135000 ;
        RECT 58.520000  46.410000 74.290000  46.480000 ;
        RECT 58.520000  69.440000 74.290000  69.510000 ;
        RECT 58.520000  92.500000 74.290000  92.570000 ;
        RECT 58.520000 115.410000 74.290000 115.480000 ;
        RECT 58.520000 138.445000 74.290000 138.515000 ;
        RECT 58.520000 161.460000 74.290000 161.530000 ;
        RECT 58.535000  80.065000 74.290000  80.135000 ;
        RECT 58.535000 103.065000 74.290000 103.135000 ;
        RECT 58.535000 126.065000 74.290000 126.135000 ;
        RECT 58.535000 149.135000 74.290000 149.205000 ;
        RECT 58.545000  28.320000 74.290000  28.390000 ;
        RECT 58.545000 172.065000 74.290000 172.135000 ;
        RECT 58.575000  57.135000 74.290000  57.205000 ;
        RECT 58.590000  46.340000 74.290000  46.410000 ;
        RECT 58.590000  69.370000 74.290000  69.440000 ;
        RECT 58.590000  92.430000 74.290000  92.500000 ;
        RECT 58.590000 115.340000 74.290000 115.410000 ;
        RECT 58.590000 138.375000 74.290000 138.445000 ;
        RECT 58.590000 161.390000 74.290000 161.460000 ;
        RECT 58.605000  80.135000 74.290000  80.205000 ;
        RECT 58.605000 103.135000 74.290000 103.205000 ;
        RECT 58.605000 126.135000 74.290000 126.205000 ;
        RECT 58.605000 149.205000 74.290000 149.275000 ;
        RECT 58.615000  28.390000 74.290000  28.460000 ;
        RECT 58.615000 172.135000 74.290000 172.205000 ;
        RECT 58.645000  57.205000 74.290000  57.275000 ;
        RECT 58.660000  46.270000 74.290000  46.340000 ;
        RECT 58.660000  69.300000 74.290000  69.370000 ;
        RECT 58.660000  92.360000 74.290000  92.430000 ;
        RECT 58.660000 115.270000 74.290000 115.340000 ;
        RECT 58.660000 138.305000 74.290000 138.375000 ;
        RECT 58.660000 161.320000 74.290000 161.390000 ;
        RECT 58.675000  80.205000 74.290000  80.275000 ;
        RECT 58.675000 103.205000 74.290000 103.275000 ;
        RECT 58.675000 126.205000 74.290000 126.275000 ;
        RECT 58.675000 149.275000 74.290000 149.345000 ;
        RECT 58.685000  28.460000 74.290000  28.530000 ;
        RECT 58.685000 172.205000 74.290000 172.275000 ;
        RECT 58.715000  57.275000 74.290000  57.345000 ;
        RECT 58.730000  46.200000 74.290000  46.270000 ;
        RECT 58.730000  69.230000 74.290000  69.300000 ;
        RECT 58.730000  92.290000 74.290000  92.360000 ;
        RECT 58.730000 115.200000 74.290000 115.270000 ;
        RECT 58.730000 138.235000 74.290000 138.305000 ;
        RECT 58.730000 161.250000 74.290000 161.320000 ;
        RECT 58.730000 185.260000 74.290000 185.295000 ;
        RECT 58.745000  80.275000 74.290000  80.345000 ;
        RECT 58.745000 103.275000 74.290000 103.345000 ;
        RECT 58.745000 126.275000 74.290000 126.345000 ;
        RECT 58.745000 149.345000 74.290000 149.415000 ;
        RECT 58.755000  28.530000 74.290000  28.600000 ;
        RECT 58.755000 172.275000 74.290000 172.345000 ;
        RECT 58.785000  57.345000 74.290000  57.415000 ;
        RECT 58.800000  46.130000 74.290000  46.200000 ;
        RECT 58.800000  69.160000 74.290000  69.230000 ;
        RECT 58.800000  92.220000 74.290000  92.290000 ;
        RECT 58.800000 115.130000 74.290000 115.200000 ;
        RECT 58.800000 138.165000 74.290000 138.235000 ;
        RECT 58.800000 161.180000 74.290000 161.250000 ;
        RECT 58.800000 185.190000 74.290000 185.260000 ;
        RECT 58.815000  80.345000 74.290000  80.415000 ;
        RECT 58.815000 103.345000 74.290000 103.415000 ;
        RECT 58.815000 126.345000 74.290000 126.415000 ;
        RECT 58.815000 149.415000 74.290000 149.485000 ;
        RECT 58.825000  28.600000 74.290000  28.670000 ;
        RECT 58.825000 172.345000 74.290000 172.415000 ;
        RECT 58.855000  57.415000 74.290000  57.485000 ;
        RECT 58.870000  46.060000 74.290000  46.130000 ;
        RECT 58.870000  69.090000 74.290000  69.160000 ;
        RECT 58.870000  92.150000 74.290000  92.220000 ;
        RECT 58.870000 115.060000 74.290000 115.130000 ;
        RECT 58.870000 138.095000 74.290000 138.165000 ;
        RECT 58.870000 161.110000 74.290000 161.180000 ;
        RECT 58.870000 185.120000 74.290000 185.190000 ;
        RECT 58.885000  80.415000 74.290000  80.485000 ;
        RECT 58.885000 103.415000 74.290000 103.485000 ;
        RECT 58.885000 126.415000 74.290000 126.485000 ;
        RECT 58.885000 149.485000 74.290000 149.555000 ;
        RECT 58.895000  28.670000 74.290000  28.740000 ;
        RECT 58.895000 172.415000 74.290000 172.485000 ;
        RECT 58.925000  57.485000 74.290000  57.555000 ;
        RECT 58.940000  45.990000 74.290000  46.060000 ;
        RECT 58.940000  69.020000 74.290000  69.090000 ;
        RECT 58.940000  92.080000 74.290000  92.150000 ;
        RECT 58.940000 114.990000 74.290000 115.060000 ;
        RECT 58.940000 138.025000 74.290000 138.095000 ;
        RECT 58.940000 161.040000 74.290000 161.110000 ;
        RECT 58.940000 185.050000 74.290000 185.120000 ;
        RECT 58.955000  80.485000 74.290000  80.555000 ;
        RECT 58.955000 103.485000 74.290000 103.555000 ;
        RECT 58.955000 126.485000 74.290000 126.555000 ;
        RECT 58.955000 149.555000 74.290000 149.625000 ;
        RECT 58.965000  28.740000 74.290000  28.810000 ;
        RECT 58.965000 172.485000 74.290000 172.555000 ;
        RECT 58.995000  57.555000 74.290000  57.625000 ;
        RECT 59.010000  45.920000 74.290000  45.990000 ;
        RECT 59.010000  68.950000 74.290000  69.020000 ;
        RECT 59.010000  92.010000 74.290000  92.080000 ;
        RECT 59.010000 114.920000 74.290000 114.990000 ;
        RECT 59.010000 137.955000 74.290000 138.025000 ;
        RECT 59.010000 160.970000 74.290000 161.040000 ;
        RECT 59.010000 184.980000 74.290000 185.050000 ;
        RECT 59.025000  80.555000 74.290000  80.625000 ;
        RECT 59.025000 103.555000 74.290000 103.625000 ;
        RECT 59.025000 126.555000 74.290000 126.625000 ;
        RECT 59.025000 149.625000 74.290000 149.695000 ;
        RECT 59.035000  28.810000 74.290000  28.880000 ;
        RECT 59.035000 172.555000 74.290000 172.625000 ;
        RECT 59.065000  57.625000 74.290000  57.695000 ;
        RECT 59.080000  45.850000 74.290000  45.920000 ;
        RECT 59.080000  68.880000 74.290000  68.950000 ;
        RECT 59.080000  91.940000 74.290000  92.010000 ;
        RECT 59.080000 114.850000 74.290000 114.920000 ;
        RECT 59.080000 137.885000 74.290000 137.955000 ;
        RECT 59.080000 160.900000 74.290000 160.970000 ;
        RECT 59.080000 184.910000 74.290000 184.980000 ;
        RECT 59.095000  80.625000 74.290000  80.695000 ;
        RECT 59.095000 103.625000 74.290000 103.695000 ;
        RECT 59.095000 126.625000 74.290000 126.695000 ;
        RECT 59.095000 149.695000 74.290000 149.765000 ;
        RECT 59.105000  28.880000 74.290000  28.950000 ;
        RECT 59.105000 172.625000 74.290000 172.695000 ;
        RECT 59.135000  57.695000 74.290000  57.765000 ;
        RECT 59.150000  45.780000 74.290000  45.850000 ;
        RECT 59.150000  68.810000 74.290000  68.880000 ;
        RECT 59.150000  91.870000 74.290000  91.940000 ;
        RECT 59.150000 114.780000 74.290000 114.850000 ;
        RECT 59.150000 137.815000 74.290000 137.885000 ;
        RECT 59.150000 160.830000 74.290000 160.900000 ;
        RECT 59.150000 184.840000 74.290000 184.910000 ;
        RECT 59.165000  80.695000 74.290000  80.765000 ;
        RECT 59.165000 103.695000 74.290000 103.765000 ;
        RECT 59.165000 126.695000 74.290000 126.765000 ;
        RECT 59.165000 149.765000 74.290000 149.835000 ;
        RECT 59.175000  28.950000 74.290000  29.020000 ;
        RECT 59.175000 172.695000 74.290000 172.765000 ;
        RECT 59.205000  57.765000 74.290000  57.835000 ;
        RECT 59.220000  45.710000 74.290000  45.780000 ;
        RECT 59.220000  68.740000 74.290000  68.810000 ;
        RECT 59.220000  91.800000 74.290000  91.870000 ;
        RECT 59.220000 114.710000 74.290000 114.780000 ;
        RECT 59.220000 137.745000 74.290000 137.815000 ;
        RECT 59.220000 160.760000 74.290000 160.830000 ;
        RECT 59.220000 184.770000 74.290000 184.840000 ;
        RECT 59.235000  80.765000 74.290000  80.835000 ;
        RECT 59.235000 103.765000 74.290000 103.835000 ;
        RECT 59.235000 126.765000 74.290000 126.835000 ;
        RECT 59.235000 149.835000 74.290000 149.905000 ;
        RECT 59.245000  29.020000 74.290000  29.090000 ;
        RECT 59.245000 172.765000 74.290000 172.835000 ;
        RECT 59.275000  57.835000 74.290000  57.905000 ;
        RECT 59.290000  45.640000 74.290000  45.710000 ;
        RECT 59.290000  68.670000 74.290000  68.740000 ;
        RECT 59.290000  91.730000 74.290000  91.800000 ;
        RECT 59.290000 114.640000 74.290000 114.710000 ;
        RECT 59.290000 137.675000 74.290000 137.745000 ;
        RECT 59.290000 160.690000 74.290000 160.760000 ;
        RECT 59.290000 184.700000 74.290000 184.770000 ;
        RECT 59.305000  80.835000 74.290000  80.905000 ;
        RECT 59.305000 103.835000 74.290000 103.905000 ;
        RECT 59.305000 126.835000 74.290000 126.905000 ;
        RECT 59.305000 149.905000 74.290000 149.975000 ;
        RECT 59.315000  29.090000 74.290000  29.160000 ;
        RECT 59.315000 172.835000 74.290000 172.905000 ;
        RECT 59.345000  57.905000 74.290000  57.975000 ;
        RECT 59.360000  45.570000 74.290000  45.640000 ;
        RECT 59.360000  68.600000 74.290000  68.670000 ;
        RECT 59.360000  91.660000 74.290000  91.730000 ;
        RECT 59.360000 114.570000 74.290000 114.640000 ;
        RECT 59.360000 137.605000 74.290000 137.675000 ;
        RECT 59.360000 160.620000 74.290000 160.690000 ;
        RECT 59.360000 184.630000 74.290000 184.700000 ;
        RECT 59.375000  80.905000 74.290000  80.975000 ;
        RECT 59.375000 103.905000 74.290000 103.975000 ;
        RECT 59.375000 126.905000 74.290000 126.975000 ;
        RECT 59.375000 149.975000 74.290000 150.045000 ;
        RECT 59.385000  29.160000 74.290000  29.230000 ;
        RECT 59.385000 172.905000 74.290000 172.975000 ;
        RECT 59.415000  57.975000 74.290000  58.045000 ;
        RECT 59.430000  45.500000 74.290000  45.570000 ;
        RECT 59.430000  68.530000 74.290000  68.600000 ;
        RECT 59.430000  91.590000 74.290000  91.660000 ;
        RECT 59.430000 114.500000 74.290000 114.570000 ;
        RECT 59.430000 137.535000 74.290000 137.605000 ;
        RECT 59.430000 160.550000 74.290000 160.620000 ;
        RECT 59.430000 184.560000 74.290000 184.630000 ;
        RECT 59.445000  80.975000 74.290000  81.045000 ;
        RECT 59.445000 103.975000 74.290000 104.045000 ;
        RECT 59.445000 126.975000 74.290000 127.045000 ;
        RECT 59.445000 150.045000 74.290000 150.115000 ;
        RECT 59.455000  29.230000 74.290000  29.300000 ;
        RECT 59.455000 172.975000 74.290000 173.045000 ;
        RECT 59.485000  58.045000 74.290000  58.115000 ;
        RECT 59.500000  45.430000 74.290000  45.500000 ;
        RECT 59.500000  68.460000 74.290000  68.530000 ;
        RECT 59.500000  91.520000 74.290000  91.590000 ;
        RECT 59.500000 114.430000 74.290000 114.500000 ;
        RECT 59.500000 137.465000 74.290000 137.535000 ;
        RECT 59.500000 160.480000 74.290000 160.550000 ;
        RECT 59.500000 184.490000 74.290000 184.560000 ;
        RECT 59.515000  81.045000 74.290000  81.115000 ;
        RECT 59.515000 104.045000 74.290000 104.115000 ;
        RECT 59.515000 127.045000 74.290000 127.115000 ;
        RECT 59.515000 150.115000 74.290000 150.185000 ;
        RECT 59.525000  29.300000 74.290000  29.370000 ;
        RECT 59.525000 173.045000 74.290000 173.115000 ;
        RECT 59.555000  58.115000 74.290000  58.185000 ;
        RECT 59.570000  45.360000 74.290000  45.430000 ;
        RECT 59.570000  68.390000 74.290000  68.460000 ;
        RECT 59.570000  91.450000 74.290000  91.520000 ;
        RECT 59.570000 114.360000 74.290000 114.430000 ;
        RECT 59.570000 137.395000 74.290000 137.465000 ;
        RECT 59.570000 160.410000 74.290000 160.480000 ;
        RECT 59.570000 184.420000 74.290000 184.490000 ;
        RECT 59.585000  81.115000 74.290000  81.185000 ;
        RECT 59.585000 104.115000 74.290000 104.185000 ;
        RECT 59.585000 127.115000 74.290000 127.185000 ;
        RECT 59.585000 150.185000 74.290000 150.255000 ;
        RECT 59.595000  29.370000 74.290000  29.440000 ;
        RECT 59.595000 173.115000 74.290000 173.185000 ;
        RECT 59.625000  58.185000 74.290000  58.255000 ;
        RECT 59.640000  45.290000 74.290000  45.360000 ;
        RECT 59.640000  68.320000 74.290000  68.390000 ;
        RECT 59.640000  91.380000 74.290000  91.450000 ;
        RECT 59.640000 114.290000 74.290000 114.360000 ;
        RECT 59.640000 137.325000 74.290000 137.395000 ;
        RECT 59.640000 160.340000 74.290000 160.410000 ;
        RECT 59.640000 184.350000 74.290000 184.420000 ;
        RECT 59.655000  81.185000 74.290000  81.255000 ;
        RECT 59.655000 104.185000 74.290000 104.255000 ;
        RECT 59.655000 127.185000 74.290000 127.255000 ;
        RECT 59.655000 150.255000 74.290000 150.325000 ;
        RECT 59.665000  29.440000 74.290000  29.510000 ;
        RECT 59.665000 173.185000 74.290000 173.255000 ;
        RECT 59.695000  58.255000 74.290000  58.325000 ;
        RECT 59.710000  45.220000 74.290000  45.290000 ;
        RECT 59.710000  68.250000 74.290000  68.320000 ;
        RECT 59.710000  91.310000 74.290000  91.380000 ;
        RECT 59.710000 114.220000 74.290000 114.290000 ;
        RECT 59.710000 137.255000 74.290000 137.325000 ;
        RECT 59.710000 160.270000 74.290000 160.340000 ;
        RECT 59.710000 184.280000 74.290000 184.350000 ;
        RECT 59.725000  81.255000 74.290000  81.325000 ;
        RECT 59.725000 104.255000 74.290000 104.325000 ;
        RECT 59.725000 127.255000 74.290000 127.325000 ;
        RECT 59.725000 150.325000 74.290000 150.395000 ;
        RECT 59.735000  29.510000 74.290000  29.580000 ;
        RECT 59.735000 173.255000 74.290000 173.325000 ;
        RECT 59.765000  58.325000 74.290000  58.395000 ;
        RECT 59.780000  45.150000 74.290000  45.220000 ;
        RECT 59.780000  68.180000 74.290000  68.250000 ;
        RECT 59.780000  91.240000 74.290000  91.310000 ;
        RECT 59.780000 114.150000 74.290000 114.220000 ;
        RECT 59.780000 137.185000 74.290000 137.255000 ;
        RECT 59.780000 160.200000 74.290000 160.270000 ;
        RECT 59.780000 184.210000 74.290000 184.280000 ;
        RECT 59.795000  81.325000 74.290000  81.395000 ;
        RECT 59.795000 104.325000 74.290000 104.395000 ;
        RECT 59.795000 127.325000 74.290000 127.395000 ;
        RECT 59.795000 150.395000 74.290000 150.465000 ;
        RECT 59.805000  29.580000 74.290000  29.650000 ;
        RECT 59.805000 173.325000 74.290000 173.395000 ;
        RECT 59.835000  58.395000 74.290000  58.465000 ;
        RECT 59.850000  45.080000 74.290000  45.150000 ;
        RECT 59.850000  68.110000 74.290000  68.180000 ;
        RECT 59.850000  91.170000 74.290000  91.240000 ;
        RECT 59.850000 114.080000 74.290000 114.150000 ;
        RECT 59.850000 137.115000 74.290000 137.185000 ;
        RECT 59.850000 160.130000 74.290000 160.200000 ;
        RECT 59.850000 184.140000 74.290000 184.210000 ;
        RECT 59.865000  81.395000 74.290000  81.465000 ;
        RECT 59.865000 104.395000 74.290000 104.465000 ;
        RECT 59.865000 127.395000 74.290000 127.465000 ;
        RECT 59.865000 150.465000 74.290000 150.535000 ;
        RECT 59.875000  29.650000 74.290000  29.720000 ;
        RECT 59.875000 173.395000 74.290000 173.465000 ;
        RECT 59.905000  58.465000 74.290000  58.535000 ;
        RECT 59.920000  45.010000 74.290000  45.080000 ;
        RECT 59.920000  68.040000 74.290000  68.110000 ;
        RECT 59.920000  91.100000 74.290000  91.170000 ;
        RECT 59.920000 114.010000 74.290000 114.080000 ;
        RECT 59.920000 137.045000 74.290000 137.115000 ;
        RECT 59.920000 160.060000 74.290000 160.130000 ;
        RECT 59.920000 184.070000 74.290000 184.140000 ;
        RECT 59.935000  81.465000 74.290000  81.535000 ;
        RECT 59.935000 104.465000 74.290000 104.535000 ;
        RECT 59.935000 127.465000 74.290000 127.535000 ;
        RECT 59.935000 150.535000 74.290000 150.605000 ;
        RECT 59.945000  29.720000 74.290000  29.790000 ;
        RECT 59.945000 173.465000 74.290000 173.535000 ;
        RECT 59.975000  58.535000 74.290000  58.605000 ;
        RECT 59.990000  44.940000 74.290000  45.010000 ;
        RECT 59.990000  67.970000 74.290000  68.040000 ;
        RECT 59.990000  91.030000 74.290000  91.100000 ;
        RECT 59.990000 113.940000 74.290000 114.010000 ;
        RECT 59.990000 136.975000 74.290000 137.045000 ;
        RECT 59.990000 159.990000 74.290000 160.060000 ;
        RECT 59.990000 184.000000 74.290000 184.070000 ;
        RECT 60.005000  81.535000 74.290000  81.605000 ;
        RECT 60.005000 104.535000 74.290000 104.605000 ;
        RECT 60.005000 127.535000 74.290000 127.605000 ;
        RECT 60.005000 150.605000 74.290000 150.675000 ;
        RECT 60.015000  29.790000 74.290000  29.860000 ;
        RECT 60.015000 173.535000 74.290000 173.605000 ;
        RECT 60.045000  58.605000 74.290000  58.675000 ;
        RECT 60.060000  44.870000 74.290000  44.940000 ;
        RECT 60.060000  67.900000 74.290000  67.970000 ;
        RECT 60.060000  90.960000 74.290000  91.030000 ;
        RECT 60.060000 113.870000 74.290000 113.940000 ;
        RECT 60.060000 136.905000 74.290000 136.975000 ;
        RECT 60.060000 159.920000 74.290000 159.990000 ;
        RECT 60.060000 183.930000 74.290000 184.000000 ;
        RECT 60.075000  81.605000 74.290000  81.675000 ;
        RECT 60.075000 104.605000 74.290000 104.675000 ;
        RECT 60.075000 127.605000 74.290000 127.675000 ;
        RECT 60.075000 150.675000 74.290000 150.745000 ;
        RECT 60.085000  29.860000 74.290000  29.930000 ;
        RECT 60.085000 173.605000 74.290000 173.675000 ;
        RECT 60.115000  58.675000 74.290000  58.745000 ;
        RECT 60.130000  44.800000 74.290000  44.870000 ;
        RECT 60.130000  67.830000 74.290000  67.900000 ;
        RECT 60.130000  90.890000 74.290000  90.960000 ;
        RECT 60.130000 113.800000 74.290000 113.870000 ;
        RECT 60.130000 136.835000 74.290000 136.905000 ;
        RECT 60.130000 159.850000 74.290000 159.920000 ;
        RECT 60.130000 183.860000 74.290000 183.930000 ;
        RECT 60.145000  81.675000 74.290000  81.745000 ;
        RECT 60.145000 104.675000 74.290000 104.745000 ;
        RECT 60.145000 127.675000 74.290000 127.745000 ;
        RECT 60.145000 150.745000 74.290000 150.815000 ;
        RECT 60.155000  29.930000 74.290000  30.000000 ;
        RECT 60.155000 173.675000 74.290000 173.745000 ;
        RECT 60.185000  58.745000 74.290000  58.815000 ;
        RECT 60.200000  44.730000 74.290000  44.800000 ;
        RECT 60.200000  67.760000 74.290000  67.830000 ;
        RECT 60.200000  90.820000 74.290000  90.890000 ;
        RECT 60.200000 113.730000 74.290000 113.800000 ;
        RECT 60.200000 136.765000 74.290000 136.835000 ;
        RECT 60.200000 159.780000 74.290000 159.850000 ;
        RECT 60.200000 183.790000 74.290000 183.860000 ;
        RECT 60.215000  81.745000 74.290000  81.815000 ;
        RECT 60.215000 104.745000 74.290000 104.815000 ;
        RECT 60.215000 127.745000 74.290000 127.815000 ;
        RECT 60.215000 150.815000 74.290000 150.885000 ;
        RECT 60.225000  30.000000 74.290000  30.070000 ;
        RECT 60.225000 173.745000 74.290000 173.815000 ;
        RECT 60.255000  58.815000 74.290000  58.885000 ;
        RECT 60.270000  44.660000 74.290000  44.730000 ;
        RECT 60.270000  67.690000 74.290000  67.760000 ;
        RECT 60.270000  90.750000 74.290000  90.820000 ;
        RECT 60.270000 113.660000 74.290000 113.730000 ;
        RECT 60.270000 136.695000 74.290000 136.765000 ;
        RECT 60.270000 159.710000 74.290000 159.780000 ;
        RECT 60.270000 183.720000 74.290000 183.790000 ;
        RECT 60.285000  81.815000 74.290000  81.885000 ;
        RECT 60.285000 104.815000 74.290000 104.885000 ;
        RECT 60.285000 127.815000 74.290000 127.885000 ;
        RECT 60.285000 150.885000 74.290000 150.955000 ;
        RECT 60.295000  30.070000 74.290000  30.140000 ;
        RECT 60.295000 173.815000 74.290000 173.885000 ;
        RECT 60.325000  58.885000 74.290000  58.955000 ;
        RECT 60.340000  44.590000 74.290000  44.660000 ;
        RECT 60.340000  67.620000 74.290000  67.690000 ;
        RECT 60.340000  90.680000 74.290000  90.750000 ;
        RECT 60.340000 113.590000 74.290000 113.660000 ;
        RECT 60.340000 136.625000 74.290000 136.695000 ;
        RECT 60.340000 159.640000 74.290000 159.710000 ;
        RECT 60.340000 183.650000 74.290000 183.720000 ;
        RECT 60.355000  81.885000 74.290000  81.955000 ;
        RECT 60.355000 104.885000 74.290000 104.955000 ;
        RECT 60.355000 127.885000 74.290000 127.955000 ;
        RECT 60.355000 150.955000 74.290000 151.025000 ;
        RECT 60.365000  30.140000 74.290000  30.210000 ;
        RECT 60.365000 173.885000 74.290000 173.955000 ;
        RECT 60.395000  58.955000 74.290000  59.025000 ;
        RECT 60.410000  44.520000 74.290000  44.590000 ;
        RECT 60.410000  67.550000 74.290000  67.620000 ;
        RECT 60.410000  90.610000 74.290000  90.680000 ;
        RECT 60.410000 113.520000 74.290000 113.590000 ;
        RECT 60.410000 136.555000 74.290000 136.625000 ;
        RECT 60.410000 159.570000 74.290000 159.640000 ;
        RECT 60.410000 183.580000 74.290000 183.650000 ;
        RECT 60.425000  81.955000 74.290000  82.025000 ;
        RECT 60.425000 104.955000 74.290000 105.025000 ;
        RECT 60.425000 127.955000 74.290000 128.025000 ;
        RECT 60.425000 151.025000 74.290000 151.095000 ;
        RECT 60.435000  30.210000 74.290000  30.280000 ;
        RECT 60.435000 173.955000 74.290000 174.025000 ;
        RECT 60.465000  59.025000 74.290000  59.095000 ;
        RECT 60.480000  44.450000 74.290000  44.520000 ;
        RECT 60.480000  67.480000 74.290000  67.550000 ;
        RECT 60.480000  90.540000 74.290000  90.610000 ;
        RECT 60.480000 113.450000 74.290000 113.520000 ;
        RECT 60.480000 136.485000 74.290000 136.555000 ;
        RECT 60.480000 159.500000 74.290000 159.570000 ;
        RECT 60.480000 183.510000 74.290000 183.580000 ;
        RECT 60.495000  82.025000 74.290000  82.095000 ;
        RECT 60.495000 105.025000 74.290000 105.095000 ;
        RECT 60.495000 128.025000 74.290000 128.095000 ;
        RECT 60.495000 151.095000 74.290000 151.165000 ;
        RECT 60.505000  30.280000 74.290000  30.350000 ;
        RECT 60.505000 174.025000 74.290000 174.095000 ;
        RECT 60.535000  59.095000 74.290000  59.165000 ;
        RECT 60.550000  44.380000 74.290000  44.450000 ;
        RECT 60.550000  67.410000 74.290000  67.480000 ;
        RECT 60.550000  90.470000 74.290000  90.540000 ;
        RECT 60.550000 113.380000 74.290000 113.450000 ;
        RECT 60.550000 136.415000 74.290000 136.485000 ;
        RECT 60.550000 159.430000 74.290000 159.500000 ;
        RECT 60.550000 183.440000 74.290000 183.510000 ;
        RECT 60.565000  82.095000 74.290000  82.165000 ;
        RECT 60.565000 105.095000 74.290000 105.165000 ;
        RECT 60.565000 128.095000 74.290000 128.165000 ;
        RECT 60.565000 151.165000 74.290000 151.235000 ;
        RECT 60.575000  30.350000 74.290000  30.420000 ;
        RECT 60.575000 174.095000 74.290000 174.165000 ;
        RECT 60.605000  59.165000 74.290000  59.235000 ;
        RECT 60.620000  44.310000 74.290000  44.380000 ;
        RECT 60.620000  67.340000 74.290000  67.410000 ;
        RECT 60.620000  90.400000 74.290000  90.470000 ;
        RECT 60.620000 113.310000 74.290000 113.380000 ;
        RECT 60.620000 136.345000 74.290000 136.415000 ;
        RECT 60.620000 159.360000 74.290000 159.430000 ;
        RECT 60.620000 183.370000 74.290000 183.440000 ;
        RECT 60.635000  82.165000 74.290000  82.235000 ;
        RECT 60.635000 105.165000 74.290000 105.235000 ;
        RECT 60.635000 128.165000 74.290000 128.235000 ;
        RECT 60.635000 151.235000 74.290000 151.305000 ;
        RECT 60.645000  30.420000 74.290000  30.490000 ;
        RECT 60.645000 174.165000 74.290000 174.235000 ;
        RECT 60.675000  59.235000 74.290000  59.305000 ;
        RECT 60.690000  44.240000 74.290000  44.310000 ;
        RECT 60.690000  67.270000 74.290000  67.340000 ;
        RECT 60.690000  90.330000 74.290000  90.400000 ;
        RECT 60.690000 113.240000 74.290000 113.310000 ;
        RECT 60.690000 136.275000 74.290000 136.345000 ;
        RECT 60.690000 159.290000 74.290000 159.360000 ;
        RECT 60.690000 183.300000 74.290000 183.370000 ;
        RECT 60.705000  82.235000 74.290000  82.305000 ;
        RECT 60.705000 105.235000 74.290000 105.305000 ;
        RECT 60.705000 128.235000 74.290000 128.305000 ;
        RECT 60.705000 151.305000 74.290000 151.375000 ;
        RECT 60.715000  30.490000 74.290000  30.560000 ;
        RECT 60.715000 174.235000 74.290000 174.305000 ;
        RECT 60.745000  59.305000 74.290000  59.375000 ;
        RECT 60.760000  44.170000 74.290000  44.240000 ;
        RECT 60.760000  67.200000 74.290000  67.270000 ;
        RECT 60.760000  90.260000 74.290000  90.330000 ;
        RECT 60.760000 113.170000 74.290000 113.240000 ;
        RECT 60.760000 136.205000 74.290000 136.275000 ;
        RECT 60.760000 159.220000 74.290000 159.290000 ;
        RECT 60.760000 183.230000 74.290000 183.300000 ;
        RECT 60.775000  82.305000 74.290000  82.375000 ;
        RECT 60.775000 105.305000 74.290000 105.375000 ;
        RECT 60.775000 128.305000 74.290000 128.375000 ;
        RECT 60.775000 151.375000 74.290000 151.445000 ;
        RECT 60.785000  30.560000 74.290000  30.630000 ;
        RECT 60.785000 174.305000 74.290000 174.375000 ;
        RECT 60.815000  59.375000 74.290000  59.445000 ;
        RECT 60.830000  44.100000 74.290000  44.170000 ;
        RECT 60.830000  67.130000 74.290000  67.200000 ;
        RECT 60.830000  90.190000 74.290000  90.260000 ;
        RECT 60.830000 113.100000 74.290000 113.170000 ;
        RECT 60.830000 136.135000 74.290000 136.205000 ;
        RECT 60.830000 159.150000 74.290000 159.220000 ;
        RECT 60.830000 183.160000 74.290000 183.230000 ;
        RECT 60.845000  82.375000 74.290000  82.445000 ;
        RECT 60.845000 105.375000 74.290000 105.445000 ;
        RECT 60.845000 128.375000 74.290000 128.445000 ;
        RECT 60.845000 151.445000 74.290000 151.515000 ;
        RECT 60.855000  30.630000 74.290000  30.700000 ;
        RECT 60.855000 174.375000 74.290000 174.445000 ;
        RECT 60.885000  59.445000 74.290000  59.515000 ;
        RECT 60.900000  44.030000 74.290000  44.100000 ;
        RECT 60.900000  67.060000 74.290000  67.130000 ;
        RECT 60.900000  90.120000 74.290000  90.190000 ;
        RECT 60.900000 113.030000 74.290000 113.100000 ;
        RECT 60.900000 136.065000 74.290000 136.135000 ;
        RECT 60.900000 159.080000 74.290000 159.150000 ;
        RECT 60.900000 183.090000 74.290000 183.160000 ;
        RECT 60.915000  82.445000 74.290000  82.515000 ;
        RECT 60.915000 105.445000 74.290000 105.515000 ;
        RECT 60.915000 128.445000 74.290000 128.515000 ;
        RECT 60.915000 151.515000 74.290000 151.585000 ;
        RECT 60.925000  30.700000 74.290000  30.770000 ;
        RECT 60.925000 174.445000 74.290000 174.515000 ;
        RECT 60.955000  59.515000 74.290000  59.585000 ;
        RECT 60.970000  43.960000 74.290000  44.030000 ;
        RECT 60.970000  66.990000 74.290000  67.060000 ;
        RECT 60.970000  90.050000 74.290000  90.120000 ;
        RECT 60.970000 112.960000 74.290000 113.030000 ;
        RECT 60.970000 135.995000 74.290000 136.065000 ;
        RECT 60.970000 159.010000 74.290000 159.080000 ;
        RECT 60.970000 183.020000 74.290000 183.090000 ;
        RECT 60.985000  82.515000 74.290000  82.585000 ;
        RECT 60.985000 105.515000 74.290000 105.585000 ;
        RECT 60.985000 128.515000 74.290000 128.585000 ;
        RECT 60.985000 151.585000 74.290000 151.655000 ;
        RECT 60.995000  30.770000 74.290000  30.840000 ;
        RECT 60.995000 174.515000 74.290000 174.585000 ;
        RECT 61.025000  59.585000 74.290000  59.655000 ;
        RECT 61.040000  43.890000 74.290000  43.960000 ;
        RECT 61.040000  66.920000 74.290000  66.990000 ;
        RECT 61.040000  89.980000 74.290000  90.050000 ;
        RECT 61.040000 112.890000 74.290000 112.960000 ;
        RECT 61.040000 135.925000 74.290000 135.995000 ;
        RECT 61.040000 158.940000 74.290000 159.010000 ;
        RECT 61.040000 182.950000 74.290000 183.020000 ;
        RECT 61.055000  82.585000 74.290000  82.655000 ;
        RECT 61.055000 105.585000 74.290000 105.655000 ;
        RECT 61.055000 128.585000 74.290000 128.655000 ;
        RECT 61.055000 151.655000 74.290000 151.725000 ;
        RECT 61.065000  30.840000 74.290000  30.910000 ;
        RECT 61.065000 174.585000 74.290000 174.655000 ;
        RECT 61.095000  59.655000 74.290000  59.725000 ;
        RECT 61.110000  30.910000 74.290000  30.955000 ;
        RECT 61.110000  30.955000 74.290000  43.820000 ;
        RECT 61.110000  43.820000 74.290000  43.890000 ;
        RECT 61.110000  59.725000 74.290000  59.740000 ;
        RECT 61.110000  59.740000 74.290000  66.850000 ;
        RECT 61.110000  66.850000 74.290000  66.920000 ;
        RECT 61.110000  82.655000 74.290000  82.710000 ;
        RECT 61.110000  82.710000 74.290000  89.910000 ;
        RECT 61.110000  89.910000 74.290000  89.980000 ;
        RECT 61.110000 105.655000 74.290000 105.710000 ;
        RECT 61.110000 105.710000 74.290000 112.820000 ;
        RECT 61.110000 112.820000 74.290000 112.890000 ;
        RECT 61.110000 128.655000 74.290000 128.710000 ;
        RECT 61.110000 128.710000 74.290000 135.855000 ;
        RECT 61.110000 135.855000 74.290000 135.925000 ;
        RECT 61.110000 151.725000 74.290000 151.780000 ;
        RECT 61.110000 151.780000 74.290000 158.870000 ;
        RECT 61.110000 158.870000 74.290000 158.940000 ;
        RECT 61.110000 174.655000 74.290000 174.700000 ;
        RECT 61.110000 174.700000 74.290000 182.880000 ;
        RECT 61.110000 182.880000 74.290000 182.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000   0.000000 48.890000  96.150000 ;
        RECT 37.890000  96.150000 48.890000  96.300000 ;
        RECT 37.890000  96.300000 49.040000  96.450000 ;
        RECT 37.890000  96.450000 49.190000  96.600000 ;
        RECT 37.890000  96.600000 49.340000  96.750000 ;
        RECT 37.890000  96.750000 49.490000  96.900000 ;
        RECT 37.890000  96.900000 49.640000  97.050000 ;
        RECT 37.890000  97.050000 49.790000  97.200000 ;
        RECT 37.890000  97.200000 49.940000  97.350000 ;
        RECT 37.890000  97.350000 50.090000  97.500000 ;
        RECT 37.890000  97.500000 50.240000  97.650000 ;
        RECT 37.890000  97.650000 50.390000  97.800000 ;
        RECT 37.890000  97.800000 50.540000  97.950000 ;
        RECT 37.890000  97.950000 50.690000  98.100000 ;
        RECT 37.890000  98.100000 50.840000  98.250000 ;
        RECT 37.890000  98.250000 50.990000  98.300000 ;
        RECT 37.890000  98.300000 51.040000  99.505000 ;
        RECT 37.890000  99.505000 43.400000  99.655000 ;
        RECT 37.890000  99.655000 43.250000  99.805000 ;
        RECT 37.890000  99.805000 43.100000  99.955000 ;
        RECT 37.890000  99.955000 42.950000 100.105000 ;
        RECT 37.890000 100.105000 42.840000 100.215000 ;
        RECT 37.890000 100.215000 42.840000 102.135000 ;
        RECT 37.890000 102.135000 42.840000 102.285000 ;
        RECT 37.890000 102.285000 42.990000 102.435000 ;
        RECT 37.890000 102.435000 43.140000 102.585000 ;
        RECT 37.890000 102.585000 43.290000 102.735000 ;
        RECT 37.890000 102.735000 43.440000 102.885000 ;
        RECT 37.890000 102.885000 43.590000 103.035000 ;
        RECT 37.890000 103.035000 43.740000 103.185000 ;
        RECT 37.890000 103.185000 43.890000 103.335000 ;
        RECT 37.890000 103.335000 44.040000 103.485000 ;
        RECT 37.890000 103.485000 44.190000 103.635000 ;
        RECT 37.890000 103.635000 44.340000 103.785000 ;
        RECT 37.890000 103.785000 44.490000 103.935000 ;
        RECT 37.890000 103.935000 44.640000 104.085000 ;
        RECT 37.890000 104.085000 44.790000 104.235000 ;
        RECT 37.890000 104.235000 44.940000 104.385000 ;
        RECT 37.890000 104.385000 45.090000 104.535000 ;
        RECT 37.890000 104.535000 45.240000 104.685000 ;
        RECT 37.890000 104.685000 45.390000 104.835000 ;
        RECT 37.890000 104.835000 45.540000 104.985000 ;
        RECT 37.890000 104.985000 45.690000 105.135000 ;
        RECT 37.890000 105.135000 45.840000 105.285000 ;
        RECT 37.890000 105.285000 45.990000 105.435000 ;
        RECT 37.890000 105.435000 46.140000 105.585000 ;
        RECT 37.890000 105.585000 46.290000 105.655000 ;
        RECT 37.965000 175.350000 48.855000 190.020000 ;
        RECT 38.040000 105.655000 46.360000 105.805000 ;
        RECT 38.055000 175.260000 48.855000 175.350000 ;
        RECT 38.190000 105.805000 46.510000 105.955000 ;
        RECT 38.205000 175.110000 48.855000 175.260000 ;
        RECT 38.340000 105.955000 46.660000 106.105000 ;
        RECT 38.355000 174.960000 48.855000 175.110000 ;
        RECT 38.490000 106.105000 46.810000 106.255000 ;
        RECT 38.505000 174.810000 48.855000 174.960000 ;
        RECT 38.640000 106.255000 46.960000 106.405000 ;
        RECT 38.655000 174.660000 48.855000 174.810000 ;
        RECT 38.790000 106.405000 47.110000 106.555000 ;
        RECT 38.805000 174.510000 48.855000 174.660000 ;
        RECT 38.940000 106.555000 47.260000 106.705000 ;
        RECT 38.955000 174.360000 48.855000 174.510000 ;
        RECT 39.090000 106.705000 47.410000 106.855000 ;
        RECT 39.105000 174.210000 48.855000 174.360000 ;
        RECT 39.240000 106.855000 47.560000 107.005000 ;
        RECT 39.255000 174.060000 48.855000 174.210000 ;
        RECT 39.390000 107.005000 47.710000 107.155000 ;
        RECT 39.405000 173.910000 48.855000 174.060000 ;
        RECT 39.540000 107.155000 47.860000 107.305000 ;
        RECT 39.555000 173.760000 48.855000 173.910000 ;
        RECT 39.690000 107.305000 48.010000 107.455000 ;
        RECT 39.705000 173.610000 48.855000 173.760000 ;
        RECT 39.840000 107.455000 48.160000 107.605000 ;
        RECT 39.855000 173.460000 48.855000 173.610000 ;
        RECT 39.990000 107.605000 48.310000 107.755000 ;
        RECT 40.005000 173.310000 48.855000 173.460000 ;
        RECT 40.140000 107.755000 48.460000 107.905000 ;
        RECT 40.155000 173.160000 48.855000 173.310000 ;
        RECT 40.290000 107.905000 48.610000 108.055000 ;
        RECT 40.305000 173.010000 48.855000 173.160000 ;
        RECT 40.385000 108.055000 48.760000 108.150000 ;
        RECT 40.455000 172.860000 48.855000 173.010000 ;
        RECT 40.535000 108.150000 48.855000 108.300000 ;
        RECT 40.605000 172.710000 48.855000 172.860000 ;
        RECT 40.685000 108.300000 48.855000 108.450000 ;
        RECT 40.755000 172.560000 48.855000 172.710000 ;
        RECT 40.835000 108.450000 48.855000 108.600000 ;
        RECT 40.905000 172.410000 48.855000 172.560000 ;
        RECT 40.985000 108.600000 48.855000 108.750000 ;
        RECT 41.055000 172.260000 48.855000 172.410000 ;
        RECT 41.135000 108.750000 48.855000 108.900000 ;
        RECT 41.205000 172.110000 48.855000 172.260000 ;
        RECT 41.285000 108.900000 48.855000 109.050000 ;
        RECT 41.355000 171.960000 48.855000 172.110000 ;
        RECT 41.435000 109.050000 48.855000 109.200000 ;
        RECT 41.505000 171.810000 48.855000 171.960000 ;
        RECT 41.585000 109.200000 48.855000 109.350000 ;
        RECT 41.655000 171.660000 48.855000 171.810000 ;
        RECT 41.735000 109.350000 48.855000 109.500000 ;
        RECT 41.805000 171.510000 48.855000 171.660000 ;
        RECT 41.885000 109.500000 48.855000 109.650000 ;
        RECT 41.955000 171.360000 48.855000 171.510000 ;
        RECT 42.035000 109.650000 48.855000 109.800000 ;
        RECT 42.105000 171.210000 48.855000 171.360000 ;
        RECT 42.185000 109.800000 48.855000 109.950000 ;
        RECT 42.255000 171.060000 48.855000 171.210000 ;
        RECT 42.335000 109.950000 48.855000 110.100000 ;
        RECT 42.405000 170.910000 48.855000 171.060000 ;
        RECT 42.485000 110.100000 48.855000 110.250000 ;
        RECT 42.555000 170.760000 48.855000 170.910000 ;
        RECT 42.635000 110.250000 48.855000 110.400000 ;
        RECT 42.705000 170.610000 48.855000 170.760000 ;
        RECT 42.785000 110.400000 48.855000 110.550000 ;
        RECT 42.855000 110.550000 48.855000 110.620000 ;
        RECT 42.855000 110.620000 48.855000 170.460000 ;
        RECT 42.855000 170.460000 48.855000 170.610000 ;
        RECT 44.655000  99.505000 51.040000  99.610000 ;
        RECT 44.760000  99.610000 51.040000  99.715000 ;
        RECT 44.910000  99.715000 51.040000  99.865000 ;
        RECT 45.060000  99.865000 51.190000 100.015000 ;
        RECT 45.210000 100.015000 51.340000 100.165000 ;
        RECT 45.260000 100.165000 51.490000 100.215000 ;
        RECT 45.260000 100.215000 51.540000 100.365000 ;
        RECT 45.260000 100.365000 51.690000 100.515000 ;
        RECT 45.260000 100.515000 51.840000 100.665000 ;
        RECT 45.260000 100.665000 51.990000 100.815000 ;
        RECT 45.260000 100.815000 52.140000 100.965000 ;
        RECT 45.260000 100.965000 52.290000 101.115000 ;
        RECT 45.260000 101.115000 52.440000 101.265000 ;
        RECT 45.260000 101.265000 52.590000 101.415000 ;
        RECT 45.260000 101.415000 52.740000 101.565000 ;
        RECT 45.260000 101.565000 52.890000 101.715000 ;
        RECT 45.260000 101.715000 53.040000 101.865000 ;
        RECT 45.260000 101.865000 53.190000 102.015000 ;
        RECT 45.260000 102.015000 53.340000 102.165000 ;
        RECT 45.260000 102.165000 53.490000 102.315000 ;
        RECT 45.260000 102.315000 53.640000 102.415000 ;
        RECT 45.410000 102.415000 53.740000 102.565000 ;
        RECT 45.560000 102.565000 53.890000 102.715000 ;
        RECT 45.710000 102.715000 54.040000 102.865000 ;
        RECT 45.860000 102.865000 54.190000 103.015000 ;
        RECT 46.010000 103.015000 54.340000 103.165000 ;
        RECT 46.160000 103.165000 54.490000 103.315000 ;
        RECT 46.310000 103.315000 54.640000 103.465000 ;
        RECT 46.460000 103.465000 54.790000 103.615000 ;
        RECT 46.610000 103.615000 54.940000 103.765000 ;
        RECT 46.760000 103.765000 55.090000 103.915000 ;
        RECT 46.910000 103.915000 55.240000 104.065000 ;
        RECT 47.060000 104.065000 55.390000 104.215000 ;
        RECT 47.210000 104.215000 55.540000 104.365000 ;
        RECT 47.360000 104.365000 55.690000 104.515000 ;
        RECT 47.510000 104.515000 55.840000 104.665000 ;
        RECT 47.660000 104.665000 55.990000 104.815000 ;
        RECT 47.810000 104.815000 56.140000 104.965000 ;
        RECT 47.960000 104.965000 56.290000 105.115000 ;
        RECT 48.110000 105.115000 56.440000 105.265000 ;
        RECT 48.260000 105.265000 56.590000 105.415000 ;
        RECT 48.410000 105.415000 56.740000 105.565000 ;
        RECT 48.560000 105.565000 56.890000 105.715000 ;
        RECT 48.710000 105.715000 57.040000 105.865000 ;
        RECT 48.860000 105.865000 57.190000 106.015000 ;
        RECT 49.010000 106.015000 57.340000 106.165000 ;
        RECT 49.160000 106.165000 57.490000 106.315000 ;
        RECT 49.310000 106.315000 57.640000 106.465000 ;
        RECT 49.460000 106.465000 57.790000 106.615000 ;
        RECT 49.610000 106.615000 57.940000 106.765000 ;
        RECT 49.760000 106.765000 58.090000 106.915000 ;
        RECT 49.775000 172.645000 59.285000 173.020000 ;
        RECT 49.775000 173.020000 59.285000 173.170000 ;
        RECT 49.775000 173.170000 59.435000 173.320000 ;
        RECT 49.775000 173.320000 59.585000 173.470000 ;
        RECT 49.775000 173.470000 59.735000 173.620000 ;
        RECT 49.775000 173.620000 59.885000 173.770000 ;
        RECT 49.775000 173.770000 60.035000 173.920000 ;
        RECT 49.775000 173.920000 60.185000 174.070000 ;
        RECT 49.775000 174.070000 60.335000 174.220000 ;
        RECT 49.775000 174.220000 60.485000 174.370000 ;
        RECT 49.775000 174.370000 60.635000 174.520000 ;
        RECT 49.775000 174.520000 60.785000 174.670000 ;
        RECT 49.775000 174.670000 60.935000 174.820000 ;
        RECT 49.775000 174.820000 61.085000 174.970000 ;
        RECT 49.775000 174.970000 61.235000 175.120000 ;
        RECT 49.775000 175.120000 61.385000 175.270000 ;
        RECT 49.775000 175.270000 61.535000 175.420000 ;
        RECT 49.775000 175.420000 61.685000 175.570000 ;
        RECT 49.775000 175.570000 61.835000 175.720000 ;
        RECT 49.775000 175.720000 61.985000 175.870000 ;
        RECT 49.775000 175.870000 62.135000 176.020000 ;
        RECT 49.775000 176.020000 62.285000 176.170000 ;
        RECT 49.775000 176.170000 62.435000 176.320000 ;
        RECT 49.775000 176.320000 62.585000 176.470000 ;
        RECT 49.775000 176.470000 62.735000 176.620000 ;
        RECT 49.775000 176.620000 62.885000 176.770000 ;
        RECT 49.775000 176.770000 63.035000 176.920000 ;
        RECT 49.775000 176.920000 63.185000 177.070000 ;
        RECT 49.775000 177.070000 63.335000 177.220000 ;
        RECT 49.775000 177.220000 63.485000 177.370000 ;
        RECT 49.775000 177.370000 63.635000 177.520000 ;
        RECT 49.775000 177.520000 63.785000 177.670000 ;
        RECT 49.775000 177.670000 63.935000 177.820000 ;
        RECT 49.775000 177.820000 64.085000 177.970000 ;
        RECT 49.775000 177.970000 64.235000 178.120000 ;
        RECT 49.775000 178.120000 64.385000 178.270000 ;
        RECT 49.775000 178.270000 64.535000 178.420000 ;
        RECT 49.775000 178.420000 64.685000 178.570000 ;
        RECT 49.775000 178.570000 64.835000 178.720000 ;
        RECT 49.775000 178.720000 64.985000 178.870000 ;
        RECT 49.775000 178.870000 65.135000 179.020000 ;
        RECT 49.775000 179.020000 65.285000 179.170000 ;
        RECT 49.775000 179.170000 65.435000 179.320000 ;
        RECT 49.775000 179.320000 65.585000 179.470000 ;
        RECT 49.775000 179.470000 65.735000 179.620000 ;
        RECT 49.775000 179.620000 65.885000 179.770000 ;
        RECT 49.775000 179.770000 66.035000 179.920000 ;
        RECT 49.775000 179.920000 66.185000 180.070000 ;
        RECT 49.775000 180.070000 66.335000 180.220000 ;
        RECT 49.775000 180.220000 66.485000 180.370000 ;
        RECT 49.775000 180.370000 66.635000 180.520000 ;
        RECT 49.775000 180.520000 66.785000 180.670000 ;
        RECT 49.775000 180.670000 66.935000 180.820000 ;
        RECT 49.775000 180.820000 67.085000 180.970000 ;
        RECT 49.775000 180.970000 67.235000 181.120000 ;
        RECT 49.775000 181.120000 67.385000 181.270000 ;
        RECT 49.775000 181.270000 67.535000 181.420000 ;
        RECT 49.775000 181.420000 67.685000 181.570000 ;
        RECT 49.775000 181.570000 67.835000 181.720000 ;
        RECT 49.775000 181.720000 67.985000 181.870000 ;
        RECT 49.775000 181.870000 68.135000 182.020000 ;
        RECT 49.775000 182.020000 68.285000 182.170000 ;
        RECT 49.775000 182.170000 68.435000 182.320000 ;
        RECT 49.775000 182.320000 68.585000 182.470000 ;
        RECT 49.775000 182.470000 68.735000 182.620000 ;
        RECT 49.775000 182.620000 68.885000 182.770000 ;
        RECT 49.775000 182.770000 69.035000 182.920000 ;
        RECT 49.775000 182.920000 69.185000 183.070000 ;
        RECT 49.775000 183.070000 69.335000 183.220000 ;
        RECT 49.775000 183.220000 69.485000 183.370000 ;
        RECT 49.775000 183.370000 69.635000 183.520000 ;
        RECT 49.775000 183.520000 69.785000 183.670000 ;
        RECT 49.775000 183.670000 69.935000 183.820000 ;
        RECT 49.775000 183.820000 70.085000 183.970000 ;
        RECT 49.775000 183.970000 70.235000 184.120000 ;
        RECT 49.775000 184.120000 70.385000 184.270000 ;
        RECT 49.775000 184.270000 70.535000 184.420000 ;
        RECT 49.775000 184.420000 70.685000 184.570000 ;
        RECT 49.775000 184.570000 70.835000 184.720000 ;
        RECT 49.775000 184.720000 70.985000 184.870000 ;
        RECT 49.775000 184.870000 71.135000 185.020000 ;
        RECT 49.775000 185.020000 71.285000 185.170000 ;
        RECT 49.775000 185.170000 71.435000 185.320000 ;
        RECT 49.775000 185.320000 71.585000 185.360000 ;
        RECT 49.775000 185.360000 71.625000 190.040000 ;
        RECT 49.835000 172.585000 59.285000 172.645000 ;
        RECT 49.910000 106.915000 58.240000 107.065000 ;
        RECT 49.985000 172.435000 59.285000 172.585000 ;
        RECT 50.060000 107.065000 58.390000 107.215000 ;
        RECT 50.135000 172.285000 59.285000 172.435000 ;
        RECT 50.210000 107.215000 58.540000 107.365000 ;
        RECT 50.285000 172.135000 59.285000 172.285000 ;
        RECT 50.360000 107.365000 58.690000 107.515000 ;
        RECT 50.435000 171.985000 59.285000 172.135000 ;
        RECT 50.510000 107.515000 58.840000 107.665000 ;
        RECT 50.585000 171.835000 59.285000 171.985000 ;
        RECT 50.660000 107.665000 58.990000 107.815000 ;
        RECT 50.735000 171.685000 59.285000 171.835000 ;
        RECT 50.805000 107.815000 59.140000 107.960000 ;
        RECT 50.885000 171.535000 59.285000 171.685000 ;
        RECT 50.955000 107.960000 59.285000 108.110000 ;
        RECT 51.035000 171.385000 59.285000 171.535000 ;
        RECT 51.105000 108.110000 59.285000 108.260000 ;
        RECT 51.185000 171.235000 59.285000 171.385000 ;
        RECT 51.255000 108.260000 59.285000 108.410000 ;
        RECT 51.335000 171.085000 59.285000 171.235000 ;
        RECT 51.405000 108.410000 59.285000 108.560000 ;
        RECT 51.485000 170.935000 59.285000 171.085000 ;
        RECT 51.555000 108.560000 59.285000 108.710000 ;
        RECT 51.635000 170.785000 59.285000 170.935000 ;
        RECT 51.705000 108.710000 59.285000 108.860000 ;
        RECT 51.785000 170.635000 59.285000 170.785000 ;
        RECT 51.855000 108.860000 59.285000 109.010000 ;
        RECT 51.935000 170.485000 59.285000 170.635000 ;
        RECT 52.005000 109.010000 59.285000 109.160000 ;
        RECT 52.085000 170.335000 59.285000 170.485000 ;
        RECT 52.155000 109.160000 59.285000 109.310000 ;
        RECT 52.235000 170.185000 59.285000 170.335000 ;
        RECT 52.305000 109.310000 59.285000 109.460000 ;
        RECT 52.385000 170.035000 59.285000 170.185000 ;
        RECT 52.455000 109.460000 59.285000 109.610000 ;
        RECT 52.535000 169.885000 59.285000 170.035000 ;
        RECT 52.605000 109.610000 59.285000 109.760000 ;
        RECT 52.685000 169.735000 59.285000 169.885000 ;
        RECT 52.755000 109.760000 59.285000 109.910000 ;
        RECT 52.835000 169.585000 59.285000 169.735000 ;
        RECT 52.905000 109.910000 59.285000 110.060000 ;
        RECT 52.985000 169.435000 59.285000 169.585000 ;
        RECT 53.055000 110.060000 59.285000 110.210000 ;
        RECT 53.135000 169.285000 59.285000 169.435000 ;
        RECT 53.205000 110.210000 59.285000 110.360000 ;
        RECT 53.285000 110.360000 59.285000 110.440000 ;
        RECT 53.285000 110.440000 59.285000 169.135000 ;
        RECT 53.285000 169.135000 59.285000 169.285000 ;
    END
  END DRN_HVC
  PIN OGC_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 25.895000 0.000000 27.895000 0.535000 ;
    END
  END OGC_HVC
  PIN P_CORE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.495000   0.000000 24.395000  36.510000 ;
        RECT 0.495000  46.960000 24.395000  90.500000 ;
        RECT 0.495000  90.500000 24.245000  90.650000 ;
        RECT 0.495000  90.650000 24.095000  90.800000 ;
        RECT 0.495000  90.800000 23.945000  90.950000 ;
        RECT 0.495000  90.950000 23.795000  91.100000 ;
        RECT 0.495000  91.100000 23.645000  91.250000 ;
        RECT 0.495000  91.250000 23.495000  91.400000 ;
        RECT 0.495000  91.400000 23.345000  91.550000 ;
        RECT 0.495000  91.550000 23.195000  91.700000 ;
        RECT 0.495000  91.700000 23.045000  91.850000 ;
        RECT 0.495000  91.850000 22.895000  92.000000 ;
        RECT 0.495000  92.000000 22.745000  92.150000 ;
        RECT 0.495000  92.150000 22.595000  92.300000 ;
        RECT 0.495000  92.300000 22.445000  92.450000 ;
        RECT 0.495000  92.450000 22.295000  92.600000 ;
        RECT 0.495000  92.600000 22.145000  92.750000 ;
        RECT 0.495000  92.750000 21.995000  92.900000 ;
        RECT 0.495000  92.900000 21.845000  93.050000 ;
        RECT 0.495000  93.050000 21.695000  93.200000 ;
        RECT 0.495000  93.200000 21.545000  93.350000 ;
        RECT 0.495000  93.350000 21.395000  93.500000 ;
        RECT 0.495000  93.500000 21.245000  93.650000 ;
        RECT 0.495000  93.650000 21.095000  93.800000 ;
        RECT 0.495000  93.800000 20.945000  93.950000 ;
        RECT 0.495000  93.950000 20.795000  94.100000 ;
        RECT 0.495000  94.100000 20.645000  94.250000 ;
        RECT 0.495000  94.250000 20.495000  94.400000 ;
        RECT 0.495000  94.400000 20.345000  94.550000 ;
        RECT 0.495000  94.550000 20.195000  94.700000 ;
        RECT 0.495000  94.700000 20.045000  94.850000 ;
        RECT 0.495000  94.850000 19.895000  95.000000 ;
        RECT 0.495000  95.000000 19.745000  95.150000 ;
        RECT 0.495000  95.150000 19.595000  95.300000 ;
        RECT 0.495000  95.300000 19.445000  95.450000 ;
        RECT 0.495000  95.450000 19.295000  95.600000 ;
        RECT 0.495000  95.600000 19.145000  95.750000 ;
        RECT 0.495000  95.750000 18.995000  95.900000 ;
        RECT 0.495000  95.900000 18.845000  96.050000 ;
        RECT 0.495000  96.050000 18.695000  96.200000 ;
        RECT 0.495000  96.200000 18.545000  96.350000 ;
        RECT 0.495000  96.350000 18.395000  96.500000 ;
        RECT 0.495000  96.500000 18.245000  96.650000 ;
        RECT 0.495000  96.650000 18.095000  96.800000 ;
        RECT 0.495000  96.800000 17.945000  96.950000 ;
        RECT 0.495000  96.950000 17.795000  97.100000 ;
        RECT 0.495000  97.100000 17.645000  97.250000 ;
        RECT 0.495000  97.250000 17.495000  97.400000 ;
        RECT 0.495000  97.400000 17.345000  97.550000 ;
        RECT 0.495000  97.550000 17.195000  97.700000 ;
        RECT 0.495000  97.700000 17.045000  97.850000 ;
        RECT 0.495000  97.850000 16.895000  98.000000 ;
        RECT 0.495000  98.000000 16.745000  98.150000 ;
        RECT 0.495000  98.150000 16.595000  98.300000 ;
        RECT 0.495000  98.300000 16.445000  98.450000 ;
        RECT 0.495000  98.450000 16.295000  98.600000 ;
        RECT 0.495000  98.600000 16.145000  98.750000 ;
        RECT 0.495000  98.750000 15.995000  98.900000 ;
        RECT 0.495000  98.900000 15.845000  99.050000 ;
        RECT 0.495000  99.050000 15.695000  99.200000 ;
        RECT 0.495000  99.200000 15.545000  99.350000 ;
        RECT 0.495000  99.350000 15.395000  99.500000 ;
        RECT 0.495000  99.500000 15.245000  99.650000 ;
        RECT 0.495000  99.650000 15.095000  99.800000 ;
        RECT 0.495000  99.800000 14.945000  99.950000 ;
        RECT 0.495000  99.950000 14.795000 100.100000 ;
        RECT 0.495000 100.100000 14.645000 100.250000 ;
        RECT 0.495000 100.250000 14.495000 100.400000 ;
        RECT 0.495000 100.400000 14.345000 100.550000 ;
        RECT 0.495000 100.550000 14.195000 100.700000 ;
        RECT 0.495000 100.700000 14.045000 100.850000 ;
        RECT 0.495000 100.850000 13.895000 101.000000 ;
        RECT 0.495000 101.000000 13.745000 101.150000 ;
        RECT 0.495000 101.150000 13.595000 101.300000 ;
        RECT 0.495000 101.300000 13.500000 101.395000 ;
        RECT 0.495000 101.395000 13.500000 173.155000 ;
        RECT 0.510000  46.945000 24.395000  46.960000 ;
        RECT 0.645000  36.510000 24.395000  36.660000 ;
        RECT 0.660000  46.795000 24.395000  46.945000 ;
        RECT 0.795000  36.660000 24.395000  36.810000 ;
        RECT 0.810000  46.645000 24.395000  46.795000 ;
        RECT 0.945000  36.810000 24.395000  36.960000 ;
        RECT 0.960000  46.495000 24.395000  46.645000 ;
        RECT 1.095000  36.960000 24.395000  37.110000 ;
        RECT 1.110000  37.110000 24.395000  37.125000 ;
        RECT 1.110000  37.125000 24.395000  46.345000 ;
        RECT 1.110000  46.345000 24.395000  46.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000   0.000000 74.290000  90.185000 ;
        RECT 50.540000  90.185000 74.290000  90.335000 ;
        RECT 50.690000  90.335000 74.290000  90.485000 ;
        RECT 50.840000  90.485000 74.290000  90.635000 ;
        RECT 50.990000  90.635000 74.290000  90.785000 ;
        RECT 51.140000  90.785000 74.290000  90.935000 ;
        RECT 51.290000  90.935000 74.290000  91.085000 ;
        RECT 51.440000  91.085000 74.290000  91.235000 ;
        RECT 51.590000  91.235000 74.290000  91.385000 ;
        RECT 51.740000  91.385000 74.290000  91.535000 ;
        RECT 51.890000  91.535000 74.290000  91.685000 ;
        RECT 52.040000  91.685000 74.290000  91.835000 ;
        RECT 52.190000  91.835000 74.290000  91.985000 ;
        RECT 52.340000  91.985000 74.290000  92.135000 ;
        RECT 52.490000  92.135000 74.290000  92.285000 ;
        RECT 52.640000  92.285000 74.290000  92.435000 ;
        RECT 52.790000  92.435000 74.290000  92.585000 ;
        RECT 52.940000  92.585000 74.290000  92.735000 ;
        RECT 53.090000  92.735000 74.290000  92.885000 ;
        RECT 53.240000  92.885000 74.290000  93.035000 ;
        RECT 53.390000  93.035000 74.290000  93.185000 ;
        RECT 53.540000  93.185000 74.290000  93.335000 ;
        RECT 53.690000  93.335000 74.290000  93.485000 ;
        RECT 53.840000  93.485000 74.290000  93.635000 ;
        RECT 53.990000  93.635000 74.290000  93.785000 ;
        RECT 54.140000  93.785000 74.290000  93.935000 ;
        RECT 54.290000  93.935000 74.290000  94.085000 ;
        RECT 54.440000  94.085000 74.290000  94.235000 ;
        RECT 54.590000  94.235000 74.290000  94.385000 ;
        RECT 54.740000  94.385000 74.290000  94.535000 ;
        RECT 54.890000  94.535000 74.290000  94.685000 ;
        RECT 55.040000  94.685000 74.290000  94.835000 ;
        RECT 55.190000  94.835000 74.290000  94.985000 ;
        RECT 55.340000  94.985000 74.290000  95.135000 ;
        RECT 55.490000  95.135000 74.290000  95.285000 ;
        RECT 55.640000  95.285000 74.290000  95.435000 ;
        RECT 55.790000  95.435000 74.290000  95.585000 ;
        RECT 55.940000  95.585000 74.290000  95.735000 ;
        RECT 56.090000  95.735000 74.290000  95.885000 ;
        RECT 56.240000  95.885000 74.290000  96.035000 ;
        RECT 56.390000  96.035000 74.290000  96.185000 ;
        RECT 56.540000  96.185000 74.290000  96.335000 ;
        RECT 56.690000  96.335000 74.290000  96.485000 ;
        RECT 56.840000  96.485000 74.290000  96.635000 ;
        RECT 56.990000  96.635000 74.290000  96.785000 ;
        RECT 57.140000  96.785000 74.290000  96.935000 ;
        RECT 57.290000  96.935000 74.290000  97.085000 ;
        RECT 57.440000  97.085000 74.290000  97.235000 ;
        RECT 57.590000  97.235000 74.290000  97.385000 ;
        RECT 57.740000  97.385000 74.290000  97.535000 ;
        RECT 57.890000  97.535000 74.290000  97.685000 ;
        RECT 58.040000  97.685000 74.290000  97.835000 ;
        RECT 58.190000  97.835000 74.290000  97.985000 ;
        RECT 58.340000  97.985000 74.290000  98.135000 ;
        RECT 58.490000  98.135000 74.290000  98.285000 ;
        RECT 58.640000  98.285000 74.290000  98.435000 ;
        RECT 58.790000  98.435000 74.290000  98.585000 ;
        RECT 58.940000  98.585000 74.290000  98.735000 ;
        RECT 59.090000  98.735000 74.290000  98.885000 ;
        RECT 59.240000  98.885000 74.290000  99.035000 ;
        RECT 59.390000  99.035000 74.290000  99.185000 ;
        RECT 59.540000  99.185000 74.290000  99.335000 ;
        RECT 59.690000  99.335000 74.290000  99.485000 ;
        RECT 59.840000  99.485000 74.290000  99.635000 ;
        RECT 59.990000  99.635000 74.290000  99.785000 ;
        RECT 60.140000  99.785000 74.290000  99.935000 ;
        RECT 60.290000  99.935000 74.290000 100.085000 ;
        RECT 60.440000 100.085000 74.290000 100.235000 ;
        RECT 60.590000 100.235000 74.290000 100.385000 ;
        RECT 60.740000 100.385000 74.290000 100.535000 ;
        RECT 60.890000 100.535000 74.290000 100.685000 ;
        RECT 61.040000 100.685000 74.290000 100.835000 ;
        RECT 61.190000 100.835000 74.290000 100.985000 ;
        RECT 61.340000 100.985000 74.290000 101.135000 ;
        RECT 61.490000 101.135000 74.290000 101.285000 ;
        RECT 61.500000 101.285000 74.290000 101.295000 ;
        RECT 61.500000 101.295000 74.290000 173.320000 ;
    END
  END P_CORE
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT  0.495000   0.000000 24.395000   2.055000 ;
        RECT  0.565000   2.055000 24.395000   2.125000 ;
        RECT  0.635000   2.125000 24.395000   2.195000 ;
        RECT  0.705000   2.195000 24.395000   2.265000 ;
        RECT  0.775000   2.265000 24.395000   2.335000 ;
        RECT  0.845000   2.335000 24.395000   2.405000 ;
        RECT  0.915000   2.405000 24.395000   2.475000 ;
        RECT  0.985000   2.475000 24.395000   2.545000 ;
        RECT  1.005000   2.545000 24.395000   2.565000 ;
        RECT  1.005000   2.565000 24.395000   8.595000 ;
        RECT  1.005000   8.595000 24.395000   8.665000 ;
        RECT  1.005000   8.665000 24.465000   8.735000 ;
        RECT  1.005000   8.735000 24.535000   8.805000 ;
        RECT  1.005000   8.805000 24.605000   8.875000 ;
        RECT  1.005000   8.875000 24.675000   8.945000 ;
        RECT  1.005000   8.945000 24.745000   9.015000 ;
        RECT  1.005000   9.015000 24.815000   9.085000 ;
        RECT  1.005000   9.085000 24.885000   9.155000 ;
        RECT  1.005000   9.155000 24.955000   9.225000 ;
        RECT  1.005000   9.225000 25.025000   9.295000 ;
        RECT  1.005000   9.295000 25.095000   9.365000 ;
        RECT  1.005000   9.365000 25.165000   9.435000 ;
        RECT  1.005000   9.435000 25.235000   9.505000 ;
        RECT  1.005000   9.505000 25.305000   9.575000 ;
        RECT  1.005000   9.575000 25.375000   9.645000 ;
        RECT  1.005000   9.645000 25.445000   9.715000 ;
        RECT  1.005000   9.715000 25.515000   9.785000 ;
        RECT  1.005000   9.785000 25.585000   9.855000 ;
        RECT  1.005000   9.855000 25.655000   9.925000 ;
        RECT  1.005000   9.925000 25.725000   9.995000 ;
        RECT  1.005000   9.995000 25.795000  10.065000 ;
        RECT  1.005000  10.065000 25.865000  10.135000 ;
        RECT  1.005000  10.135000 25.935000  10.205000 ;
        RECT  1.005000  10.205000 26.005000  10.275000 ;
        RECT  1.005000  10.275000 26.075000  10.345000 ;
        RECT  1.005000  10.345000 26.145000  10.415000 ;
        RECT  1.005000  10.415000 26.215000  10.485000 ;
        RECT  1.005000  10.485000 26.285000  10.555000 ;
        RECT  1.005000  10.555000 26.355000  10.625000 ;
        RECT  1.005000  10.625000 26.425000  10.695000 ;
        RECT  1.005000  10.695000 26.495000  10.765000 ;
        RECT  1.005000  10.765000 26.565000  10.835000 ;
        RECT  1.005000  10.835000 26.635000  10.905000 ;
        RECT  1.005000  10.905000 26.705000  10.975000 ;
        RECT  1.005000  10.975000 26.775000  11.045000 ;
        RECT  1.005000  11.045000 26.845000  11.115000 ;
        RECT  1.005000  11.115000 26.915000  11.185000 ;
        RECT  1.005000  11.185000 26.985000  11.255000 ;
        RECT  1.005000  11.255000 27.055000  11.325000 ;
        RECT  1.005000  11.325000 27.125000  11.395000 ;
        RECT  1.005000  11.395000 27.195000  11.465000 ;
        RECT  1.005000  11.465000 27.265000  11.535000 ;
        RECT  1.005000  11.535000 27.335000  11.605000 ;
        RECT  1.005000  11.605000 27.405000  11.675000 ;
        RECT  1.005000  11.675000 27.475000  11.745000 ;
        RECT  1.005000  11.745000 27.545000  11.815000 ;
        RECT  1.005000  11.815000 27.615000  11.885000 ;
        RECT  1.005000  11.885000 27.685000  11.955000 ;
        RECT  1.005000  11.955000 27.755000  12.025000 ;
        RECT  1.005000  12.025000 27.825000  12.095000 ;
        RECT  1.005000  12.095000 27.895000  12.165000 ;
        RECT  1.005000  12.165000 27.965000  12.235000 ;
        RECT  1.005000  12.235000 28.035000  12.305000 ;
        RECT  1.005000  12.305000 28.105000  12.375000 ;
        RECT  1.005000  12.375000 28.175000  12.400000 ;
        RECT  1.005000  12.400000 36.895000  25.700000 ;
        RECT  1.005000  25.700000 18.750000  25.770000 ;
        RECT  1.005000  25.770000 18.680000  25.840000 ;
        RECT  1.005000  25.840000 18.610000  25.910000 ;
        RECT  1.005000  25.910000 18.540000  25.980000 ;
        RECT  1.005000  25.980000 18.470000  26.050000 ;
        RECT  1.005000  26.050000 18.400000  26.120000 ;
        RECT  1.005000  26.120000 18.330000  26.190000 ;
        RECT  1.005000  26.190000 18.260000  26.260000 ;
        RECT  1.005000  26.260000 18.190000  26.330000 ;
        RECT  1.005000  26.330000 18.120000  26.400000 ;
        RECT  1.005000  26.400000 18.050000  26.470000 ;
        RECT  1.005000  26.470000 17.980000  26.540000 ;
        RECT  1.005000  26.540000 17.910000  26.610000 ;
        RECT  1.005000  26.610000 17.840000  26.680000 ;
        RECT  1.005000  26.680000 17.770000  26.750000 ;
        RECT  1.005000  26.750000 17.700000  26.820000 ;
        RECT  1.005000  26.820000 17.630000  26.890000 ;
        RECT  1.005000  26.890000 17.560000  26.960000 ;
        RECT  1.005000  26.960000 17.490000  27.030000 ;
        RECT  1.005000  27.030000 17.420000  27.100000 ;
        RECT  1.005000  27.100000 17.350000  27.170000 ;
        RECT  1.005000  27.170000 17.280000  27.240000 ;
        RECT  1.005000  27.240000 17.210000  27.310000 ;
        RECT  1.005000  27.310000 17.140000  27.380000 ;
        RECT  1.005000  27.380000 17.070000  27.450000 ;
        RECT  1.005000  27.450000 17.000000  27.520000 ;
        RECT  1.005000  27.520000 16.930000  27.590000 ;
        RECT  1.005000  27.590000 16.860000  27.660000 ;
        RECT  1.005000  27.660000 16.790000  27.730000 ;
        RECT  1.005000  27.730000 16.720000  27.800000 ;
        RECT  1.005000  27.800000 16.650000  27.870000 ;
        RECT  1.005000  27.870000 16.580000  27.940000 ;
        RECT  1.005000  27.940000 16.510000  28.010000 ;
        RECT  1.005000  28.010000 16.440000  28.080000 ;
        RECT  1.005000  28.080000 16.370000  28.150000 ;
        RECT  1.005000  28.150000 16.300000  28.220000 ;
        RECT  1.005000  28.220000 16.230000  28.290000 ;
        RECT  1.005000  28.290000 16.160000  28.360000 ;
        RECT  1.005000  28.360000 16.090000  28.430000 ;
        RECT  1.005000  28.430000 16.020000  28.500000 ;
        RECT  1.005000  28.500000 15.950000  28.570000 ;
        RECT  1.005000  28.570000 15.880000  28.640000 ;
        RECT  1.005000  28.640000 15.810000  28.710000 ;
        RECT  1.005000  28.710000 15.740000  28.780000 ;
        RECT  1.005000  28.780000 15.670000  28.850000 ;
        RECT  1.005000  28.850000 15.600000  28.920000 ;
        RECT  1.005000  28.920000 15.530000  28.990000 ;
        RECT  1.005000  28.990000 15.460000  29.060000 ;
        RECT  1.005000  29.060000 15.390000  29.130000 ;
        RECT  1.005000  29.130000 15.320000  29.200000 ;
        RECT  1.005000  29.200000 15.250000  29.270000 ;
        RECT  1.005000  29.270000 15.205000  29.315000 ;
        RECT  1.005000  29.315000 15.205000  35.665000 ;
        RECT  1.005000  35.665000 15.205000  35.735000 ;
        RECT  1.005000  35.735000 15.275000  35.805000 ;
        RECT  1.005000  35.805000 15.345000  35.875000 ;
        RECT  1.005000  35.875000 15.415000  35.945000 ;
        RECT  1.005000  35.945000 15.485000  36.015000 ;
        RECT  1.005000  36.015000 15.555000  36.085000 ;
        RECT  1.005000  36.085000 15.625000  36.155000 ;
        RECT  1.005000  36.155000 15.695000  36.225000 ;
        RECT  1.005000  36.225000 15.765000  36.295000 ;
        RECT  1.005000  36.295000 15.835000  36.365000 ;
        RECT  1.005000  36.365000 15.905000  36.435000 ;
        RECT  1.005000  36.435000 15.975000  36.505000 ;
        RECT  1.005000  36.505000 16.045000  36.575000 ;
        RECT  1.005000  36.575000 16.115000  36.645000 ;
        RECT  1.005000  36.645000 16.185000  36.715000 ;
        RECT  1.005000  36.715000 16.255000  36.785000 ;
        RECT  1.005000  36.785000 16.325000  36.855000 ;
        RECT  1.005000  47.100000 14.120000  54.215000 ;
        RECT  1.005000  54.215000 14.120000  54.285000 ;
        RECT  1.005000  54.285000 14.190000  54.355000 ;
        RECT  1.005000  54.355000 14.260000  54.425000 ;
        RECT  1.005000  54.425000 14.330000  54.495000 ;
        RECT  1.005000  54.495000 14.400000  54.565000 ;
        RECT  1.005000  54.565000 14.470000  54.635000 ;
        RECT  1.005000  54.635000 14.540000  54.705000 ;
        RECT  1.005000  54.705000 14.610000  54.775000 ;
        RECT  1.005000  54.775000 14.680000  54.845000 ;
        RECT  1.005000  54.845000 14.750000  54.915000 ;
        RECT  1.005000  54.915000 14.820000  54.985000 ;
        RECT  1.005000  54.985000 14.890000  55.055000 ;
        RECT  1.005000  55.055000 14.960000  55.125000 ;
        RECT  1.005000  55.125000 15.030000  55.195000 ;
        RECT  1.005000  55.195000 15.100000  55.265000 ;
        RECT  1.005000  55.265000 15.170000  55.335000 ;
        RECT  1.005000  55.335000 15.240000  55.405000 ;
        RECT  1.005000  55.405000 15.310000  55.475000 ;
        RECT  1.005000  55.475000 15.380000  55.545000 ;
        RECT  1.005000  55.545000 15.450000  55.615000 ;
        RECT  1.005000  55.615000 15.520000  55.685000 ;
        RECT  1.005000  55.685000 15.590000  55.755000 ;
        RECT  1.005000  55.755000 15.660000  55.825000 ;
        RECT  1.005000  55.825000 15.730000  55.895000 ;
        RECT  1.005000  55.895000 15.800000  55.965000 ;
        RECT  1.005000  55.965000 15.870000  56.035000 ;
        RECT  1.005000  56.035000 15.940000  56.105000 ;
        RECT  1.005000  56.105000 16.010000  56.175000 ;
        RECT  1.005000  56.175000 16.080000  56.245000 ;
        RECT  1.005000  56.245000 16.150000  56.315000 ;
        RECT  1.005000  56.315000 16.220000  56.385000 ;
        RECT  1.005000  56.385000 16.290000  56.455000 ;
        RECT  1.005000  56.455000 16.360000  56.525000 ;
        RECT  1.005000  56.525000 16.430000  56.595000 ;
        RECT  1.005000  56.595000 16.500000  56.665000 ;
        RECT  1.005000  56.665000 16.570000  56.735000 ;
        RECT  1.005000  56.735000 16.640000  56.805000 ;
        RECT  1.005000  56.805000 16.710000  56.875000 ;
        RECT  1.005000  56.875000 16.780000  56.945000 ;
        RECT  1.005000  56.945000 16.850000  57.015000 ;
        RECT  1.005000  57.015000 16.920000  57.085000 ;
        RECT  1.005000  57.085000 16.990000  57.155000 ;
        RECT  1.005000  57.155000 17.060000  57.225000 ;
        RECT  1.005000  57.225000 17.130000  57.295000 ;
        RECT  1.005000  57.295000 17.200000  57.365000 ;
        RECT  1.005000  57.365000 17.270000  57.435000 ;
        RECT  1.005000  57.435000 17.340000  57.505000 ;
        RECT  1.005000  57.505000 17.410000  57.575000 ;
        RECT  1.005000  57.575000 17.480000  57.645000 ;
        RECT  1.005000  57.645000 17.550000  57.715000 ;
        RECT  1.005000  57.715000 17.620000  57.780000 ;
        RECT  1.005000  57.780000 56.710000  66.480000 ;
        RECT  1.005000  66.480000 17.595000  66.550000 ;
        RECT  1.005000  66.550000 17.525000  66.620000 ;
        RECT  1.005000  66.620000 17.455000  66.690000 ;
        RECT  1.005000  66.690000 17.385000  66.760000 ;
        RECT  1.005000  66.760000 17.315000  66.830000 ;
        RECT  1.005000  66.830000 17.245000  66.900000 ;
        RECT  1.005000  66.900000 17.175000  66.970000 ;
        RECT  1.005000  66.970000 17.105000  67.040000 ;
        RECT  1.005000  67.040000 17.035000  67.110000 ;
        RECT  1.005000  67.110000 16.965000  67.180000 ;
        RECT  1.005000  67.180000 16.895000  67.250000 ;
        RECT  1.005000  67.250000 16.825000  67.320000 ;
        RECT  1.005000  67.320000 16.755000  67.390000 ;
        RECT  1.005000  67.390000 16.685000  67.460000 ;
        RECT  1.005000  67.460000 16.615000  67.530000 ;
        RECT  1.005000  67.530000 16.545000  67.600000 ;
        RECT  1.005000  67.600000 16.475000  67.670000 ;
        RECT  1.005000  67.670000 16.405000  67.740000 ;
        RECT  1.005000  67.740000 16.335000  67.810000 ;
        RECT  1.005000  67.810000 16.265000  67.880000 ;
        RECT  1.005000  67.880000 16.195000  67.950000 ;
        RECT  1.005000  67.950000 16.125000  68.020000 ;
        RECT  1.005000  68.020000 16.055000  68.090000 ;
        RECT  1.005000  68.090000 15.985000  68.160000 ;
        RECT  1.005000  68.160000 15.915000  68.230000 ;
        RECT  1.005000  68.230000 15.845000  68.300000 ;
        RECT  1.005000  68.300000 15.775000  68.370000 ;
        RECT  1.005000  68.370000 15.705000  68.440000 ;
        RECT  1.005000  68.440000 15.635000  68.510000 ;
        RECT  1.005000  68.510000 15.565000  68.580000 ;
        RECT  1.005000  68.580000 15.495000  68.650000 ;
        RECT  1.005000  68.650000 15.425000  68.720000 ;
        RECT  1.005000  68.720000 15.355000  68.790000 ;
        RECT  1.005000  68.790000 15.285000  68.860000 ;
        RECT  1.005000  68.860000 15.215000  68.930000 ;
        RECT  1.005000  68.930000 15.145000  69.000000 ;
        RECT  1.005000  69.000000 15.075000  69.070000 ;
        RECT  1.005000  69.070000 15.005000  69.140000 ;
        RECT  1.005000  69.140000 14.935000  69.210000 ;
        RECT  1.005000  69.210000 14.865000  69.280000 ;
        RECT  1.005000  69.280000 14.795000  69.350000 ;
        RECT  1.005000  69.350000 14.725000  69.420000 ;
        RECT  1.005000  69.420000 14.655000  69.490000 ;
        RECT  1.005000  69.490000 14.585000  69.560000 ;
        RECT  1.005000  69.560000 14.515000  69.630000 ;
        RECT  1.005000  69.630000 14.445000  69.700000 ;
        RECT  1.005000  69.700000 14.375000  69.770000 ;
        RECT  1.005000  69.770000 14.305000  69.840000 ;
        RECT  1.005000  69.840000 14.235000  69.910000 ;
        RECT  1.005000  69.910000 14.165000  69.980000 ;
        RECT  1.005000  69.980000 14.120000  70.025000 ;
        RECT  1.005000  70.025000 14.120000  77.240000 ;
        RECT  1.005000  77.240000 14.120000  77.310000 ;
        RECT  1.005000  77.310000 14.190000  77.380000 ;
        RECT  1.005000  77.380000 14.260000  77.450000 ;
        RECT  1.005000  77.450000 14.330000  77.520000 ;
        RECT  1.005000  77.520000 14.400000  77.590000 ;
        RECT  1.005000  77.590000 14.470000  77.660000 ;
        RECT  1.005000  77.660000 14.540000  77.730000 ;
        RECT  1.005000  77.730000 14.610000  77.800000 ;
        RECT  1.005000  77.800000 14.680000  77.870000 ;
        RECT  1.005000  77.870000 14.750000  77.940000 ;
        RECT  1.005000  77.940000 14.820000  78.010000 ;
        RECT  1.005000  78.010000 14.890000  78.080000 ;
        RECT  1.005000  78.080000 14.960000  78.150000 ;
        RECT  1.005000  78.150000 15.030000  78.220000 ;
        RECT  1.005000  78.220000 15.100000  78.290000 ;
        RECT  1.005000  78.290000 15.170000  78.360000 ;
        RECT  1.005000  78.360000 15.240000  78.430000 ;
        RECT  1.005000  78.430000 15.310000  78.500000 ;
        RECT  1.005000  78.500000 15.380000  78.570000 ;
        RECT  1.005000  78.570000 15.450000  78.640000 ;
        RECT  1.005000  78.640000 15.520000  78.710000 ;
        RECT  1.005000  78.710000 15.590000  78.780000 ;
        RECT  1.005000  78.780000 15.660000  78.850000 ;
        RECT  1.005000  78.850000 15.730000  78.920000 ;
        RECT  1.005000  78.920000 15.800000  78.990000 ;
        RECT  1.005000  78.990000 15.870000  79.060000 ;
        RECT  1.005000  79.060000 15.940000  79.130000 ;
        RECT  1.005000  79.130000 16.010000  79.200000 ;
        RECT  1.005000  79.200000 16.080000  79.270000 ;
        RECT  1.005000  79.270000 16.150000  79.340000 ;
        RECT  1.005000  79.340000 16.220000  79.410000 ;
        RECT  1.005000  79.410000 16.290000  79.480000 ;
        RECT  1.005000  79.480000 16.360000  79.550000 ;
        RECT  1.005000  79.550000 16.430000  79.620000 ;
        RECT  1.005000  79.620000 16.500000  79.690000 ;
        RECT  1.005000  79.690000 16.570000  79.760000 ;
        RECT  1.005000  79.760000 16.640000  79.830000 ;
        RECT  1.005000  79.830000 16.710000  79.900000 ;
        RECT  1.005000  79.900000 16.780000  79.970000 ;
        RECT  1.005000  79.970000 16.850000  80.040000 ;
        RECT  1.005000  80.040000 16.920000  80.110000 ;
        RECT  1.005000  80.110000 16.990000  80.180000 ;
        RECT  1.005000  80.180000 17.060000  80.250000 ;
        RECT  1.005000  80.250000 17.130000  80.320000 ;
        RECT  1.005000  80.320000 17.200000  80.390000 ;
        RECT  1.005000  80.390000 17.270000  80.460000 ;
        RECT  1.005000  80.460000 17.340000  80.530000 ;
        RECT  1.005000  80.530000 17.410000  80.600000 ;
        RECT  1.005000  80.600000 17.480000  80.670000 ;
        RECT  1.005000  80.670000 17.550000  80.740000 ;
        RECT  1.005000  80.740000 17.620000  80.780000 ;
        RECT  1.005000  80.780000 56.705000  89.480000 ;
        RECT  1.005000  89.480000 17.595000  89.550000 ;
        RECT  1.005000  89.550000 17.525000  89.620000 ;
        RECT  1.005000  89.620000 17.455000  89.690000 ;
        RECT  1.005000  89.690000 17.385000  89.760000 ;
        RECT  1.005000  89.760000 17.315000  89.830000 ;
        RECT  1.005000  89.830000 17.245000  89.900000 ;
        RECT  1.005000  89.900000 17.175000  89.970000 ;
        RECT  1.005000  89.970000 17.105000  90.040000 ;
        RECT  1.005000  90.040000 17.035000  90.110000 ;
        RECT  1.005000  90.110000 16.965000  90.180000 ;
        RECT  1.005000  90.180000 16.895000  90.250000 ;
        RECT  1.005000  90.250000 16.825000  90.320000 ;
        RECT  1.005000  90.320000 16.755000  90.390000 ;
        RECT  1.005000  90.390000 16.685000  90.460000 ;
        RECT  1.005000  90.460000 16.615000  90.530000 ;
        RECT  1.005000  90.530000 16.545000  90.600000 ;
        RECT  1.005000  90.600000 16.475000  90.670000 ;
        RECT  1.005000  90.670000 16.405000  90.740000 ;
        RECT  1.005000  90.740000 16.335000  90.810000 ;
        RECT  1.005000  90.810000 16.265000  90.880000 ;
        RECT  1.005000  90.880000 16.195000  90.950000 ;
        RECT  1.005000  90.950000 16.125000  91.020000 ;
        RECT  1.005000  91.020000 16.055000  91.090000 ;
        RECT  1.005000  91.090000 15.985000  91.160000 ;
        RECT  1.005000  91.160000 15.915000  91.230000 ;
        RECT  1.005000  91.230000 15.845000  91.300000 ;
        RECT  1.005000  91.300000 15.775000  91.370000 ;
        RECT  1.005000  91.370000 15.705000  91.440000 ;
        RECT  1.005000  91.440000 15.635000  91.510000 ;
        RECT  1.005000  91.510000 15.565000  91.580000 ;
        RECT  1.005000  91.580000 15.495000  91.650000 ;
        RECT  1.005000  91.650000 15.425000  91.720000 ;
        RECT  1.005000  91.720000 15.355000  91.790000 ;
        RECT  1.005000  91.790000 15.285000  91.860000 ;
        RECT  1.005000  91.860000 15.215000  91.930000 ;
        RECT  1.005000  91.930000 15.145000  92.000000 ;
        RECT  1.005000  92.000000 15.075000  92.070000 ;
        RECT  1.005000  92.070000 15.005000  92.140000 ;
        RECT  1.005000  92.140000 14.935000  92.210000 ;
        RECT  1.005000  92.210000 14.865000  92.280000 ;
        RECT  1.005000  92.280000 14.795000  92.350000 ;
        RECT  1.005000  92.350000 14.725000  92.420000 ;
        RECT  1.005000  92.420000 14.655000  92.490000 ;
        RECT  1.005000  92.490000 14.585000  92.560000 ;
        RECT  1.005000  92.560000 14.515000  92.630000 ;
        RECT  1.005000  92.630000 14.445000  92.700000 ;
        RECT  1.005000  92.700000 14.375000  92.770000 ;
        RECT  1.005000  92.770000 14.305000  92.840000 ;
        RECT  1.005000  92.840000 14.235000  92.910000 ;
        RECT  1.005000  92.910000 14.165000  92.980000 ;
        RECT  1.005000  92.980000 14.120000  93.025000 ;
        RECT  1.005000  93.025000 14.120000 100.240000 ;
        RECT  1.005000 100.240000 14.120000 100.310000 ;
        RECT  1.005000 100.310000 14.190000 100.380000 ;
        RECT  1.005000 100.380000 14.260000 100.450000 ;
        RECT  1.005000 100.450000 14.330000 100.520000 ;
        RECT  1.005000 100.520000 14.400000 100.590000 ;
        RECT  1.005000 100.590000 14.470000 100.660000 ;
        RECT  1.005000 100.660000 14.540000 100.730000 ;
        RECT  1.005000 100.730000 14.610000 100.800000 ;
        RECT  1.005000 100.800000 14.680000 100.870000 ;
        RECT  1.005000 100.870000 14.750000 100.940000 ;
        RECT  1.005000 100.940000 14.820000 101.010000 ;
        RECT  1.005000 101.010000 14.890000 101.080000 ;
        RECT  1.005000 101.080000 14.960000 101.150000 ;
        RECT  1.005000 101.150000 15.030000 101.220000 ;
        RECT  1.005000 101.220000 15.100000 101.290000 ;
        RECT  1.005000 101.290000 15.170000 101.360000 ;
        RECT  1.005000 101.360000 15.240000 101.430000 ;
        RECT  1.005000 101.430000 15.310000 101.500000 ;
        RECT  1.005000 101.500000 15.380000 101.570000 ;
        RECT  1.005000 101.570000 15.450000 101.640000 ;
        RECT  1.005000 101.640000 15.520000 101.710000 ;
        RECT  1.005000 101.710000 15.590000 101.780000 ;
        RECT  1.005000 101.780000 15.660000 101.850000 ;
        RECT  1.005000 101.850000 15.730000 101.920000 ;
        RECT  1.005000 101.920000 15.800000 101.990000 ;
        RECT  1.005000 101.990000 15.870000 102.060000 ;
        RECT  1.005000 102.060000 15.940000 102.130000 ;
        RECT  1.005000 102.130000 16.010000 102.200000 ;
        RECT  1.005000 102.200000 16.080000 102.270000 ;
        RECT  1.005000 102.270000 16.150000 102.340000 ;
        RECT  1.005000 102.340000 16.220000 102.410000 ;
        RECT  1.005000 102.410000 16.290000 102.480000 ;
        RECT  1.005000 102.480000 16.360000 102.550000 ;
        RECT  1.005000 102.550000 16.430000 102.620000 ;
        RECT  1.005000 102.620000 16.500000 102.690000 ;
        RECT  1.005000 102.690000 16.570000 102.760000 ;
        RECT  1.005000 102.760000 16.640000 102.830000 ;
        RECT  1.005000 102.830000 16.710000 102.900000 ;
        RECT  1.005000 102.900000 16.780000 102.970000 ;
        RECT  1.005000 102.970000 16.850000 103.040000 ;
        RECT  1.005000 103.040000 16.920000 103.110000 ;
        RECT  1.005000 103.110000 16.990000 103.180000 ;
        RECT  1.005000 103.180000 17.060000 103.250000 ;
        RECT  1.005000 103.250000 17.130000 103.320000 ;
        RECT  1.005000 103.320000 17.200000 103.390000 ;
        RECT  1.005000 103.390000 17.270000 103.460000 ;
        RECT  1.005000 103.460000 17.340000 103.530000 ;
        RECT  1.005000 103.530000 17.410000 103.600000 ;
        RECT  1.005000 103.600000 17.480000 103.670000 ;
        RECT  1.005000 103.670000 17.550000 103.740000 ;
        RECT  1.005000 103.740000 17.620000 103.780000 ;
        RECT  1.005000 103.780000 56.705000 112.480000 ;
        RECT  1.005000 112.480000 17.635000 112.550000 ;
        RECT  1.005000 112.550000 17.565000 112.620000 ;
        RECT  1.005000 112.620000 17.495000 112.690000 ;
        RECT  1.005000 112.690000 17.425000 112.760000 ;
        RECT  1.005000 112.760000 17.355000 112.830000 ;
        RECT  1.005000 112.830000 17.285000 112.900000 ;
        RECT  1.005000 112.900000 17.215000 112.970000 ;
        RECT  1.005000 112.970000 17.145000 113.040000 ;
        RECT  1.005000 113.040000 17.075000 113.110000 ;
        RECT  1.005000 113.110000 17.005000 113.180000 ;
        RECT  1.005000 113.180000 16.935000 113.250000 ;
        RECT  1.005000 113.250000 16.865000 113.320000 ;
        RECT  1.005000 113.320000 16.795000 113.390000 ;
        RECT  1.005000 113.390000 16.725000 113.460000 ;
        RECT  1.005000 113.460000 16.655000 113.530000 ;
        RECT  1.005000 113.530000 16.585000 113.600000 ;
        RECT  1.005000 113.600000 16.515000 113.670000 ;
        RECT  1.005000 113.670000 16.445000 113.740000 ;
        RECT  1.005000 113.740000 16.375000 113.810000 ;
        RECT  1.005000 113.810000 16.305000 113.880000 ;
        RECT  1.005000 113.880000 16.235000 113.950000 ;
        RECT  1.005000 113.950000 16.165000 114.020000 ;
        RECT  1.005000 114.020000 16.095000 114.090000 ;
        RECT  1.005000 114.090000 16.025000 114.160000 ;
        RECT  1.005000 114.160000 15.955000 114.230000 ;
        RECT  1.005000 114.230000 15.885000 114.300000 ;
        RECT  1.005000 114.300000 15.815000 114.370000 ;
        RECT  1.005000 114.370000 15.745000 114.440000 ;
        RECT  1.005000 114.440000 15.675000 114.510000 ;
        RECT  1.005000 114.510000 15.605000 114.580000 ;
        RECT  1.005000 114.580000 15.535000 114.650000 ;
        RECT  1.005000 114.650000 15.465000 114.720000 ;
        RECT  1.005000 114.720000 15.395000 114.790000 ;
        RECT  1.005000 114.790000 15.325000 114.860000 ;
        RECT  1.005000 114.860000 15.255000 114.930000 ;
        RECT  1.005000 114.930000 15.185000 115.000000 ;
        RECT  1.005000 115.000000 15.115000 115.070000 ;
        RECT  1.005000 115.070000 15.045000 115.140000 ;
        RECT  1.005000 115.140000 14.975000 115.210000 ;
        RECT  1.005000 115.210000 14.905000 115.280000 ;
        RECT  1.005000 115.280000 14.835000 115.350000 ;
        RECT  1.005000 115.350000 14.765000 115.420000 ;
        RECT  1.005000 115.420000 14.695000 115.490000 ;
        RECT  1.005000 115.490000 14.625000 115.560000 ;
        RECT  1.005000 115.560000 14.555000 115.630000 ;
        RECT  1.005000 115.630000 14.485000 115.700000 ;
        RECT  1.005000 115.700000 14.415000 115.770000 ;
        RECT  1.005000 115.770000 14.345000 115.840000 ;
        RECT  1.005000 115.840000 14.275000 115.910000 ;
        RECT  1.005000 115.910000 14.205000 115.980000 ;
        RECT  1.005000 115.980000 14.135000 116.050000 ;
        RECT  1.005000 116.050000 14.120000 116.065000 ;
        RECT  1.005000 116.065000 14.120000 123.145000 ;
        RECT  1.005000 123.145000 14.120000 123.215000 ;
        RECT  1.005000 123.215000 14.190000 123.285000 ;
        RECT  1.005000 123.285000 14.260000 123.355000 ;
        RECT  1.005000 123.355000 14.330000 123.425000 ;
        RECT  1.005000 123.425000 14.400000 123.495000 ;
        RECT  1.005000 123.495000 14.470000 123.565000 ;
        RECT  1.005000 123.565000 14.540000 123.635000 ;
        RECT  1.005000 123.635000 14.610000 123.705000 ;
        RECT  1.005000 123.705000 14.680000 123.775000 ;
        RECT  1.005000 123.775000 14.750000 123.845000 ;
        RECT  1.005000 123.845000 14.820000 123.915000 ;
        RECT  1.005000 123.915000 14.890000 123.985000 ;
        RECT  1.005000 123.985000 14.960000 124.055000 ;
        RECT  1.005000 124.055000 15.030000 124.125000 ;
        RECT  1.005000 124.125000 15.100000 124.195000 ;
        RECT  1.005000 124.195000 15.170000 124.265000 ;
        RECT  1.005000 124.265000 15.240000 124.335000 ;
        RECT  1.005000 124.335000 15.310000 124.405000 ;
        RECT  1.005000 124.405000 15.380000 124.475000 ;
        RECT  1.005000 124.475000 15.450000 124.545000 ;
        RECT  1.005000 124.545000 15.520000 124.615000 ;
        RECT  1.005000 124.615000 15.590000 124.685000 ;
        RECT  1.005000 124.685000 15.660000 124.755000 ;
        RECT  1.005000 124.755000 15.730000 124.825000 ;
        RECT  1.005000 124.825000 15.800000 124.895000 ;
        RECT  1.005000 124.895000 15.870000 124.965000 ;
        RECT  1.005000 124.965000 15.940000 125.035000 ;
        RECT  1.005000 125.035000 16.010000 125.105000 ;
        RECT  1.005000 125.105000 16.080000 125.175000 ;
        RECT  1.005000 125.175000 16.150000 125.245000 ;
        RECT  1.005000 125.245000 16.220000 125.315000 ;
        RECT  1.005000 125.315000 16.290000 125.385000 ;
        RECT  1.005000 125.385000 16.360000 125.455000 ;
        RECT  1.005000 125.455000 16.430000 125.525000 ;
        RECT  1.005000 125.525000 16.500000 125.595000 ;
        RECT  1.005000 125.595000 16.570000 125.665000 ;
        RECT  1.005000 125.665000 16.640000 125.735000 ;
        RECT  1.005000 125.735000 16.710000 125.805000 ;
        RECT  1.005000 125.805000 16.780000 125.875000 ;
        RECT  1.005000 125.875000 16.850000 125.945000 ;
        RECT  1.005000 125.945000 16.920000 126.015000 ;
        RECT  1.005000 126.015000 16.990000 126.085000 ;
        RECT  1.005000 126.085000 17.060000 126.155000 ;
        RECT  1.005000 126.155000 17.130000 126.225000 ;
        RECT  1.005000 126.225000 17.200000 126.295000 ;
        RECT  1.005000 126.295000 17.270000 126.365000 ;
        RECT  1.005000 126.365000 17.340000 126.435000 ;
        RECT  1.005000 126.435000 17.410000 126.505000 ;
        RECT  1.005000 126.505000 17.480000 126.575000 ;
        RECT  1.005000 126.575000 17.550000 126.645000 ;
        RECT  1.005000 126.645000 17.620000 126.715000 ;
        RECT  1.005000 126.715000 17.690000 126.780000 ;
        RECT  1.005000 126.780000 56.705000 135.480000 ;
        RECT  1.005000 135.480000 17.740000 135.550000 ;
        RECT  1.005000 135.550000 17.670000 135.620000 ;
        RECT  1.005000 135.620000 17.600000 135.690000 ;
        RECT  1.005000 135.690000 17.530000 135.760000 ;
        RECT  1.005000 135.760000 17.460000 135.830000 ;
        RECT  1.005000 135.830000 17.390000 135.900000 ;
        RECT  1.005000 135.900000 17.320000 135.970000 ;
        RECT  1.005000 135.970000 17.250000 136.040000 ;
        RECT  1.005000 136.040000 17.180000 136.110000 ;
        RECT  1.005000 136.110000 17.110000 136.180000 ;
        RECT  1.005000 136.180000 17.040000 136.250000 ;
        RECT  1.005000 136.250000 16.970000 136.320000 ;
        RECT  1.005000 136.320000 16.900000 136.390000 ;
        RECT  1.005000 136.390000 16.830000 136.460000 ;
        RECT  1.005000 136.460000 16.760000 136.530000 ;
        RECT  1.005000 136.530000 16.690000 136.600000 ;
        RECT  1.005000 136.600000 16.620000 136.670000 ;
        RECT  1.005000 136.670000 16.550000 136.740000 ;
        RECT  1.005000 136.740000 16.480000 136.810000 ;
        RECT  1.005000 136.810000 16.410000 136.880000 ;
        RECT  1.005000 136.880000 16.340000 136.950000 ;
        RECT  1.005000 136.950000 16.270000 137.020000 ;
        RECT  1.005000 137.020000 16.200000 137.090000 ;
        RECT  1.005000 137.090000 16.130000 137.160000 ;
        RECT  1.005000 137.160000 16.060000 137.230000 ;
        RECT  1.005000 137.230000 15.990000 137.300000 ;
        RECT  1.005000 137.300000 15.920000 137.370000 ;
        RECT  1.005000 137.370000 15.850000 137.440000 ;
        RECT  1.005000 137.440000 15.780000 137.510000 ;
        RECT  1.005000 137.510000 15.710000 137.580000 ;
        RECT  1.005000 137.580000 15.640000 137.650000 ;
        RECT  1.005000 137.650000 15.570000 137.720000 ;
        RECT  1.005000 137.720000 15.500000 137.790000 ;
        RECT  1.005000 137.790000 15.430000 137.860000 ;
        RECT  1.005000 137.860000 15.360000 137.930000 ;
        RECT  1.005000 137.930000 15.290000 138.000000 ;
        RECT  1.005000 138.000000 15.220000 138.070000 ;
        RECT  1.005000 138.070000 15.150000 138.140000 ;
        RECT  1.005000 138.140000 15.080000 138.210000 ;
        RECT  1.005000 138.210000 15.010000 138.280000 ;
        RECT  1.005000 138.280000 14.940000 138.350000 ;
        RECT  1.005000 138.350000 14.870000 138.420000 ;
        RECT  1.005000 138.420000 14.800000 138.490000 ;
        RECT  1.005000 138.490000 14.730000 138.560000 ;
        RECT  1.005000 138.560000 14.660000 138.630000 ;
        RECT  1.005000 138.630000 14.590000 138.700000 ;
        RECT  1.005000 138.700000 14.520000 138.770000 ;
        RECT  1.005000 138.770000 14.450000 138.840000 ;
        RECT  1.005000 138.840000 14.380000 138.910000 ;
        RECT  1.005000 138.910000 14.310000 138.980000 ;
        RECT  1.005000 138.980000 14.240000 139.050000 ;
        RECT  1.005000 139.050000 14.170000 139.120000 ;
        RECT  1.005000 139.120000 14.120000 139.170000 ;
        RECT  1.005000 139.170000 14.120000 146.215000 ;
        RECT  1.005000 146.215000 14.120000 146.285000 ;
        RECT  1.005000 146.285000 14.190000 146.355000 ;
        RECT  1.005000 146.355000 14.260000 146.425000 ;
        RECT  1.005000 146.425000 14.330000 146.495000 ;
        RECT  1.005000 146.495000 14.400000 146.565000 ;
        RECT  1.005000 146.565000 14.470000 146.635000 ;
        RECT  1.005000 146.635000 14.540000 146.705000 ;
        RECT  1.005000 146.705000 14.610000 146.775000 ;
        RECT  1.005000 146.775000 14.680000 146.845000 ;
        RECT  1.005000 146.845000 14.750000 146.915000 ;
        RECT  1.005000 146.915000 14.820000 146.985000 ;
        RECT  1.005000 146.985000 14.890000 147.055000 ;
        RECT  1.005000 147.055000 14.960000 147.125000 ;
        RECT  1.005000 147.125000 15.030000 147.195000 ;
        RECT  1.005000 147.195000 15.100000 147.265000 ;
        RECT  1.005000 147.265000 15.170000 147.335000 ;
        RECT  1.005000 147.335000 15.240000 147.405000 ;
        RECT  1.005000 147.405000 15.310000 147.475000 ;
        RECT  1.005000 147.475000 15.380000 147.545000 ;
        RECT  1.005000 147.545000 15.450000 147.615000 ;
        RECT  1.005000 147.615000 15.520000 147.685000 ;
        RECT  1.005000 147.685000 15.590000 147.755000 ;
        RECT  1.005000 147.755000 15.660000 147.825000 ;
        RECT  1.005000 147.825000 15.730000 147.895000 ;
        RECT  1.005000 147.895000 15.800000 147.965000 ;
        RECT  1.005000 147.965000 15.870000 148.035000 ;
        RECT  1.005000 148.035000 15.940000 148.105000 ;
        RECT  1.005000 148.105000 16.010000 148.175000 ;
        RECT  1.005000 148.175000 16.080000 148.245000 ;
        RECT  1.005000 148.245000 16.150000 148.315000 ;
        RECT  1.005000 148.315000 16.220000 148.385000 ;
        RECT  1.005000 148.385000 16.290000 148.455000 ;
        RECT  1.005000 148.455000 16.360000 148.525000 ;
        RECT  1.005000 148.525000 16.430000 148.595000 ;
        RECT  1.005000 148.595000 16.500000 148.665000 ;
        RECT  1.005000 148.665000 16.570000 148.735000 ;
        RECT  1.005000 148.735000 16.640000 148.805000 ;
        RECT  1.005000 148.805000 16.710000 148.875000 ;
        RECT  1.005000 148.875000 16.780000 148.945000 ;
        RECT  1.005000 148.945000 16.850000 149.015000 ;
        RECT  1.005000 149.015000 16.920000 149.085000 ;
        RECT  1.005000 149.085000 16.990000 149.155000 ;
        RECT  1.005000 149.155000 17.060000 149.225000 ;
        RECT  1.005000 149.225000 17.130000 149.295000 ;
        RECT  1.005000 149.295000 17.200000 149.365000 ;
        RECT  1.005000 149.365000 17.270000 149.435000 ;
        RECT  1.005000 149.435000 17.340000 149.505000 ;
        RECT  1.005000 149.505000 17.410000 149.575000 ;
        RECT  1.005000 149.575000 17.480000 149.645000 ;
        RECT  1.005000 149.645000 17.550000 149.715000 ;
        RECT  1.005000 149.715000 17.620000 149.780000 ;
        RECT  1.005000 149.780000 56.705000 158.480000 ;
        RECT  1.005000 158.480000 17.650000 158.550000 ;
        RECT  1.005000 158.550000 17.580000 158.620000 ;
        RECT  1.005000 158.620000 17.510000 158.690000 ;
        RECT  1.005000 158.690000 17.440000 158.760000 ;
        RECT  1.005000 158.760000 17.370000 158.830000 ;
        RECT  1.005000 158.830000 17.300000 158.900000 ;
        RECT  1.005000 158.900000 17.230000 158.970000 ;
        RECT  1.005000 158.970000 17.160000 159.040000 ;
        RECT  1.005000 159.040000 17.090000 159.110000 ;
        RECT  1.005000 159.110000 17.020000 159.180000 ;
        RECT  1.005000 159.180000 16.950000 159.250000 ;
        RECT  1.005000 159.250000 16.880000 159.320000 ;
        RECT  1.005000 159.320000 16.810000 159.390000 ;
        RECT  1.005000 159.390000 16.740000 159.460000 ;
        RECT  1.005000 159.460000 16.670000 159.530000 ;
        RECT  1.005000 159.530000 16.600000 159.600000 ;
        RECT  1.005000 159.600000 16.530000 159.670000 ;
        RECT  1.005000 159.670000 16.460000 159.740000 ;
        RECT  1.005000 159.740000 16.390000 159.810000 ;
        RECT  1.005000 159.810000 16.320000 159.880000 ;
        RECT  1.005000 159.880000 16.250000 159.950000 ;
        RECT  1.005000 159.950000 16.180000 160.020000 ;
        RECT  1.005000 160.020000 16.110000 160.090000 ;
        RECT  1.005000 160.090000 16.040000 160.160000 ;
        RECT  1.005000 160.160000 15.970000 160.230000 ;
        RECT  1.005000 160.230000 15.900000 160.300000 ;
        RECT  1.005000 160.300000 15.830000 160.370000 ;
        RECT  1.005000 160.370000 15.760000 160.440000 ;
        RECT  1.005000 160.440000 15.690000 160.510000 ;
        RECT  1.005000 160.510000 15.620000 160.580000 ;
        RECT  1.005000 160.580000 15.550000 160.650000 ;
        RECT  1.005000 160.650000 15.480000 160.720000 ;
        RECT  1.005000 160.720000 15.410000 160.790000 ;
        RECT  1.005000 160.790000 15.340000 160.860000 ;
        RECT  1.005000 160.860000 15.270000 160.930000 ;
        RECT  1.005000 160.930000 15.200000 161.000000 ;
        RECT  1.005000 161.000000 15.130000 161.070000 ;
        RECT  1.005000 161.070000 15.060000 161.140000 ;
        RECT  1.005000 161.140000 14.990000 161.210000 ;
        RECT  1.005000 161.210000 14.920000 161.280000 ;
        RECT  1.005000 161.280000 14.850000 161.350000 ;
        RECT  1.005000 161.350000 14.780000 161.420000 ;
        RECT  1.005000 161.420000 14.710000 161.490000 ;
        RECT  1.005000 161.490000 14.640000 161.560000 ;
        RECT  1.005000 161.560000 14.570000 161.630000 ;
        RECT  1.005000 161.630000 14.500000 161.700000 ;
        RECT  1.005000 161.700000 14.430000 161.770000 ;
        RECT  1.005000 161.770000 14.360000 161.840000 ;
        RECT  1.005000 161.840000 14.290000 161.910000 ;
        RECT  1.005000 161.910000 14.220000 161.980000 ;
        RECT  1.005000 161.980000 14.150000 162.050000 ;
        RECT  1.005000 162.050000 14.120000 162.080000 ;
        RECT  1.005000 162.080000 14.120000 169.220000 ;
        RECT  1.005000 169.220000 14.120000 169.290000 ;
        RECT  1.005000 169.290000 14.190000 169.360000 ;
        RECT  1.005000 169.360000 14.260000 169.430000 ;
        RECT  1.005000 169.430000 14.330000 169.500000 ;
        RECT  1.005000 169.500000 14.400000 169.570000 ;
        RECT  1.005000 169.570000 14.470000 169.640000 ;
        RECT  1.005000 169.640000 14.540000 169.710000 ;
        RECT  1.005000 169.710000 14.610000 169.780000 ;
        RECT  1.005000 169.780000 14.680000 169.850000 ;
        RECT  1.005000 169.850000 14.750000 169.920000 ;
        RECT  1.005000 169.920000 14.820000 169.990000 ;
        RECT  1.005000 169.990000 14.890000 170.060000 ;
        RECT  1.005000 170.060000 14.960000 170.130000 ;
        RECT  1.005000 170.130000 15.030000 170.200000 ;
        RECT  1.005000 170.200000 15.100000 170.270000 ;
        RECT  1.005000 170.270000 15.170000 170.340000 ;
        RECT  1.005000 170.340000 15.240000 170.410000 ;
        RECT  1.005000 170.410000 15.310000 170.480000 ;
        RECT  1.005000 170.480000 15.380000 170.550000 ;
        RECT  1.005000 170.550000 15.450000 170.620000 ;
        RECT  1.005000 170.620000 15.520000 170.690000 ;
        RECT  1.005000 170.690000 15.590000 170.760000 ;
        RECT  1.005000 170.760000 15.660000 170.830000 ;
        RECT  1.005000 170.830000 15.730000 170.900000 ;
        RECT  1.005000 170.900000 15.800000 170.970000 ;
        RECT  1.005000 170.970000 15.870000 171.040000 ;
        RECT  1.005000 171.040000 15.940000 171.110000 ;
        RECT  1.005000 171.110000 16.010000 171.180000 ;
        RECT  1.005000 171.180000 16.080000 171.250000 ;
        RECT  1.005000 171.250000 16.150000 171.320000 ;
        RECT  1.005000 171.320000 16.220000 171.390000 ;
        RECT  1.005000 171.390000 16.290000 171.460000 ;
        RECT  1.005000 171.460000 16.360000 171.530000 ;
        RECT  1.005000 171.530000 16.430000 171.600000 ;
        RECT  1.005000 171.600000 16.500000 171.670000 ;
        RECT  1.005000 171.670000 16.570000 171.740000 ;
        RECT  1.005000 171.740000 16.640000 171.810000 ;
        RECT  1.005000 171.810000 16.710000 171.880000 ;
        RECT  1.005000 171.880000 16.780000 171.950000 ;
        RECT  1.005000 171.950000 16.850000 172.020000 ;
        RECT  1.005000 172.020000 16.920000 172.090000 ;
        RECT  1.005000 172.090000 16.990000 172.160000 ;
        RECT  1.005000 172.160000 17.060000 172.230000 ;
        RECT  1.005000 172.230000 17.130000 172.300000 ;
        RECT  1.005000 172.300000 17.200000 172.370000 ;
        RECT  1.005000 172.370000 17.270000 172.440000 ;
        RECT  1.005000 172.440000 17.340000 172.510000 ;
        RECT  1.005000 172.510000 17.410000 172.580000 ;
        RECT  1.005000 172.580000 17.480000 172.650000 ;
        RECT  1.005000 172.650000 17.550000 172.720000 ;
        RECT  1.005000 172.720000 17.620000 172.780000 ;
        RECT  1.005000 172.780000 57.960000 181.480000 ;
        RECT  1.005000 181.480000 17.625000 181.550000 ;
        RECT  1.005000 181.550000 17.555000 181.620000 ;
        RECT  1.005000 181.620000 17.485000 181.690000 ;
        RECT  1.005000 181.690000 17.415000 181.760000 ;
        RECT  1.005000 181.760000 17.345000 181.830000 ;
        RECT  1.005000 181.830000 17.275000 181.900000 ;
        RECT  1.005000 181.900000 17.205000 181.970000 ;
        RECT  1.005000 181.970000 17.135000 182.040000 ;
        RECT  1.005000 182.040000 17.065000 182.110000 ;
        RECT  1.005000 182.110000 16.995000 182.180000 ;
        RECT  1.005000 182.180000 16.925000 182.250000 ;
        RECT  1.005000 182.250000 16.855000 182.320000 ;
        RECT  1.005000 182.320000 16.785000 182.390000 ;
        RECT  1.005000 182.390000 16.715000 182.460000 ;
        RECT  1.005000 182.460000 16.645000 182.530000 ;
        RECT  1.005000 182.530000 16.575000 182.600000 ;
        RECT  1.005000 182.600000 16.505000 182.670000 ;
        RECT  1.005000 182.670000 16.435000 182.740000 ;
        RECT  1.005000 182.740000 16.365000 182.810000 ;
        RECT  1.005000 182.810000 16.295000 182.880000 ;
        RECT  1.005000 182.880000 16.225000 182.950000 ;
        RECT  1.005000 182.950000 16.155000 183.020000 ;
        RECT  1.005000 183.020000 16.085000 183.090000 ;
        RECT  1.005000 183.090000 16.015000 183.160000 ;
        RECT  1.005000 183.160000 15.945000 183.230000 ;
        RECT  1.005000 183.230000 15.875000 183.300000 ;
        RECT  1.005000 183.300000 15.805000 183.370000 ;
        RECT  1.005000 183.370000 15.735000 183.440000 ;
        RECT  1.005000 183.440000 15.665000 183.510000 ;
        RECT  1.005000 183.510000 15.595000 183.580000 ;
        RECT  1.005000 183.580000 15.525000 183.650000 ;
        RECT  1.005000 183.650000 15.455000 183.720000 ;
        RECT  1.005000 183.720000 15.385000 183.790000 ;
        RECT  1.005000 183.790000 15.315000 183.860000 ;
        RECT  1.005000 183.860000 15.245000 183.930000 ;
        RECT  1.005000 183.930000 15.175000 184.000000 ;
        RECT  1.005000 184.000000 15.105000 184.070000 ;
        RECT  1.005000 184.070000 15.035000 184.140000 ;
        RECT  1.005000 184.140000 14.965000 184.210000 ;
        RECT  1.005000 184.210000 14.895000 184.280000 ;
        RECT  1.005000 184.280000 14.825000 184.350000 ;
        RECT  1.005000 184.350000 14.755000 184.420000 ;
        RECT  1.005000 184.420000 14.685000 184.490000 ;
        RECT  1.005000 184.490000 14.615000 184.560000 ;
        RECT  1.005000 184.560000 14.545000 184.630000 ;
        RECT  1.005000 184.630000 14.475000 184.700000 ;
        RECT  1.005000 184.700000 14.405000 184.770000 ;
        RECT  1.005000 184.770000 14.335000 184.840000 ;
        RECT  1.005000 184.840000 14.265000 184.910000 ;
        RECT  1.005000 184.910000 14.195000 184.980000 ;
        RECT  1.005000 184.980000 14.125000 185.050000 ;
        RECT  1.005000 185.050000 14.120000 185.055000 ;
        RECT  1.005000 185.055000 14.120000 189.585000 ;
        RECT  1.005000 189.585000 14.120000 189.655000 ;
        RECT  1.005000 189.655000 14.190000 189.725000 ;
        RECT  1.005000 189.725000 14.260000 189.795000 ;
        RECT  1.005000 189.795000 14.330000 189.865000 ;
        RECT  1.005000 189.865000 14.400000 189.935000 ;
        RECT  1.005000 189.935000 14.470000 190.005000 ;
        RECT  1.005000 190.005000 14.540000 190.075000 ;
        RECT  1.005000 190.075000 14.610000 190.145000 ;
        RECT  1.005000 190.145000 14.680000 190.215000 ;
        RECT  1.005000 190.215000 14.750000 190.285000 ;
        RECT  1.005000 190.285000 14.820000 190.355000 ;
        RECT  1.005000 190.355000 14.890000 190.425000 ;
        RECT  1.005000 190.425000 14.960000 190.495000 ;
        RECT  1.005000 190.495000 15.030000 190.560000 ;
        RECT  1.005000 190.560000 67.200000 195.075000 ;
        RECT  1.010000  47.095000 14.120000  47.100000 ;
        RECT  1.045000  36.855000 16.395000  36.895000 ;
        RECT  1.050000  47.055000 14.120000  47.095000 ;
        RECT  1.085000  36.895000 16.435000  36.935000 ;
        RECT  1.090000  36.935000 16.475000  36.940000 ;
        RECT  1.090000  36.940000 16.480000  37.010000 ;
        RECT  1.090000  37.010000 16.550000  37.080000 ;
        RECT  1.090000  37.080000 16.620000  37.150000 ;
        RECT  1.090000  37.150000 16.690000  37.220000 ;
        RECT  1.090000  37.220000 16.760000  37.290000 ;
        RECT  1.090000  37.290000 16.830000  37.360000 ;
        RECT  1.090000  37.360000 16.900000  37.430000 ;
        RECT  1.090000  37.430000 16.970000  37.500000 ;
        RECT  1.090000  37.500000 17.040000  37.570000 ;
        RECT  1.090000  37.570000 17.110000  37.640000 ;
        RECT  1.090000  37.640000 17.180000  37.710000 ;
        RECT  1.090000  37.710000 17.250000  37.780000 ;
        RECT  1.090000  37.780000 17.320000  37.850000 ;
        RECT  1.090000  37.850000 17.390000  37.920000 ;
        RECT  1.090000  37.920000 17.460000  37.990000 ;
        RECT  1.090000  37.990000 17.530000  38.060000 ;
        RECT  1.090000  38.060000 17.600000  38.130000 ;
        RECT  1.090000  38.130000 17.670000  38.200000 ;
        RECT  1.090000  38.200000 17.740000  38.270000 ;
        RECT  1.090000  38.270000 17.810000  38.340000 ;
        RECT  1.090000  38.340000 17.880000  38.410000 ;
        RECT  1.090000  38.410000 17.950000  38.480000 ;
        RECT  1.090000  38.480000 18.020000  38.550000 ;
        RECT  1.090000  38.550000 18.090000  38.620000 ;
        RECT  1.090000  38.620000 18.160000  38.690000 ;
        RECT  1.090000  38.690000 18.230000  38.760000 ;
        RECT  1.090000  38.760000 18.300000  38.830000 ;
        RECT  1.090000  38.830000 18.370000  38.900000 ;
        RECT  1.090000  38.900000 18.440000  38.970000 ;
        RECT  1.090000  38.970000 18.510000  39.040000 ;
        RECT  1.090000  39.040000 18.580000  39.110000 ;
        RECT  1.090000  39.110000 18.650000  39.180000 ;
        RECT  1.090000  39.180000 18.720000  39.250000 ;
        RECT  1.090000  39.250000 18.790000  39.320000 ;
        RECT  1.090000  39.320000 18.860000  39.390000 ;
        RECT  1.090000  39.390000 18.930000  39.460000 ;
        RECT  1.090000  39.460000 19.000000  39.530000 ;
        RECT  1.090000  39.530000 19.070000  39.600000 ;
        RECT  1.090000  39.600000 19.140000  39.670000 ;
        RECT  1.090000  39.670000 19.210000  39.740000 ;
        RECT  1.090000  39.740000 19.280000  39.810000 ;
        RECT  1.090000  39.810000 19.350000  39.880000 ;
        RECT  1.090000  39.880000 19.420000  39.950000 ;
        RECT  1.090000  39.950000 19.490000  40.020000 ;
        RECT  1.090000  40.020000 19.560000  40.090000 ;
        RECT  1.090000  40.090000 19.630000  40.160000 ;
        RECT  1.090000  40.160000 19.700000  40.230000 ;
        RECT  1.090000  40.230000 19.770000  40.300000 ;
        RECT  1.090000  40.300000 19.840000  40.350000 ;
        RECT  1.090000  40.350000 56.160000  40.420000 ;
        RECT  1.090000  40.420000 56.090000  40.490000 ;
        RECT  1.090000  40.490000 56.020000  40.560000 ;
        RECT  1.090000  40.560000 55.950000  40.630000 ;
        RECT  1.090000  40.630000 55.880000  40.700000 ;
        RECT  1.090000  40.700000 55.810000  40.770000 ;
        RECT  1.090000  40.770000 55.740000  40.840000 ;
        RECT  1.090000  40.840000 55.670000  40.910000 ;
        RECT  1.090000  40.910000 55.600000  40.980000 ;
        RECT  1.090000  40.980000 55.530000  41.050000 ;
        RECT  1.090000  41.050000 55.460000  41.120000 ;
        RECT  1.090000  41.120000 55.390000  41.190000 ;
        RECT  1.090000  41.190000 55.320000  41.260000 ;
        RECT  1.090000  41.260000 55.250000  41.330000 ;
        RECT  1.090000  41.330000 55.180000  41.400000 ;
        RECT  1.090000  41.400000 55.110000  41.470000 ;
        RECT  1.090000  41.470000 55.040000  41.540000 ;
        RECT  1.090000  41.540000 54.970000  41.610000 ;
        RECT  1.090000  41.610000 54.900000  41.680000 ;
        RECT  1.090000  41.680000 54.830000  41.750000 ;
        RECT  1.090000  41.750000 54.760000  41.820000 ;
        RECT  1.090000  41.820000 54.690000  41.890000 ;
        RECT  1.090000  41.890000 54.620000  41.960000 ;
        RECT  1.090000  41.960000 54.550000  42.030000 ;
        RECT  1.090000  42.030000 54.480000  42.100000 ;
        RECT  1.090000  42.100000 54.410000  42.170000 ;
        RECT  1.090000  42.170000 54.340000  42.240000 ;
        RECT  1.090000  42.240000 54.270000  42.310000 ;
        RECT  1.090000  42.310000 54.200000  42.380000 ;
        RECT  1.090000  42.380000 16.985000  42.450000 ;
        RECT  1.090000  42.450000 16.915000  42.520000 ;
        RECT  1.090000  42.520000 16.845000  42.590000 ;
        RECT  1.090000  42.590000 16.775000  42.660000 ;
        RECT  1.090000  42.660000 16.705000  42.730000 ;
        RECT  1.090000  42.730000 16.635000  42.800000 ;
        RECT  1.090000  42.800000 16.565000  42.870000 ;
        RECT  1.090000  42.870000 16.495000  42.940000 ;
        RECT  1.090000  42.940000 16.425000  43.010000 ;
        RECT  1.090000  43.010000 16.355000  43.080000 ;
        RECT  1.090000  43.080000 16.285000  43.150000 ;
        RECT  1.090000  43.150000 16.215000  43.220000 ;
        RECT  1.090000  43.220000 16.145000  43.290000 ;
        RECT  1.090000  43.290000 16.075000  43.360000 ;
        RECT  1.090000  43.360000 16.005000  43.430000 ;
        RECT  1.090000  43.430000 15.935000  43.500000 ;
        RECT  1.090000  43.500000 15.865000  43.570000 ;
        RECT  1.090000  43.570000 15.795000  43.640000 ;
        RECT  1.090000  43.640000 15.725000  43.710000 ;
        RECT  1.090000  43.710000 15.655000  43.780000 ;
        RECT  1.090000  43.780000 15.585000  43.850000 ;
        RECT  1.090000  43.850000 15.515000  43.920000 ;
        RECT  1.090000  43.920000 15.445000  43.990000 ;
        RECT  1.090000  43.990000 15.375000  44.060000 ;
        RECT  1.090000  44.060000 15.305000  44.130000 ;
        RECT  1.090000  44.130000 15.235000  44.200000 ;
        RECT  1.090000  44.200000 15.165000  44.270000 ;
        RECT  1.090000  44.270000 15.095000  44.340000 ;
        RECT  1.090000  44.340000 15.025000  44.410000 ;
        RECT  1.090000  44.410000 14.955000  44.480000 ;
        RECT  1.090000  44.480000 14.885000  44.550000 ;
        RECT  1.090000  44.550000 14.815000  44.620000 ;
        RECT  1.090000  44.620000 14.745000  44.690000 ;
        RECT  1.090000  44.690000 14.675000  44.760000 ;
        RECT  1.090000  44.760000 14.605000  44.830000 ;
        RECT  1.090000  44.830000 14.535000  44.900000 ;
        RECT  1.090000  44.900000 14.465000  44.970000 ;
        RECT  1.090000  44.970000 14.395000  45.040000 ;
        RECT  1.090000  45.040000 14.325000  45.110000 ;
        RECT  1.090000  45.110000 14.255000  45.180000 ;
        RECT  1.090000  45.180000 14.185000  45.250000 ;
        RECT  1.090000  45.250000 14.120000  45.315000 ;
        RECT  1.090000  45.315000 14.120000  47.015000 ;
        RECT  1.090000  47.015000 14.120000  47.055000 ;
        RECT 52.630000  40.295000 56.230000  40.350000 ;
        RECT 52.700000  40.225000 56.285000  40.295000 ;
        RECT 52.770000  40.155000 56.355000  40.225000 ;
        RECT 52.840000  40.085000 56.425000  40.155000 ;
        RECT 52.910000  40.015000 56.495000  40.085000 ;
        RECT 52.980000  39.945000 56.565000  40.015000 ;
        RECT 53.050000  39.875000 56.635000  39.945000 ;
        RECT 53.120000  39.805000 56.705000  39.875000 ;
        RECT 53.190000  39.735000 56.775000  39.805000 ;
        RECT 53.260000  39.665000 56.845000  39.735000 ;
        RECT 53.270000  39.655000 56.915000  39.665000 ;
        RECT 53.340000  39.585000 56.915000  39.655000 ;
        RECT 53.410000  39.515000 56.915000  39.585000 ;
        RECT 53.480000  39.445000 56.915000  39.515000 ;
        RECT 53.550000  39.375000 56.915000  39.445000 ;
        RECT 53.620000  39.305000 56.915000  39.375000 ;
        RECT 53.690000  39.235000 56.915000  39.305000 ;
        RECT 53.760000  39.165000 56.915000  39.235000 ;
        RECT 53.830000  39.095000 56.915000  39.165000 ;
        RECT 53.900000  39.025000 56.915000  39.095000 ;
        RECT 53.970000  38.955000 56.915000  39.025000 ;
        RECT 54.040000  38.885000 56.915000  38.955000 ;
        RECT 54.110000  38.815000 56.915000  38.885000 ;
        RECT 54.180000  38.745000 56.915000  38.815000 ;
        RECT 54.250000  38.675000 56.915000  38.745000 ;
        RECT 54.320000  38.605000 56.915000  38.675000 ;
        RECT 54.390000  38.535000 56.915000  38.605000 ;
        RECT 54.460000  38.465000 56.915000  38.535000 ;
        RECT 54.530000  38.395000 56.915000  38.465000 ;
        RECT 54.600000  38.325000 56.915000  38.395000 ;
        RECT 54.670000  36.115000 56.915000  38.255000 ;
        RECT 54.670000  38.255000 56.915000  38.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT  3.160000 185.360000 25.010000 200.000000 ;
        RECT  3.200000 185.320000 25.010000 185.360000 ;
        RECT  3.350000 185.170000 25.010000 185.320000 ;
        RECT  3.500000 185.020000 25.010000 185.170000 ;
        RECT  3.650000 184.870000 25.010000 185.020000 ;
        RECT  3.800000 184.720000 25.010000 184.870000 ;
        RECT  3.950000 184.570000 25.010000 184.720000 ;
        RECT  4.100000 184.420000 25.010000 184.570000 ;
        RECT  4.250000 184.270000 25.010000 184.420000 ;
        RECT  4.400000 184.120000 25.010000 184.270000 ;
        RECT  4.550000 183.970000 25.010000 184.120000 ;
        RECT  4.700000 183.820000 25.010000 183.970000 ;
        RECT  4.850000 183.670000 25.010000 183.820000 ;
        RECT  5.000000 183.520000 25.010000 183.670000 ;
        RECT  5.150000 183.370000 25.010000 183.520000 ;
        RECT  5.300000 183.220000 25.010000 183.370000 ;
        RECT  5.450000 183.070000 25.010000 183.220000 ;
        RECT  5.600000 182.920000 25.010000 183.070000 ;
        RECT  5.750000 182.770000 25.010000 182.920000 ;
        RECT  5.900000 182.620000 25.010000 182.770000 ;
        RECT  6.050000 182.470000 25.010000 182.620000 ;
        RECT  6.200000 182.320000 25.010000 182.470000 ;
        RECT  6.350000 182.170000 25.010000 182.320000 ;
        RECT  6.500000 182.020000 25.010000 182.170000 ;
        RECT  6.650000 181.870000 25.010000 182.020000 ;
        RECT  6.800000 181.720000 25.010000 181.870000 ;
        RECT  6.950000 181.570000 25.010000 181.720000 ;
        RECT  7.100000 181.420000 25.010000 181.570000 ;
        RECT  7.250000 181.270000 25.010000 181.420000 ;
        RECT  7.400000 181.120000 25.010000 181.270000 ;
        RECT  7.550000 180.970000 25.010000 181.120000 ;
        RECT  7.700000 180.820000 25.010000 180.970000 ;
        RECT  7.850000 180.670000 25.010000 180.820000 ;
        RECT  8.000000 180.520000 25.010000 180.670000 ;
        RECT  8.150000 180.370000 25.010000 180.520000 ;
        RECT  8.300000 180.220000 25.010000 180.370000 ;
        RECT  8.450000 180.070000 25.010000 180.220000 ;
        RECT  8.600000 179.920000 25.010000 180.070000 ;
        RECT  8.750000 179.770000 25.010000 179.920000 ;
        RECT  8.900000 179.620000 25.010000 179.770000 ;
        RECT  9.050000 179.470000 25.010000 179.620000 ;
        RECT  9.200000 179.320000 25.010000 179.470000 ;
        RECT  9.350000 179.170000 25.010000 179.320000 ;
        RECT  9.500000 179.020000 25.010000 179.170000 ;
        RECT  9.650000 178.870000 25.010000 179.020000 ;
        RECT  9.800000 178.720000 25.010000 178.870000 ;
        RECT  9.950000 178.570000 25.010000 178.720000 ;
        RECT 10.100000 178.420000 25.010000 178.570000 ;
        RECT 10.250000 178.270000 25.010000 178.420000 ;
        RECT 10.400000 178.120000 25.010000 178.270000 ;
        RECT 10.550000 177.970000 25.010000 178.120000 ;
        RECT 10.700000 177.820000 25.010000 177.970000 ;
        RECT 10.850000 177.670000 25.010000 177.820000 ;
        RECT 11.000000 177.520000 25.010000 177.670000 ;
        RECT 11.150000 177.370000 25.010000 177.520000 ;
        RECT 11.300000 177.220000 25.010000 177.370000 ;
        RECT 11.450000 177.070000 25.010000 177.220000 ;
        RECT 11.600000 176.920000 25.010000 177.070000 ;
        RECT 11.750000 176.770000 25.010000 176.920000 ;
        RECT 11.900000 176.620000 25.010000 176.770000 ;
        RECT 12.050000 176.470000 25.010000 176.620000 ;
        RECT 12.200000 176.320000 25.010000 176.470000 ;
        RECT 12.350000 176.170000 25.010000 176.320000 ;
        RECT 12.500000 176.020000 25.010000 176.170000 ;
        RECT 12.650000 175.870000 25.010000 176.020000 ;
        RECT 12.800000 175.720000 25.010000 175.870000 ;
        RECT 12.950000 175.570000 25.010000 175.720000 ;
        RECT 13.100000 175.420000 25.010000 175.570000 ;
        RECT 13.250000 175.270000 25.010000 175.420000 ;
        RECT 13.400000 175.120000 25.010000 175.270000 ;
        RECT 13.550000 174.970000 25.010000 175.120000 ;
        RECT 13.700000 174.820000 25.010000 174.970000 ;
        RECT 13.850000 174.670000 25.010000 174.820000 ;
        RECT 14.000000 174.520000 25.010000 174.670000 ;
        RECT 14.150000 174.370000 25.010000 174.520000 ;
        RECT 14.300000 174.220000 25.010000 174.370000 ;
        RECT 14.450000 174.070000 25.010000 174.220000 ;
        RECT 14.600000 173.920000 25.010000 174.070000 ;
        RECT 14.750000 173.770000 25.010000 173.920000 ;
        RECT 14.900000 173.620000 25.010000 173.770000 ;
        RECT 15.050000 173.470000 25.010000 173.620000 ;
        RECT 15.200000 173.320000 25.010000 173.470000 ;
        RECT 15.350000 173.170000 25.010000 173.320000 ;
        RECT 15.500000 102.200000 23.830000 102.350000 ;
        RECT 15.500000 102.350000 23.680000 102.500000 ;
        RECT 15.500000 102.500000 23.530000 102.650000 ;
        RECT 15.500000 102.650000 23.380000 102.800000 ;
        RECT 15.500000 102.800000 23.230000 102.950000 ;
        RECT 15.500000 102.950000 23.080000 103.100000 ;
        RECT 15.500000 103.100000 22.930000 103.250000 ;
        RECT 15.500000 103.250000 22.780000 103.400000 ;
        RECT 15.500000 103.400000 22.630000 103.550000 ;
        RECT 15.500000 103.550000 22.480000 103.700000 ;
        RECT 15.500000 103.700000 22.330000 103.850000 ;
        RECT 15.500000 103.850000 22.180000 104.000000 ;
        RECT 15.500000 104.000000 22.030000 104.150000 ;
        RECT 15.500000 104.150000 21.880000 104.300000 ;
        RECT 15.500000 104.300000 21.730000 104.450000 ;
        RECT 15.500000 104.450000 21.580000 104.600000 ;
        RECT 15.500000 104.600000 21.500000 104.680000 ;
        RECT 15.500000 104.680000 21.500000 169.130000 ;
        RECT 15.500000 169.130000 21.500000 169.280000 ;
        RECT 15.500000 169.280000 21.650000 169.430000 ;
        RECT 15.500000 169.430000 21.800000 169.580000 ;
        RECT 15.500000 169.580000 21.950000 169.730000 ;
        RECT 15.500000 169.730000 22.100000 169.880000 ;
        RECT 15.500000 169.880000 22.250000 170.030000 ;
        RECT 15.500000 170.030000 22.400000 170.180000 ;
        RECT 15.500000 170.180000 22.550000 170.330000 ;
        RECT 15.500000 170.330000 22.700000 170.480000 ;
        RECT 15.500000 170.480000 22.850000 170.630000 ;
        RECT 15.500000 170.630000 23.000000 170.780000 ;
        RECT 15.500000 170.780000 23.150000 170.930000 ;
        RECT 15.500000 170.930000 23.300000 171.080000 ;
        RECT 15.500000 171.080000 23.450000 171.230000 ;
        RECT 15.500000 171.230000 23.600000 171.380000 ;
        RECT 15.500000 171.380000 23.750000 171.530000 ;
        RECT 15.500000 171.530000 23.900000 171.680000 ;
        RECT 15.500000 171.680000 24.050000 171.830000 ;
        RECT 15.500000 171.830000 24.200000 171.980000 ;
        RECT 15.500000 171.980000 24.350000 172.130000 ;
        RECT 15.500000 172.130000 24.500000 172.280000 ;
        RECT 15.500000 172.280000 24.650000 172.430000 ;
        RECT 15.500000 172.430000 24.800000 172.580000 ;
        RECT 15.500000 172.580000 24.950000 172.640000 ;
        RECT 15.500000 172.640000 25.010000 173.020000 ;
        RECT 15.500000 173.020000 25.010000 173.170000 ;
        RECT 15.645000 102.055000 23.980000 102.200000 ;
        RECT 15.795000 101.905000 24.125000 102.055000 ;
        RECT 15.945000 101.755000 24.275000 101.905000 ;
        RECT 16.095000 101.605000 24.425000 101.755000 ;
        RECT 16.245000 101.455000 24.575000 101.605000 ;
        RECT 16.395000 101.305000 24.725000 101.455000 ;
        RECT 16.545000 101.155000 24.875000 101.305000 ;
        RECT 16.695000 101.005000 25.025000 101.155000 ;
        RECT 16.845000 100.855000 25.175000 101.005000 ;
        RECT 16.995000 100.705000 25.325000 100.855000 ;
        RECT 17.145000 100.555000 25.475000 100.705000 ;
        RECT 17.295000 100.405000 25.625000 100.555000 ;
        RECT 17.445000 100.255000 25.775000 100.405000 ;
        RECT 17.595000 100.105000 25.925000 100.255000 ;
        RECT 17.745000  99.955000 26.075000 100.105000 ;
        RECT 17.895000  99.805000 26.225000  99.955000 ;
        RECT 18.045000  99.655000 26.375000  99.805000 ;
        RECT 18.195000  99.505000 26.525000  99.655000 ;
        RECT 18.345000  99.355000 26.675000  99.505000 ;
        RECT 18.495000  99.205000 26.825000  99.355000 ;
        RECT 18.645000  99.055000 26.975000  99.205000 ;
        RECT 18.795000  98.905000 27.125000  99.055000 ;
        RECT 18.945000  98.755000 27.275000  98.905000 ;
        RECT 19.095000  98.605000 27.425000  98.755000 ;
        RECT 19.245000  98.455000 27.575000  98.605000 ;
        RECT 19.395000  98.305000 27.725000  98.455000 ;
        RECT 19.545000  98.155000 27.875000  98.305000 ;
        RECT 19.695000  98.005000 28.025000  98.155000 ;
        RECT 19.845000  97.855000 28.175000  98.005000 ;
        RECT 19.995000  97.705000 28.325000  97.855000 ;
        RECT 20.145000  97.555000 28.475000  97.705000 ;
        RECT 20.295000  97.405000 28.625000  97.555000 ;
        RECT 20.445000  97.255000 28.775000  97.405000 ;
        RECT 20.595000  97.105000 28.925000  97.255000 ;
        RECT 20.745000  96.955000 29.075000  97.105000 ;
        RECT 20.895000  96.805000 29.225000  96.955000 ;
        RECT 21.045000  96.655000 29.375000  96.805000 ;
        RECT 21.195000  96.505000 29.525000  96.655000 ;
        RECT 21.345000  96.355000 29.525000  96.505000 ;
        RECT 21.495000  96.205000 29.525000  96.355000 ;
        RECT 21.645000  96.055000 29.525000  96.205000 ;
        RECT 21.795000  95.905000 29.525000  96.055000 ;
        RECT 21.945000  95.755000 29.525000  95.905000 ;
        RECT 22.095000  95.605000 29.525000  95.755000 ;
        RECT 22.245000  95.455000 29.525000  95.605000 ;
        RECT 22.395000  95.305000 29.525000  95.455000 ;
        RECT 22.545000  95.155000 29.525000  95.305000 ;
        RECT 22.695000  95.005000 29.525000  95.155000 ;
        RECT 22.845000  94.855000 29.525000  95.005000 ;
        RECT 22.995000  94.705000 29.525000  94.855000 ;
        RECT 23.145000  94.555000 29.525000  94.705000 ;
        RECT 23.295000  94.405000 29.525000  94.555000 ;
        RECT 23.445000  94.255000 29.525000  94.405000 ;
        RECT 23.595000  94.105000 29.525000  94.255000 ;
        RECT 23.745000  92.540000 29.935000  92.690000 ;
        RECT 23.745000  92.690000 29.785000  92.840000 ;
        RECT 23.745000  92.840000 29.635000  92.990000 ;
        RECT 23.745000  92.990000 29.525000  93.100000 ;
        RECT 23.745000  93.100000 29.525000  93.955000 ;
        RECT 23.745000  93.955000 29.525000  94.105000 ;
        RECT 23.820000  92.465000 30.085000  92.540000 ;
        RECT 23.895000  92.390000 30.160000  92.465000 ;
        RECT 23.945000  92.340000 36.895000  92.390000 ;
        RECT 24.095000  92.190000 36.895000  92.340000 ;
        RECT 24.245000  92.040000 36.895000  92.190000 ;
        RECT 24.395000  91.890000 36.895000  92.040000 ;
        RECT 24.545000  91.740000 36.895000  91.890000 ;
        RECT 24.695000  91.590000 36.895000  91.740000 ;
        RECT 24.845000  91.440000 36.895000  91.590000 ;
        RECT 24.995000  91.290000 36.895000  91.440000 ;
        RECT 25.145000  91.140000 36.895000  91.290000 ;
        RECT 25.295000  90.990000 36.895000  91.140000 ;
        RECT 25.445000  90.840000 36.895000  90.990000 ;
        RECT 25.595000  90.690000 36.895000  90.840000 ;
        RECT 25.745000  90.540000 36.895000  90.690000 ;
        RECT 25.895000   0.000000 36.895000  90.390000 ;
        RECT 25.895000  90.390000 36.895000  90.540000 ;
        RECT 25.930000 102.390000 34.250000 102.540000 ;
        RECT 25.930000 102.540000 34.100000 102.690000 ;
        RECT 25.930000 102.690000 33.950000 102.840000 ;
        RECT 25.930000 102.840000 33.800000 102.990000 ;
        RECT 25.930000 102.990000 33.650000 103.140000 ;
        RECT 25.930000 103.140000 33.500000 103.290000 ;
        RECT 25.930000 103.290000 33.350000 103.440000 ;
        RECT 25.930000 103.440000 33.200000 103.590000 ;
        RECT 25.930000 103.590000 33.050000 103.740000 ;
        RECT 25.930000 103.740000 32.900000 103.890000 ;
        RECT 25.930000 103.890000 32.750000 104.040000 ;
        RECT 25.930000 104.040000 32.600000 104.190000 ;
        RECT 25.930000 104.190000 32.450000 104.340000 ;
        RECT 25.930000 104.340000 32.300000 104.490000 ;
        RECT 25.930000 104.490000 32.150000 104.640000 ;
        RECT 25.930000 104.640000 32.000000 104.790000 ;
        RECT 25.930000 104.790000 31.930000 104.860000 ;
        RECT 25.930000 104.860000 31.930000 170.460000 ;
        RECT 25.930000 170.460000 31.930000 170.610000 ;
        RECT 25.930000 170.610000 32.080000 170.760000 ;
        RECT 25.930000 170.760000 32.230000 170.910000 ;
        RECT 25.930000 170.910000 32.380000 171.060000 ;
        RECT 25.930000 171.060000 32.530000 171.210000 ;
        RECT 25.930000 171.210000 32.680000 171.360000 ;
        RECT 25.930000 171.360000 32.830000 171.510000 ;
        RECT 25.930000 171.510000 32.980000 171.660000 ;
        RECT 25.930000 171.660000 33.130000 171.810000 ;
        RECT 25.930000 171.810000 33.280000 171.960000 ;
        RECT 25.930000 171.960000 33.430000 172.110000 ;
        RECT 25.930000 172.110000 33.580000 172.260000 ;
        RECT 25.930000 172.260000 33.730000 172.410000 ;
        RECT 25.930000 172.410000 33.880000 172.560000 ;
        RECT 25.930000 172.560000 34.030000 172.710000 ;
        RECT 25.930000 172.710000 34.180000 172.860000 ;
        RECT 25.930000 172.860000 34.330000 173.010000 ;
        RECT 25.930000 173.010000 34.480000 173.160000 ;
        RECT 25.930000 173.160000 34.630000 173.310000 ;
        RECT 25.930000 173.310000 34.780000 173.460000 ;
        RECT 25.930000 173.460000 34.930000 173.610000 ;
        RECT 25.930000 173.610000 35.080000 173.760000 ;
        RECT 25.930000 173.760000 35.230000 173.910000 ;
        RECT 25.930000 173.910000 35.380000 174.060000 ;
        RECT 25.930000 174.060000 35.530000 174.210000 ;
        RECT 25.930000 174.210000 35.680000 174.360000 ;
        RECT 25.930000 174.360000 35.830000 174.510000 ;
        RECT 25.930000 174.510000 35.980000 174.660000 ;
        RECT 25.930000 174.660000 36.130000 174.810000 ;
        RECT 25.930000 174.810000 36.280000 174.960000 ;
        RECT 25.930000 174.960000 36.430000 175.110000 ;
        RECT 25.930000 175.110000 36.580000 175.260000 ;
        RECT 25.930000 175.260000 36.730000 175.350000 ;
        RECT 25.930000 175.350000 36.820000 200.000000 ;
        RECT 26.025000 102.295000 34.400000 102.390000 ;
        RECT 26.175000 102.145000 34.495000 102.295000 ;
        RECT 26.325000 101.995000 34.645000 102.145000 ;
        RECT 26.475000 101.845000 34.795000 101.995000 ;
        RECT 26.625000 101.695000 34.945000 101.845000 ;
        RECT 26.775000 101.545000 35.095000 101.695000 ;
        RECT 26.925000 101.395000 35.245000 101.545000 ;
        RECT 27.075000 101.245000 35.395000 101.395000 ;
        RECT 27.225000 101.095000 35.545000 101.245000 ;
        RECT 27.375000 100.945000 35.695000 101.095000 ;
        RECT 27.525000 100.795000 35.845000 100.945000 ;
        RECT 27.675000 100.645000 35.995000 100.795000 ;
        RECT 27.825000 100.495000 36.145000 100.645000 ;
        RECT 27.975000 100.345000 36.295000 100.495000 ;
        RECT 28.125000 100.195000 36.445000 100.345000 ;
        RECT 28.275000 100.045000 36.595000 100.195000 ;
        RECT 28.425000  99.895000 36.745000 100.045000 ;
        RECT 28.495000  99.825000 36.895000  99.895000 ;
        RECT 28.645000  99.675000 36.895000  99.825000 ;
        RECT 28.795000  99.525000 36.895000  99.675000 ;
        RECT 28.945000  99.375000 36.895000  99.525000 ;
        RECT 29.095000  99.225000 36.895000  99.375000 ;
        RECT 29.245000  99.075000 36.895000  99.225000 ;
        RECT 29.395000  98.925000 36.895000  99.075000 ;
        RECT 29.545000  98.775000 36.895000  98.925000 ;
        RECT 29.695000  98.625000 36.895000  98.775000 ;
        RECT 29.845000  98.475000 36.895000  98.625000 ;
        RECT 29.995000  98.325000 36.895000  98.475000 ;
        RECT 30.145000  98.175000 36.895000  98.325000 ;
        RECT 30.295000  98.025000 36.895000  98.175000 ;
        RECT 30.445000  97.875000 36.895000  98.025000 ;
        RECT 30.595000  97.725000 36.895000  97.875000 ;
        RECT 30.745000  97.575000 36.895000  97.725000 ;
        RECT 30.895000  97.425000 36.895000  97.575000 ;
        RECT 31.045000  97.275000 36.895000  97.425000 ;
        RECT 31.195000  97.125000 36.895000  97.275000 ;
        RECT 31.345000  96.975000 36.895000  97.125000 ;
        RECT 31.385000  92.390000 36.895000  92.540000 ;
        RECT 31.495000  96.825000 36.895000  96.975000 ;
        RECT 31.535000  92.540000 36.895000  92.690000 ;
        RECT 31.645000  96.675000 36.895000  96.825000 ;
        RECT 31.685000  92.690000 36.895000  92.840000 ;
        RECT 31.795000  96.525000 36.895000  96.675000 ;
        RECT 31.835000  92.840000 36.895000  92.990000 ;
        RECT 31.945000  92.990000 36.895000  93.100000 ;
        RECT 31.945000  93.100000 36.895000  96.375000 ;
        RECT 31.945000  96.375000 36.895000  96.525000 ;
    END
  END SRC_BDY_HVC
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.835000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  1.070000  43.270000  1.400000  43.440000 ;
      RECT  1.145000  43.440000  1.315000  43.810000 ;
      RECT  3.100000  27.160000 48.200000  28.030000 ;
      RECT  3.100000  28.030000  4.020000  38.695000 ;
      RECT  3.100000  38.695000 48.200000  39.565000 ;
      RECT  3.130000  27.140000 48.200000  27.160000 ;
      RECT  3.130000  39.565000 48.200000  39.585000 ;
      RECT  4.735000  29.230000 45.955000  29.430000 ;
      RECT  4.735000  29.430000  4.905000  37.425000 ;
      RECT  4.735000  37.425000 45.955000  37.595000 ;
      RECT  6.115000  29.780000  6.285000  36.570000 ;
      RECT  6.340000  36.970000 45.060000  37.230000 ;
      RECT  6.895000  29.775000  7.065000  36.570000 ;
      RECT  7.675000  29.780000  7.845000  36.570000 ;
      RECT  8.050000  43.270000  8.690000  43.440000 ;
      RECT  8.455000  29.770000  8.625000  36.570000 ;
      RECT  8.510000 162.655000 10.360000 169.150000 ;
      RECT  9.135000  43.505000 70.125000  44.755000 ;
      RECT  9.135000  44.755000 10.385000  71.570000 ;
      RECT  9.135000  71.570000 21.085000  72.820000 ;
      RECT  9.150000 169.400000 10.400000 198.445000 ;
      RECT  9.150000 198.445000 70.125000 199.695000 ;
      RECT  9.170000 133.350000 20.990000 134.540000 ;
      RECT  9.170000 134.540000 10.360000 162.655000 ;
      RECT  9.170000 169.150000 10.360000 169.400000 ;
      RECT  9.200000 133.205000 14.190000 133.350000 ;
      RECT  9.235000  29.780000  9.405000  36.570000 ;
      RECT  9.405000  74.180000  9.935000  74.350000 ;
      RECT  9.500000  74.350000  9.830000  74.355000 ;
      RECT 10.015000  29.775000 10.185000  36.570000 ;
      RECT 10.770000 162.655000 11.975000 169.905000 ;
      RECT 10.795000  29.780000 10.965000  36.570000 ;
      RECT 11.100000 170.415000 11.990000 196.835000 ;
      RECT 11.100000 196.835000 68.155000 197.725000 ;
      RECT 11.105000  45.460000 68.155000  46.350000 ;
      RECT 11.105000  46.350000 11.995000  69.975000 ;
      RECT 11.105000  69.975000 22.680000  70.865000 ;
      RECT 11.125000 135.315000 22.660000 136.165000 ;
      RECT 11.125000 136.165000 12.100000 158.915000 ;
      RECT 11.125000 158.915000 11.975000 162.655000 ;
      RECT 11.125000 169.905000 11.975000 170.415000 ;
      RECT 11.575000  29.770000 11.745000  36.570000 ;
      RECT 12.065000   1.000000 70.650000   1.890000 ;
      RECT 12.065000   1.890000 13.045000  22.230000 ;
      RECT 12.065000  22.230000 56.085000  22.350000 ;
      RECT 12.065000  22.350000 56.105000  23.240000 ;
      RECT 12.355000  29.780000 12.525000  36.570000 ;
      RECT 12.400000 159.555000 64.500000 161.990000 ;
      RECT 12.830000 182.570000 66.685000 184.990000 ;
      RECT 13.085000  46.815000 64.500000  46.990000 ;
      RECT 13.085000  46.990000 13.255000  67.965000 ;
      RECT 13.090000  46.740000 64.500000  46.815000 ;
      RECT 13.135000  29.775000 13.305000  36.570000 ;
      RECT 13.780000   4.820000 14.010000   8.825000 ;
      RECT 13.780000   8.825000 68.570000   9.055000 ;
      RECT 13.780000  11.040000 14.010000  15.045000 ;
      RECT 13.780000  15.045000 68.570000  15.275000 ;
      RECT 13.780000  17.260000 14.010000  21.265000 ;
      RECT 13.780000  21.265000 68.570000  21.495000 ;
      RECT 13.810000   2.635000 68.540000   2.835000 ;
      RECT 13.810000   2.835000 13.980000   4.820000 ;
      RECT 13.810000   9.055000 13.980000  11.040000 ;
      RECT 13.810000  15.275000 13.980000  17.260000 ;
      RECT 13.915000  29.780000 14.085000  36.570000 ;
      RECT 13.980000   2.605000 19.570000   2.635000 ;
      RECT 14.385000  47.160000 15.435000  66.930000 ;
      RECT 14.385000 139.160000 15.435000 158.930000 ;
      RECT 14.385000 162.160000 15.435000 181.930000 ;
      RECT 14.385000 185.160000 15.435000 195.185000 ;
      RECT 14.515000   4.820000 14.745000   7.770000 ;
      RECT 14.515000  11.040000 14.745000  13.990000 ;
      RECT 14.515000  17.260000 14.745000  20.210000 ;
      RECT 14.550000   3.755000 14.720000   4.820000 ;
      RECT 14.550000   7.770000 14.720000   8.505000 ;
      RECT 14.550000   9.975000 14.720000  11.040000 ;
      RECT 14.550000  13.990000 14.720000  14.725000 ;
      RECT 14.550000  16.195000 14.720000  17.260000 ;
      RECT 14.550000  20.210000 14.720000  20.945000 ;
      RECT 14.695000  29.770000 14.865000  36.570000 ;
      RECT 14.775000   3.075000 18.775000   3.305000 ;
      RECT 14.775000   9.295000 18.775000   9.525000 ;
      RECT 14.775000  15.515000 18.775000  15.745000 ;
      RECT 15.475000  29.780000 15.645000  36.570000 ;
      RECT 15.705000  67.340000 64.500000  68.995000 ;
      RECT 15.780000 136.540000 64.500000 138.990000 ;
      RECT 15.780000 159.340000 64.500000 159.555000 ;
      RECT 15.780000 182.340000 66.685000 182.570000 ;
      RECT 15.780000 195.370000 16.490000 195.540000 ;
      RECT 16.255000  29.770000 16.425000  36.570000 ;
      RECT 16.865000  47.525000 17.395000  65.695000 ;
      RECT 16.865000 139.525000 17.395000 157.695000 ;
      RECT 16.865000 162.525000 17.395000 180.695000 ;
      RECT 16.865000 185.525000 17.395000 195.055000 ;
      RECT 16.885000  47.325000 17.395000  47.525000 ;
      RECT 16.885000  65.695000 17.395000  67.035000 ;
      RECT 16.885000 139.325000 17.395000 139.525000 ;
      RECT 16.885000 157.695000 17.395000 159.035000 ;
      RECT 16.885000 162.325000 17.395000 162.525000 ;
      RECT 16.885000 180.695000 17.395000 182.035000 ;
      RECT 16.885000 185.325000 17.395000 185.525000 ;
      RECT 17.035000  29.780000 17.205000  36.570000 ;
      RECT 17.790000 195.370000 18.500000 195.540000 ;
      RECT 17.815000  29.770000 17.985000  36.570000 ;
      RECT 17.835000 133.145000 20.990000 133.350000 ;
      RECT 18.410000  74.185000 18.740000  74.200000 ;
      RECT 18.410000  74.200000 19.000000  74.370000 ;
      RECT 18.410000  74.370000 18.740000  74.385000 ;
      RECT 18.595000  29.780000 18.765000  36.570000 ;
      RECT 18.810000   4.820000 19.040000   7.770000 ;
      RECT 18.810000  11.040000 19.040000  13.990000 ;
      RECT 18.810000  17.260000 19.040000  20.210000 ;
      RECT 18.830000   3.755000 19.000000   4.820000 ;
      RECT 18.830000   7.770000 19.000000   8.505000 ;
      RECT 18.830000   9.975000 19.000000  11.040000 ;
      RECT 18.830000  13.990000 19.000000  14.725000 ;
      RECT 18.830000  16.195000 19.000000  17.260000 ;
      RECT 18.830000  20.210000 19.000000  20.945000 ;
      RECT 18.845000  47.160000 20.035000  66.870000 ;
      RECT 18.845000 139.160000 20.035000 158.870000 ;
      RECT 18.845000 162.160000 20.035000 181.870000 ;
      RECT 18.845000 185.160000 20.035000 195.010000 ;
      RECT 18.985000 195.010000 19.875000 195.075000 ;
      RECT 19.375000  29.775000 19.545000  36.570000 ;
      RECT 19.540000   4.820000 19.770000   8.825000 ;
      RECT 19.540000  11.040000 19.770000  15.045000 ;
      RECT 19.540000  17.260000 19.770000  21.265000 ;
      RECT 19.565000  97.500000 20.990000 133.145000 ;
      RECT 19.570000   2.835000 19.740000   4.820000 ;
      RECT 19.570000   9.055000 19.740000  11.040000 ;
      RECT 19.570000  15.275000 19.740000  17.260000 ;
      RECT 19.740000   2.605000 29.330000   2.635000 ;
      RECT 19.800000  72.820000 21.085000  96.895000 ;
      RECT 19.800000  96.895000 20.990000  97.500000 ;
      RECT 20.155000  29.780000 20.325000  36.570000 ;
      RECT 20.275000   4.820000 20.505000   7.770000 ;
      RECT 20.275000  11.040000 20.505000  13.990000 ;
      RECT 20.275000  17.260000 20.505000  20.210000 ;
      RECT 20.310000   3.755000 20.480000   4.820000 ;
      RECT 20.310000   7.770000 20.480000   8.505000 ;
      RECT 20.310000   9.975000 20.480000  11.040000 ;
      RECT 20.310000  13.990000 20.480000  14.725000 ;
      RECT 20.310000  16.195000 20.480000  17.260000 ;
      RECT 20.310000  20.210000 20.480000  20.945000 ;
      RECT 20.380000 195.370000 21.090000 195.540000 ;
      RECT 20.535000   3.075000 28.535000   3.305000 ;
      RECT 20.535000   9.295000 28.535000   9.525000 ;
      RECT 20.535000  15.515000 28.535000  15.745000 ;
      RECT 20.935000  29.770000 21.105000  36.570000 ;
      RECT 21.465000  47.525000 21.995000  65.695000 ;
      RECT 21.465000 139.525000 21.995000 157.695000 ;
      RECT 21.465000 162.525000 21.995000 180.695000 ;
      RECT 21.465000 185.525000 21.995000 195.055000 ;
      RECT 21.485000  47.325000 21.995000  47.525000 ;
      RECT 21.485000  65.695000 21.995000  67.035000 ;
      RECT 21.485000 139.325000 21.995000 139.525000 ;
      RECT 21.485000 157.695000 21.995000 159.035000 ;
      RECT 21.485000 162.325000 21.995000 162.525000 ;
      RECT 21.485000 180.695000 21.995000 182.035000 ;
      RECT 21.485000 185.325000 21.995000 185.525000 ;
      RECT 21.715000  29.780000 21.885000  36.570000 ;
      RECT 21.790000  70.865000 22.680000  97.450000 ;
      RECT 21.810000  97.450000 22.660000 135.315000 ;
      RECT 22.390000 195.370000 23.100000 195.540000 ;
      RECT 22.495000  29.775000 22.665000  36.570000 ;
      RECT 23.025000  90.495000 64.500000  92.990000 ;
      RECT 23.055000 113.340000 64.500000 115.990000 ;
      RECT 23.275000  29.780000 23.445000  36.570000 ;
      RECT 23.445000  47.160000 24.635000  66.870000 ;
      RECT 23.445000 139.160000 24.635000 158.870000 ;
      RECT 23.445000 162.160000 24.635000 181.870000 ;
      RECT 23.445000 185.160000 24.635000 195.010000 ;
      RECT 23.510000  68.995000 64.500000  69.990000 ;
      RECT 23.585000  70.160000 24.635000  89.930000 ;
      RECT 23.585000  93.160000 24.635000 112.930000 ;
      RECT 23.585000 116.160000 24.635000 135.930000 ;
      RECT 23.585000 195.010000 24.475000 195.030000 ;
      RECT 24.055000  29.770000 24.225000  36.570000 ;
      RECT 24.835000  29.780000 25.005000  36.570000 ;
      RECT 24.980000  90.370000 64.500000  90.495000 ;
      RECT 24.980000 136.370000 64.500000 136.540000 ;
      RECT 24.980000 195.370000 25.690000 195.540000 ;
      RECT 25.615000  29.775000 25.785000  36.570000 ;
      RECT 25.670000  90.340000 64.500000  90.370000 ;
      RECT 25.670000 136.340000 64.500000 136.370000 ;
      RECT 26.065000  47.525000 26.595000  65.695000 ;
      RECT 26.065000  70.525000 26.595000  88.695000 ;
      RECT 26.065000  93.525000 26.595000 111.695000 ;
      RECT 26.065000 116.525000 26.595000 134.695000 ;
      RECT 26.065000 139.525000 26.595000 157.695000 ;
      RECT 26.065000 162.525000 26.595000 180.695000 ;
      RECT 26.065000 185.525000 26.595000 195.055000 ;
      RECT 26.085000  47.325000 26.595000  47.525000 ;
      RECT 26.085000  65.695000 26.595000  67.035000 ;
      RECT 26.085000  70.325000 26.595000  70.525000 ;
      RECT 26.085000  88.695000 26.595000  90.035000 ;
      RECT 26.085000  93.325000 26.595000  93.525000 ;
      RECT 26.085000 111.695000 26.595000 113.035000 ;
      RECT 26.085000 116.325000 26.595000 116.525000 ;
      RECT 26.085000 134.695000 26.595000 136.035000 ;
      RECT 26.085000 139.325000 26.595000 139.525000 ;
      RECT 26.085000 157.695000 26.595000 159.035000 ;
      RECT 26.085000 162.325000 26.595000 162.525000 ;
      RECT 26.085000 180.695000 26.595000 182.035000 ;
      RECT 26.085000 185.325000 26.595000 185.525000 ;
      RECT 26.395000  29.780000 26.565000  36.570000 ;
      RECT 26.990000 195.370000 27.700000 195.540000 ;
      RECT 27.175000  29.770000 27.345000  36.570000 ;
      RECT 27.955000  29.780000 28.125000  36.570000 ;
      RECT 28.045000  47.160000 29.235000  66.870000 ;
      RECT 28.045000  70.160000 29.235000  89.870000 ;
      RECT 28.045000  93.160000 29.235000 112.870000 ;
      RECT 28.045000 116.160000 29.235000 135.870000 ;
      RECT 28.045000 139.160000 29.235000 158.870000 ;
      RECT 28.045000 162.160000 29.235000 181.870000 ;
      RECT 28.045000 185.160000 29.235000 195.010000 ;
      RECT 28.185000 195.010000 29.075000 195.030000 ;
      RECT 28.570000   4.820000 28.800000   7.770000 ;
      RECT 28.570000  11.040000 28.800000  13.990000 ;
      RECT 28.570000  17.260000 28.800000  20.210000 ;
      RECT 28.590000   3.755000 28.760000   4.820000 ;
      RECT 28.590000   7.770000 28.760000   8.505000 ;
      RECT 28.590000   9.975000 28.760000  11.040000 ;
      RECT 28.590000  13.990000 28.760000  14.725000 ;
      RECT 28.590000  16.195000 28.760000  17.260000 ;
      RECT 28.590000  20.210000 28.760000  20.945000 ;
      RECT 28.735000  29.775000 28.905000  36.570000 ;
      RECT 29.300000   4.820000 29.530000   8.825000 ;
      RECT 29.300000  11.040000 29.530000  15.045000 ;
      RECT 29.300000  17.260000 29.530000  21.265000 ;
      RECT 29.330000   2.835000 29.500000   4.820000 ;
      RECT 29.330000   9.055000 29.500000  11.040000 ;
      RECT 29.330000  15.275000 29.500000  17.260000 ;
      RECT 29.500000   2.605000 39.090000   2.635000 ;
      RECT 29.515000  29.780000 29.685000  36.570000 ;
      RECT 29.580000 195.370000 30.290000 195.540000 ;
      RECT 30.035000   4.820000 30.265000   7.770000 ;
      RECT 30.035000  11.040000 30.265000  13.990000 ;
      RECT 30.035000  17.260000 30.265000  20.210000 ;
      RECT 30.070000   3.755000 30.240000   4.820000 ;
      RECT 30.070000   7.770000 30.240000   8.505000 ;
      RECT 30.070000   9.975000 30.240000  11.040000 ;
      RECT 30.070000  13.990000 30.240000  14.725000 ;
      RECT 30.070000  16.195000 30.240000  17.260000 ;
      RECT 30.070000  20.210000 30.240000  20.945000 ;
      RECT 30.295000   3.075000 38.295000   3.305000 ;
      RECT 30.295000   9.295000 38.295000   9.525000 ;
      RECT 30.295000  15.515000 38.295000  15.745000 ;
      RECT 30.295000  29.770000 30.465000  36.570000 ;
      RECT 30.665000  47.525000 31.195000  65.695000 ;
      RECT 30.665000  70.525000 31.195000  88.695000 ;
      RECT 30.665000  93.525000 31.195000 111.695000 ;
      RECT 30.665000 116.525000 31.195000 134.695000 ;
      RECT 30.665000 139.525000 31.195000 157.695000 ;
      RECT 30.665000 162.525000 31.195000 180.695000 ;
      RECT 30.665000 185.525000 31.195000 195.055000 ;
      RECT 30.685000  47.325000 31.195000  47.525000 ;
      RECT 30.685000  65.695000 31.195000  67.035000 ;
      RECT 30.685000  70.325000 31.195000  70.525000 ;
      RECT 30.685000  88.695000 31.195000  90.035000 ;
      RECT 30.685000  93.325000 31.195000  93.525000 ;
      RECT 30.685000 111.695000 31.195000 113.035000 ;
      RECT 30.685000 116.325000 31.195000 116.525000 ;
      RECT 30.685000 134.695000 31.195000 136.035000 ;
      RECT 30.685000 139.325000 31.195000 139.525000 ;
      RECT 30.685000 157.695000 31.195000 159.035000 ;
      RECT 30.685000 162.325000 31.195000 162.525000 ;
      RECT 30.685000 180.695000 31.195000 182.035000 ;
      RECT 30.685000 185.325000 31.195000 185.525000 ;
      RECT 31.075000  29.780000 31.245000  36.570000 ;
      RECT 31.590000 195.370000 32.300000 195.540000 ;
      RECT 31.855000  29.775000 32.025000  36.570000 ;
      RECT 32.635000  29.780000 32.805000  36.570000 ;
      RECT 32.645000  47.160000 33.835000  66.870000 ;
      RECT 32.645000  70.160000 33.835000  89.870000 ;
      RECT 32.645000  93.160000 33.835000 112.870000 ;
      RECT 32.645000 116.160000 33.835000 135.870000 ;
      RECT 32.645000 139.160000 33.835000 158.870000 ;
      RECT 32.645000 162.160000 33.835000 181.870000 ;
      RECT 32.645000 185.160000 33.835000 195.010000 ;
      RECT 32.785000 195.010000 33.675000 195.030000 ;
      RECT 33.415000  29.770000 33.585000  36.570000 ;
      RECT 34.180000 195.370000 34.890000 195.540000 ;
      RECT 34.195000  29.780000 34.365000  36.570000 ;
      RECT 34.975000  29.775000 35.145000  36.570000 ;
      RECT 35.265000  47.525000 35.795000  65.695000 ;
      RECT 35.265000  70.525000 35.795000  88.695000 ;
      RECT 35.265000  93.525000 35.795000 111.695000 ;
      RECT 35.265000 116.525000 35.795000 134.695000 ;
      RECT 35.265000 139.525000 35.795000 157.695000 ;
      RECT 35.265000 162.525000 35.795000 180.695000 ;
      RECT 35.265000 185.525000 35.795000 195.055000 ;
      RECT 35.285000  47.325000 35.795000  47.525000 ;
      RECT 35.285000  65.695000 35.795000  67.035000 ;
      RECT 35.285000  70.325000 35.795000  70.525000 ;
      RECT 35.285000  88.695000 35.795000  90.035000 ;
      RECT 35.285000  93.325000 35.795000  93.525000 ;
      RECT 35.285000 111.695000 35.795000 113.035000 ;
      RECT 35.285000 116.325000 35.795000 116.525000 ;
      RECT 35.285000 134.695000 35.795000 136.035000 ;
      RECT 35.285000 139.325000 35.795000 139.525000 ;
      RECT 35.285000 157.695000 35.795000 159.035000 ;
      RECT 35.285000 162.325000 35.795000 162.525000 ;
      RECT 35.285000 180.695000 35.795000 182.035000 ;
      RECT 35.285000 185.325000 35.795000 185.525000 ;
      RECT 35.755000  29.780000 35.925000  36.570000 ;
      RECT 36.190000 195.370000 36.900000 195.540000 ;
      RECT 36.535000  29.770000 36.705000  36.570000 ;
      RECT 37.245000  47.160000 38.435000  66.870000 ;
      RECT 37.245000  70.160000 38.435000  89.870000 ;
      RECT 37.245000  93.160000 38.435000 112.870000 ;
      RECT 37.245000 116.160000 38.435000 135.870000 ;
      RECT 37.245000 139.160000 38.435000 158.870000 ;
      RECT 37.245000 162.160000 38.435000 181.870000 ;
      RECT 37.245000 185.160000 38.435000 195.010000 ;
      RECT 37.315000  29.780000 37.485000  36.570000 ;
      RECT 37.385000 195.010000 38.275000 195.030000 ;
      RECT 38.095000  29.775000 38.265000  36.570000 ;
      RECT 38.330000   4.820000 38.560000   7.770000 ;
      RECT 38.330000  11.040000 38.560000  13.990000 ;
      RECT 38.330000  17.260000 38.560000  20.210000 ;
      RECT 38.350000   3.755000 38.520000   4.820000 ;
      RECT 38.350000   7.770000 38.520000   8.505000 ;
      RECT 38.350000   9.975000 38.520000  11.040000 ;
      RECT 38.350000  13.990000 38.520000  14.725000 ;
      RECT 38.350000  16.195000 38.520000  17.260000 ;
      RECT 38.350000  20.210000 38.520000  20.945000 ;
      RECT 38.780000 195.370000 39.490000 195.540000 ;
      RECT 38.875000  29.780000 39.045000  36.570000 ;
      RECT 39.060000   4.820000 39.290000   8.825000 ;
      RECT 39.060000  11.040000 39.290000  15.045000 ;
      RECT 39.060000  17.260000 39.290000  21.265000 ;
      RECT 39.090000   2.835000 39.260000   4.820000 ;
      RECT 39.090000   9.055000 39.260000  11.040000 ;
      RECT 39.090000  15.275000 39.260000  17.260000 ;
      RECT 39.260000   2.605000 48.850000   2.635000 ;
      RECT 39.655000  29.770000 39.825000  36.570000 ;
      RECT 39.795000   4.820000 40.025000   7.770000 ;
      RECT 39.795000  11.040000 40.025000  13.990000 ;
      RECT 39.795000  17.260000 40.025000  20.210000 ;
      RECT 39.830000   3.755000 40.000000   4.820000 ;
      RECT 39.830000   7.770000 40.000000   8.505000 ;
      RECT 39.830000   9.975000 40.000000  11.040000 ;
      RECT 39.830000  13.990000 40.000000  14.725000 ;
      RECT 39.830000  16.195000 40.000000  17.260000 ;
      RECT 39.830000  20.210000 40.000000  20.945000 ;
      RECT 39.865000  47.525000 40.395000  65.695000 ;
      RECT 39.865000  70.525000 40.395000  88.695000 ;
      RECT 39.865000  93.525000 40.395000 111.695000 ;
      RECT 39.865000 116.525000 40.395000 134.695000 ;
      RECT 39.865000 139.525000 40.395000 157.695000 ;
      RECT 39.865000 162.525000 40.395000 180.695000 ;
      RECT 39.865000 185.525000 40.395000 195.055000 ;
      RECT 39.885000  47.325000 40.395000  47.525000 ;
      RECT 39.885000  65.695000 40.395000  67.035000 ;
      RECT 39.885000  70.325000 40.395000  70.525000 ;
      RECT 39.885000  88.695000 40.395000  90.035000 ;
      RECT 39.885000  93.325000 40.395000  93.525000 ;
      RECT 39.885000 111.695000 40.395000 113.035000 ;
      RECT 39.885000 116.325000 40.395000 116.525000 ;
      RECT 39.885000 134.695000 40.395000 136.035000 ;
      RECT 39.885000 139.325000 40.395000 139.525000 ;
      RECT 39.885000 157.695000 40.395000 159.035000 ;
      RECT 39.885000 162.325000 40.395000 162.525000 ;
      RECT 39.885000 180.695000 40.395000 182.035000 ;
      RECT 39.885000 185.325000 40.395000 185.525000 ;
      RECT 40.055000   3.075000 48.055000   3.305000 ;
      RECT 40.055000   9.295000 48.055000   9.525000 ;
      RECT 40.055000  15.515000 48.055000  15.745000 ;
      RECT 40.435000  29.780000 40.605000  36.570000 ;
      RECT 40.790000 195.370000 41.500000 195.540000 ;
      RECT 41.215000  29.770000 41.385000  36.570000 ;
      RECT 41.845000  47.160000 43.035000  66.870000 ;
      RECT 41.845000  70.160000 43.035000  89.870000 ;
      RECT 41.845000  93.160000 43.035000 112.870000 ;
      RECT 41.845000 116.160000 43.035000 135.870000 ;
      RECT 41.845000 139.160000 43.035000 158.870000 ;
      RECT 41.845000 162.160000 43.035000 181.870000 ;
      RECT 41.845000 185.160000 43.035000 195.010000 ;
      RECT 41.985000 195.010000 42.875000 195.030000 ;
      RECT 41.995000  29.780000 42.165000  36.570000 ;
      RECT 42.775000  29.775000 42.945000  36.570000 ;
      RECT 43.380000 195.370000 44.090000 195.540000 ;
      RECT 43.555000  29.780000 43.725000  36.570000 ;
      RECT 44.335000  29.770000 44.505000  36.570000 ;
      RECT 44.465000  47.525000 44.995000  65.695000 ;
      RECT 44.465000  70.525000 44.995000  88.695000 ;
      RECT 44.465000  93.525000 44.995000 111.695000 ;
      RECT 44.465000 116.525000 44.995000 134.695000 ;
      RECT 44.465000 139.525000 44.995000 157.695000 ;
      RECT 44.465000 162.525000 44.995000 180.695000 ;
      RECT 44.465000 185.525000 44.995000 195.055000 ;
      RECT 44.485000  47.325000 44.995000  47.525000 ;
      RECT 44.485000  65.695000 44.995000  67.035000 ;
      RECT 44.485000  70.325000 44.995000  70.525000 ;
      RECT 44.485000  88.695000 44.995000  90.035000 ;
      RECT 44.485000  93.325000 44.995000  93.525000 ;
      RECT 44.485000 111.695000 44.995000 113.035000 ;
      RECT 44.485000 116.325000 44.995000 116.525000 ;
      RECT 44.485000 134.695000 44.995000 136.035000 ;
      RECT 44.485000 139.325000 44.995000 139.525000 ;
      RECT 44.485000 157.695000 44.995000 159.035000 ;
      RECT 44.485000 162.325000 44.995000 162.525000 ;
      RECT 44.485000 180.695000 44.995000 182.035000 ;
      RECT 44.485000 185.325000 44.995000 185.525000 ;
      RECT 45.115000  29.780000 45.285000  36.570000 ;
      RECT 45.390000 195.370000 46.100000 195.540000 ;
      RECT 45.755000  29.430000 45.955000  37.425000 ;
      RECT 46.445000  47.160000 47.635000  66.870000 ;
      RECT 46.445000  70.160000 47.635000  89.870000 ;
      RECT 46.445000  93.160000 47.635000 112.870000 ;
      RECT 46.445000 116.160000 47.635000 135.870000 ;
      RECT 46.445000 139.160000 47.635000 158.870000 ;
      RECT 46.445000 162.160000 47.635000 181.870000 ;
      RECT 46.445000 185.160000 47.635000 195.010000 ;
      RECT 46.585000 195.010000 47.475000 195.030000 ;
      RECT 47.310000  28.030000 48.200000  29.215000 ;
      RECT 47.310000  29.525000 48.200000  38.695000 ;
      RECT 47.330000  29.215000 48.180000  29.525000 ;
      RECT 47.980000 195.370000 48.690000 195.540000 ;
      RECT 48.090000   4.820000 48.320000   7.770000 ;
      RECT 48.090000  11.040000 48.320000  13.990000 ;
      RECT 48.090000  17.260000 48.320000  20.210000 ;
      RECT 48.110000   3.755000 48.280000   4.820000 ;
      RECT 48.110000   7.770000 48.280000   8.505000 ;
      RECT 48.110000   9.975000 48.280000  11.040000 ;
      RECT 48.110000  13.990000 48.280000  14.725000 ;
      RECT 48.110000  16.195000 48.280000  17.260000 ;
      RECT 48.110000  20.210000 48.280000  20.945000 ;
      RECT 48.820000   4.820000 49.050000   8.825000 ;
      RECT 48.820000  11.040000 49.050000  15.045000 ;
      RECT 48.820000  17.260000 49.050000  21.265000 ;
      RECT 48.850000   2.835000 49.020000   4.820000 ;
      RECT 48.850000   9.055000 49.020000  11.040000 ;
      RECT 48.850000  15.275000 49.020000  17.260000 ;
      RECT 49.020000   2.605000 58.610000   2.635000 ;
      RECT 49.065000  47.525000 49.595000  65.695000 ;
      RECT 49.065000  70.525000 49.595000  88.695000 ;
      RECT 49.065000  93.525000 49.595000 111.695000 ;
      RECT 49.065000 116.525000 49.595000 134.695000 ;
      RECT 49.065000 139.525000 49.595000 157.695000 ;
      RECT 49.065000 162.525000 49.595000 180.695000 ;
      RECT 49.065000 185.525000 49.595000 195.055000 ;
      RECT 49.085000  47.325000 49.595000  47.525000 ;
      RECT 49.085000  65.695000 49.595000  67.035000 ;
      RECT 49.085000  70.325000 49.595000  70.525000 ;
      RECT 49.085000  88.695000 49.595000  90.035000 ;
      RECT 49.085000  93.325000 49.595000  93.525000 ;
      RECT 49.085000 111.695000 49.595000 113.035000 ;
      RECT 49.085000 116.325000 49.595000 116.525000 ;
      RECT 49.085000 134.695000 49.595000 136.035000 ;
      RECT 49.085000 139.325000 49.595000 139.525000 ;
      RECT 49.085000 157.695000 49.595000 159.035000 ;
      RECT 49.085000 162.325000 49.595000 162.525000 ;
      RECT 49.085000 180.695000 49.595000 182.035000 ;
      RECT 49.085000 185.325000 49.595000 185.525000 ;
      RECT 49.555000   4.820000 49.785000   7.770000 ;
      RECT 49.555000  11.040000 49.785000  13.990000 ;
      RECT 49.555000  17.260000 49.785000  20.210000 ;
      RECT 49.590000   3.755000 49.760000   4.820000 ;
      RECT 49.590000   7.770000 49.760000   8.505000 ;
      RECT 49.590000   9.975000 49.760000  11.040000 ;
      RECT 49.590000  13.990000 49.760000  14.725000 ;
      RECT 49.590000  16.195000 49.760000  17.260000 ;
      RECT 49.590000  20.210000 49.760000  20.945000 ;
      RECT 49.815000   3.075000 57.815000   3.305000 ;
      RECT 49.815000   9.295000 57.815000   9.525000 ;
      RECT 49.815000  15.515000 57.815000  15.745000 ;
      RECT 49.990000 195.370000 50.700000 195.540000 ;
      RECT 51.045000  47.160000 52.235000  66.870000 ;
      RECT 51.045000  70.160000 52.235000  89.870000 ;
      RECT 51.045000  93.160000 52.235000 112.870000 ;
      RECT 51.045000 116.160000 52.235000 135.870000 ;
      RECT 51.045000 139.160000 52.235000 158.870000 ;
      RECT 51.045000 162.160000 52.235000 181.870000 ;
      RECT 51.045000 185.160000 52.235000 195.010000 ;
      RECT 51.185000 195.010000 52.075000 195.030000 ;
      RECT 52.320000  29.300000 68.865000  31.060000 ;
      RECT 52.320000  31.060000 53.210000  41.455000 ;
      RECT 52.320000  41.455000 68.865000  42.495000 ;
      RECT 52.580000 195.370000 53.290000 195.540000 ;
      RECT 53.665000  47.525000 54.195000  65.695000 ;
      RECT 53.665000  70.525000 54.195000  88.695000 ;
      RECT 53.665000  93.525000 54.195000 111.695000 ;
      RECT 53.665000 116.525000 54.195000 134.695000 ;
      RECT 53.665000 139.525000 54.195000 157.695000 ;
      RECT 53.665000 162.525000 54.195000 180.695000 ;
      RECT 53.665000 185.525000 54.195000 195.055000 ;
      RECT 53.685000  47.325000 54.195000  47.525000 ;
      RECT 53.685000  65.695000 54.195000  67.035000 ;
      RECT 53.685000  70.325000 54.195000  70.525000 ;
      RECT 53.685000  88.695000 54.195000  90.035000 ;
      RECT 53.685000  93.325000 54.195000  93.525000 ;
      RECT 53.685000 111.695000 54.195000 113.035000 ;
      RECT 53.685000 116.325000 54.195000 116.525000 ;
      RECT 53.685000 134.695000 54.195000 136.035000 ;
      RECT 53.685000 139.325000 54.195000 139.525000 ;
      RECT 53.685000 157.695000 54.195000 159.035000 ;
      RECT 53.685000 162.325000 54.195000 162.525000 ;
      RECT 53.685000 180.695000 54.195000 182.035000 ;
      RECT 53.685000 185.325000 54.195000 185.525000 ;
      RECT 53.960000  31.835000 67.140000  32.005000 ;
      RECT 53.960000  32.005000 54.130000  40.410000 ;
      RECT 53.960000  40.410000 67.140000  40.580000 ;
      RECT 54.590000 195.370000 55.300000 195.540000 ;
      RECT 54.690000  32.560000 54.860000  36.190000 ;
      RECT 54.690000  36.190000 54.865000  39.290000 ;
      RECT 54.690000  39.290000 54.860000  39.350000 ;
      RECT 54.940000  39.770000 66.335000  39.940000 ;
      RECT 55.215000  23.240000 56.105000  28.345000 ;
      RECT 55.215000  28.345000 70.630000  29.300000 ;
      RECT 55.465000  32.620000 55.640000  35.770000 ;
      RECT 55.470000  32.560000 55.640000  32.620000 ;
      RECT 55.470000  35.770000 55.640000  39.350000 ;
      RECT 55.645000  47.160000 56.835000  66.870000 ;
      RECT 55.645000  70.160000 56.835000  89.870000 ;
      RECT 55.645000  93.160000 56.835000 112.870000 ;
      RECT 55.645000 116.160000 56.835000 135.870000 ;
      RECT 55.645000 139.160000 56.835000 158.870000 ;
      RECT 55.645000 162.160000 56.835000 181.870000 ;
      RECT 55.645000 185.160000 56.835000 195.010000 ;
      RECT 55.785000 195.010000 56.675000 195.140000 ;
      RECT 56.250000  32.560000 56.420000  36.190000 ;
      RECT 56.250000  36.190000 56.425000  39.290000 ;
      RECT 56.250000  39.290000 56.420000  39.350000 ;
      RECT 56.820000  23.480000 57.050000  27.485000 ;
      RECT 56.820000  27.485000 68.570000  27.715000 ;
      RECT 56.850000  21.495000 57.020000  23.480000 ;
      RECT 57.025000  32.620000 57.200000  35.770000 ;
      RECT 57.030000  32.560000 57.200000  32.620000 ;
      RECT 57.030000  35.770000 57.200000  39.350000 ;
      RECT 57.180000 195.370000 57.890000 195.540000 ;
      RECT 57.555000  23.480000 57.785000  26.430000 ;
      RECT 57.590000  22.415000 57.760000  23.480000 ;
      RECT 57.590000  26.430000 57.760000  27.165000 ;
      RECT 57.810000  32.560000 57.980000  36.190000 ;
      RECT 57.810000  36.190000 57.985000  39.290000 ;
      RECT 57.810000  39.290000 57.980000  39.350000 ;
      RECT 57.815000  21.735000 61.815000  21.965000 ;
      RECT 57.850000   4.820000 58.080000   7.770000 ;
      RECT 57.850000  11.040000 58.080000  13.990000 ;
      RECT 57.850000  17.260000 58.080000  20.210000 ;
      RECT 57.870000   3.755000 58.040000   4.820000 ;
      RECT 57.870000   7.770000 58.040000   8.505000 ;
      RECT 57.870000   9.975000 58.040000  11.040000 ;
      RECT 57.870000  13.990000 58.040000  14.725000 ;
      RECT 57.870000  16.195000 58.040000  17.260000 ;
      RECT 57.870000  20.210000 58.040000  20.945000 ;
      RECT 58.265000  47.525000 58.795000  65.695000 ;
      RECT 58.265000  70.525000 58.795000  88.695000 ;
      RECT 58.265000  93.525000 58.795000 111.695000 ;
      RECT 58.265000 116.525000 58.795000 134.695000 ;
      RECT 58.265000 139.525000 58.795000 157.695000 ;
      RECT 58.265000 162.525000 58.795000 180.695000 ;
      RECT 58.265000 185.525000 58.795000 195.055000 ;
      RECT 58.285000  47.325000 58.795000  47.525000 ;
      RECT 58.285000  65.695000 58.795000  67.035000 ;
      RECT 58.285000  70.325000 58.795000  70.525000 ;
      RECT 58.285000  88.695000 58.795000  90.035000 ;
      RECT 58.285000  93.325000 58.795000  93.525000 ;
      RECT 58.285000 111.695000 58.795000 113.035000 ;
      RECT 58.285000 116.325000 58.795000 116.525000 ;
      RECT 58.285000 134.695000 58.795000 136.035000 ;
      RECT 58.285000 139.325000 58.795000 139.525000 ;
      RECT 58.285000 157.695000 58.795000 159.035000 ;
      RECT 58.285000 162.325000 58.795000 162.525000 ;
      RECT 58.285000 180.695000 58.795000 182.035000 ;
      RECT 58.285000 185.325000 58.795000 185.525000 ;
      RECT 58.580000   4.820000 58.810000   8.825000 ;
      RECT 58.580000  11.040000 58.810000  15.045000 ;
      RECT 58.580000  17.260000 58.810000  21.265000 ;
      RECT 58.585000  32.620000 58.760000  35.770000 ;
      RECT 58.590000  32.560000 58.760000  32.620000 ;
      RECT 58.590000  35.770000 58.760000  39.350000 ;
      RECT 58.610000   2.835000 58.780000   4.820000 ;
      RECT 58.610000   9.055000 58.780000  11.040000 ;
      RECT 58.610000  15.275000 58.780000  17.260000 ;
      RECT 58.780000   2.605000 68.370000   2.635000 ;
      RECT 59.190000 195.370000 59.900000 195.540000 ;
      RECT 59.315000   4.820000 59.545000   7.770000 ;
      RECT 59.315000  11.040000 59.545000  13.990000 ;
      RECT 59.315000  17.260000 59.545000  20.210000 ;
      RECT 59.350000   3.755000 59.520000   4.820000 ;
      RECT 59.350000   7.770000 59.520000   8.505000 ;
      RECT 59.350000   9.975000 59.520000  11.040000 ;
      RECT 59.350000  13.990000 59.520000  14.725000 ;
      RECT 59.350000  16.195000 59.520000  17.260000 ;
      RECT 59.350000  20.210000 59.520000  20.945000 ;
      RECT 59.370000  32.560000 59.540000  36.190000 ;
      RECT 59.370000  36.190000 59.545000  39.290000 ;
      RECT 59.370000  39.290000 59.540000  39.350000 ;
      RECT 59.575000   3.075000 67.575000   3.305000 ;
      RECT 59.575000   9.295000 67.575000   9.525000 ;
      RECT 59.575000  15.515000 67.575000  15.745000 ;
      RECT 60.145000  32.620000 60.320000  35.770000 ;
      RECT 60.150000  32.560000 60.320000  32.620000 ;
      RECT 60.150000  35.770000 60.320000  39.350000 ;
      RECT 60.245000  47.160000 61.435000  66.870000 ;
      RECT 60.245000  70.160000 61.435000  89.870000 ;
      RECT 60.245000  93.160000 61.435000 112.870000 ;
      RECT 60.245000 116.160000 61.435000 135.870000 ;
      RECT 60.245000 139.160000 61.435000 158.870000 ;
      RECT 60.245000 162.160000 61.435000 181.870000 ;
      RECT 60.245000 185.160000 61.435000 195.010000 ;
      RECT 60.385000 195.010000 61.275000 195.140000 ;
      RECT 60.930000  32.560000 61.100000  36.190000 ;
      RECT 60.930000  36.190000 61.105000  39.290000 ;
      RECT 60.930000  39.290000 61.100000  39.350000 ;
      RECT 61.705000  32.620000 61.880000  35.770000 ;
      RECT 61.710000  32.560000 61.880000  32.620000 ;
      RECT 61.710000  35.770000 61.880000  39.350000 ;
      RECT 61.780000 195.370000 62.490000 195.540000 ;
      RECT 61.850000  23.480000 62.080000  26.430000 ;
      RECT 61.870000  22.415000 62.040000  23.480000 ;
      RECT 61.870000  26.430000 62.040000  27.165000 ;
      RECT 62.490000  32.560000 62.660000  36.190000 ;
      RECT 62.490000  36.190000 62.665000  39.290000 ;
      RECT 62.490000  39.290000 62.660000  39.350000 ;
      RECT 62.580000  23.480000 62.810000  27.485000 ;
      RECT 62.610000  21.495000 62.780000  23.480000 ;
      RECT 62.865000  47.525000 63.395000  65.695000 ;
      RECT 62.865000  70.525000 63.395000  88.695000 ;
      RECT 62.865000  93.525000 63.395000 111.695000 ;
      RECT 62.865000 116.525000 63.395000 134.695000 ;
      RECT 62.865000 139.525000 63.395000 157.695000 ;
      RECT 62.865000 162.525000 63.395000 180.695000 ;
      RECT 62.865000 185.525000 63.395000 195.055000 ;
      RECT 62.885000  47.325000 63.395000  47.525000 ;
      RECT 62.885000  65.695000 63.395000  67.035000 ;
      RECT 62.885000  70.325000 63.395000  70.525000 ;
      RECT 62.885000  88.695000 63.395000  90.035000 ;
      RECT 62.885000  93.325000 63.395000  93.525000 ;
      RECT 62.885000 111.695000 63.395000 113.035000 ;
      RECT 62.885000 116.325000 63.395000 116.525000 ;
      RECT 62.885000 134.695000 63.395000 136.035000 ;
      RECT 62.885000 139.325000 63.395000 139.525000 ;
      RECT 62.885000 157.695000 63.395000 159.035000 ;
      RECT 62.885000 162.325000 63.395000 162.525000 ;
      RECT 62.885000 180.695000 63.395000 182.035000 ;
      RECT 62.885000 185.325000 63.395000 185.525000 ;
      RECT 63.265000  32.620000 63.440000  35.770000 ;
      RECT 63.270000  32.560000 63.440000  32.620000 ;
      RECT 63.270000  35.770000 63.440000  39.350000 ;
      RECT 63.315000  23.480000 63.545000  26.430000 ;
      RECT 63.350000  22.415000 63.520000  23.480000 ;
      RECT 63.350000  26.430000 63.520000  27.165000 ;
      RECT 63.575000  21.735000 67.575000  21.965000 ;
      RECT 63.790000 195.370000 64.500000 195.540000 ;
      RECT 64.050000  32.560000 64.220000  36.190000 ;
      RECT 64.050000  36.190000 64.225000  39.290000 ;
      RECT 64.050000  39.290000 64.220000  39.350000 ;
      RECT 64.825000  32.620000 65.000000  35.770000 ;
      RECT 64.830000  32.560000 65.000000  32.620000 ;
      RECT 64.830000  35.770000 65.000000  39.350000 ;
      RECT 64.845000  47.160000 65.875000  66.930000 ;
      RECT 64.845000  70.160000 65.875000  89.930000 ;
      RECT 64.845000  93.160000 65.875000 112.935000 ;
      RECT 64.845000 116.160000 65.875000 135.930000 ;
      RECT 64.845000 139.160000 65.875000 158.930000 ;
      RECT 64.845000 162.160000 65.875000 181.930000 ;
      RECT 64.845000 185.160000 65.875000 195.180000 ;
      RECT 65.610000  32.560000 65.780000  36.190000 ;
      RECT 65.610000  36.190000 65.785000  39.290000 ;
      RECT 65.610000  39.290000 65.780000  39.350000 ;
      RECT 66.385000  32.620000 66.560000  35.770000 ;
      RECT 66.390000  32.560000 66.560000  32.620000 ;
      RECT 66.390000  35.770000 66.560000  39.350000 ;
      RECT 66.935000  32.005000 67.140000  36.065000 ;
      RECT 66.935000  36.275000 67.140000  40.410000 ;
      RECT 66.970000  36.065000 67.140000  36.275000 ;
      RECT 67.265000  46.350000 68.155000 101.315000 ;
      RECT 67.265000 166.045000 68.155000 196.835000 ;
      RECT 67.290000 101.315000 68.140000 101.710000 ;
      RECT 67.290000 101.710000 68.155000 165.645000 ;
      RECT 67.290000 165.645000 68.140000 166.045000 ;
      RECT 67.610000   4.820000 67.840000   7.770000 ;
      RECT 67.610000  11.040000 67.840000  13.990000 ;
      RECT 67.610000  17.260000 67.840000  20.210000 ;
      RECT 67.610000  23.480000 67.840000  26.430000 ;
      RECT 67.630000   3.755000 67.800000   4.820000 ;
      RECT 67.630000   7.770000 67.800000   8.505000 ;
      RECT 67.630000   9.975000 67.800000  11.040000 ;
      RECT 67.630000  13.990000 67.800000  14.725000 ;
      RECT 67.630000  16.195000 67.800000  17.260000 ;
      RECT 67.630000  20.210000 67.800000  20.945000 ;
      RECT 67.630000  22.415000 67.800000  23.480000 ;
      RECT 67.630000  26.430000 67.800000  27.165000 ;
      RECT 67.975000  31.060000 68.865000  40.480000 ;
      RECT 67.975000  41.315000 68.865000  41.455000 ;
      RECT 68.000000  40.480000 68.830000  41.315000 ;
      RECT 68.340000   4.820000 68.570000   8.825000 ;
      RECT 68.340000  11.040000 68.570000  15.045000 ;
      RECT 68.340000  17.260000 68.570000  21.265000 ;
      RECT 68.340000  23.480000 68.570000  27.485000 ;
      RECT 68.370000   2.835000 68.540000   4.820000 ;
      RECT 68.370000   9.055000 68.540000  11.040000 ;
      RECT 68.370000  15.275000 68.540000  17.260000 ;
      RECT 68.370000  21.495000 68.540000  23.480000 ;
      RECT 68.875000  44.755000 70.125000  45.995000 ;
      RECT 68.875000  46.185000 70.125000 198.445000 ;
      RECT 68.905000  45.995000 70.095000  46.185000 ;
      RECT 69.740000  22.520000 70.630000  28.345000 ;
      RECT 69.760000   1.890000 70.650000   2.770000 ;
      RECT 69.765000   3.845000 70.630000   8.915000 ;
      RECT 69.765000   9.845000 70.630000  14.915000 ;
      RECT 69.765000  16.165000 70.630000  21.235000 ;
      RECT 69.780000   2.770000 70.630000   3.845000 ;
      RECT 69.780000   8.915000 70.630000   9.845000 ;
      RECT 69.780000  14.915000 70.630000  16.165000 ;
      RECT 69.780000  21.235000 70.630000  22.520000 ;
      RECT 70.470000  42.820000 71.055000  42.990000 ;
      RECT 70.725000  42.735000 71.055000  42.820000 ;
      RECT 70.725000  42.990000 71.055000  43.015000 ;
      RECT 72.245000 199.210000 72.775000 199.380000 ;
      RECT 72.345000 199.380000 72.675000 199.420000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  0.215000   2.170000 ;
      RECT  0.000000   0.000000  0.215000   2.170000 ;
      RECT  0.000000   2.170000  0.215000   2.240000 ;
      RECT  0.000000   2.170000  0.725000   2.680000 ;
      RECT  0.000000   2.240000  0.285000   2.310000 ;
      RECT  0.000000   2.310000  0.355000   2.380000 ;
      RECT  0.000000   2.380000  0.425000   2.450000 ;
      RECT  0.000000   2.450000  0.495000   2.520000 ;
      RECT  0.000000   2.520000  0.565000   2.590000 ;
      RECT  0.000000   2.590000  0.635000   2.660000 ;
      RECT  0.000000   2.660000  0.705000   2.680000 ;
      RECT  0.000000   2.680000  0.725000  36.970000 ;
      RECT  0.000000   2.680000  0.725000  36.970000 ;
      RECT  0.000000  36.970000  0.725000  37.015000 ;
      RECT  0.000000  36.970000  0.810000  37.055000 ;
      RECT  0.000000  37.015000  0.770000  37.055000 ;
      RECT  0.000000  37.055000  0.810000  46.900000 ;
      RECT  0.000000  37.055000  0.810000  46.900000 ;
      RECT  0.000000  46.900000  0.725000  46.985000 ;
      RECT  0.000000  46.900000  0.770000  46.940000 ;
      RECT  0.000000  46.940000  0.730000  46.980000 ;
      RECT  0.000000  46.980000  0.725000  46.985000 ;
      RECT  0.000000  46.985000  0.725000 195.355000 ;
      RECT  0.000000  46.985000  0.725000 195.355000 ;
      RECT  0.000000 195.355000 67.480000 200.000000 ;
      RECT  0.000000 195.355000 75.000000 200.000000 ;
      RECT 14.400000  45.430000 57.415000  47.315000 ;
      RECT 14.400000  45.430000 59.035000  45.500000 ;
      RECT 14.400000  45.430000 59.035000  45.500000 ;
      RECT 14.400000  45.500000 58.965000  45.570000 ;
      RECT 14.400000  45.500000 58.965000  45.570000 ;
      RECT 14.400000  45.570000 58.895000  45.640000 ;
      RECT 14.400000  45.570000 58.895000  45.640000 ;
      RECT 14.400000  45.640000 58.825000  45.710000 ;
      RECT 14.400000  45.640000 58.825000  45.710000 ;
      RECT 14.400000  45.710000 58.755000  45.780000 ;
      RECT 14.400000  45.710000 58.755000  45.780000 ;
      RECT 14.400000  45.780000 58.685000  45.850000 ;
      RECT 14.400000  45.780000 58.685000  45.850000 ;
      RECT 14.400000  45.850000 58.615000  45.920000 ;
      RECT 14.400000  45.850000 58.615000  45.920000 ;
      RECT 14.400000  45.920000 58.545000  45.990000 ;
      RECT 14.400000  45.920000 58.545000  45.990000 ;
      RECT 14.400000  45.990000 58.475000  46.060000 ;
      RECT 14.400000  45.990000 58.475000  46.060000 ;
      RECT 14.400000  46.060000 58.405000  46.130000 ;
      RECT 14.400000  46.060000 58.405000  46.130000 ;
      RECT 14.400000  46.130000 58.335000  46.200000 ;
      RECT 14.400000  46.130000 58.335000  46.200000 ;
      RECT 14.400000  46.200000 58.265000  46.270000 ;
      RECT 14.400000  46.200000 58.265000  46.270000 ;
      RECT 14.400000  46.270000 58.195000  46.340000 ;
      RECT 14.400000  46.270000 58.195000  46.340000 ;
      RECT 14.400000  46.340000 58.125000  46.410000 ;
      RECT 14.400000  46.340000 58.125000  46.410000 ;
      RECT 14.400000  46.410000 58.055000  46.480000 ;
      RECT 14.400000  46.410000 58.055000  46.480000 ;
      RECT 14.400000  46.480000 57.985000  46.550000 ;
      RECT 14.400000  46.480000 57.985000  46.550000 ;
      RECT 14.400000  46.550000 57.915000  46.620000 ;
      RECT 14.400000  46.550000 57.915000  46.620000 ;
      RECT 14.400000  46.620000 57.845000  46.690000 ;
      RECT 14.400000  46.620000 57.845000  46.690000 ;
      RECT 14.400000  46.690000 57.775000  46.760000 ;
      RECT 14.400000  46.690000 57.775000  46.760000 ;
      RECT 14.400000  46.760000 57.705000  46.830000 ;
      RECT 14.400000  46.760000 57.705000  46.830000 ;
      RECT 14.400000  46.830000 57.635000  46.900000 ;
      RECT 14.400000  46.830000 57.635000  46.900000 ;
      RECT 14.400000  46.900000 57.565000  46.970000 ;
      RECT 14.400000  46.900000 57.565000  46.970000 ;
      RECT 14.400000  46.970000 57.495000  47.040000 ;
      RECT 14.400000  46.970000 57.495000  47.040000 ;
      RECT 14.400000  47.040000 57.425000  47.110000 ;
      RECT 14.400000  47.040000 57.425000  47.110000 ;
      RECT 14.400000  47.110000 57.360000  47.175000 ;
      RECT 14.400000  47.110000 57.360000  47.175000 ;
      RECT 14.400000  47.175000 16.525000  54.100000 ;
      RECT 14.400000  47.315000 16.665000  54.100000 ;
      RECT 14.400000  54.100000 16.665000  54.905000 ;
      RECT 14.400000  70.140000 57.405000  70.160000 ;
      RECT 14.400000  70.140000 57.405000  70.160000 ;
      RECT 14.400000  70.140000 57.445000  70.315000 ;
      RECT 14.400000  70.160000 57.390000  70.175000 ;
      RECT 14.400000  70.160000 57.390000  70.175000 ;
      RECT 14.400000  70.175000 24.540000  72.870000 ;
      RECT 14.400000  70.315000 24.680000  72.925000 ;
      RECT 14.400000  72.870000 24.470000  72.940000 ;
      RECT 14.400000  72.870000 24.470000  72.940000 ;
      RECT 14.400000  72.925000 23.590000  74.015000 ;
      RECT 14.400000  72.940000 24.400000  73.010000 ;
      RECT 14.400000  72.940000 24.400000  73.010000 ;
      RECT 14.400000  73.010000 24.330000  73.080000 ;
      RECT 14.400000  73.010000 24.330000  73.080000 ;
      RECT 14.400000  73.080000 24.260000  73.150000 ;
      RECT 14.400000  73.080000 24.260000  73.150000 ;
      RECT 14.400000  73.150000 24.190000  73.220000 ;
      RECT 14.400000  73.150000 24.190000  73.220000 ;
      RECT 14.400000  73.220000 24.120000  73.290000 ;
      RECT 14.400000  73.220000 24.120000  73.290000 ;
      RECT 14.400000  73.290000 24.050000  73.360000 ;
      RECT 14.400000  73.290000 24.050000  73.360000 ;
      RECT 14.400000  73.360000 23.980000  73.430000 ;
      RECT 14.400000  73.360000 23.980000  73.430000 ;
      RECT 14.400000  73.430000 23.910000  73.500000 ;
      RECT 14.400000  73.430000 23.910000  73.500000 ;
      RECT 14.400000  73.500000 23.840000  73.570000 ;
      RECT 14.400000  73.500000 23.840000  73.570000 ;
      RECT 14.400000  73.570000 23.770000  73.640000 ;
      RECT 14.400000  73.570000 23.770000  73.640000 ;
      RECT 14.400000  73.640000 23.700000  73.710000 ;
      RECT 14.400000  73.640000 23.700000  73.710000 ;
      RECT 14.400000  73.710000 23.630000  73.780000 ;
      RECT 14.400000  73.710000 23.630000  73.780000 ;
      RECT 14.400000  73.780000 23.560000  73.850000 ;
      RECT 14.400000  73.780000 23.560000  73.850000 ;
      RECT 14.400000  73.850000 23.535000  73.875000 ;
      RECT 14.400000  73.850000 23.535000  73.875000 ;
      RECT 14.400000  73.875000 18.130000  74.695000 ;
      RECT 14.400000  74.015000 18.270000  74.555000 ;
      RECT 14.400000  74.555000 24.680000  75.675000 ;
      RECT 14.400000  74.695000 23.505000  74.765000 ;
      RECT 14.400000  74.695000 23.505000  74.765000 ;
      RECT 14.400000  74.765000 23.575000  74.835000 ;
      RECT 14.400000  74.765000 23.575000  74.835000 ;
      RECT 14.400000  74.835000 23.645000  74.905000 ;
      RECT 14.400000  74.835000 23.645000  74.905000 ;
      RECT 14.400000  74.905000 23.715000  74.975000 ;
      RECT 14.400000  74.905000 23.715000  74.975000 ;
      RECT 14.400000  74.975000 23.785000  75.045000 ;
      RECT 14.400000  74.975000 23.785000  75.045000 ;
      RECT 14.400000  75.045000 23.855000  75.115000 ;
      RECT 14.400000  75.045000 23.855000  75.115000 ;
      RECT 14.400000  75.115000 23.925000  75.185000 ;
      RECT 14.400000  75.115000 23.925000  75.185000 ;
      RECT 14.400000  75.185000 23.995000  75.255000 ;
      RECT 14.400000  75.185000 23.995000  75.255000 ;
      RECT 14.400000  75.255000 24.065000  75.325000 ;
      RECT 14.400000  75.255000 24.065000  75.325000 ;
      RECT 14.400000  75.325000 24.135000  75.395000 ;
      RECT 14.400000  75.325000 24.135000  75.395000 ;
      RECT 14.400000  75.395000 24.205000  75.465000 ;
      RECT 14.400000  75.395000 24.205000  75.465000 ;
      RECT 14.400000  75.465000 24.275000  75.535000 ;
      RECT 14.400000  75.465000 24.275000  75.535000 ;
      RECT 14.400000  75.535000 24.345000  75.605000 ;
      RECT 14.400000  75.535000 24.345000  75.605000 ;
      RECT 14.400000  75.605000 24.415000  75.675000 ;
      RECT 14.400000  75.605000 24.415000  75.675000 ;
      RECT 14.400000  75.675000 24.485000  75.730000 ;
      RECT 14.400000  75.675000 24.485000  75.730000 ;
      RECT 14.400000  75.675000 24.680000  77.125000 ;
      RECT 14.400000  75.730000 24.540000  77.125000 ;
      RECT 14.400000  77.125000 24.680000  79.295000 ;
      RECT 14.400000  93.140000 57.465000  93.160000 ;
      RECT 14.400000  93.140000 57.465000  93.160000 ;
      RECT 14.400000  93.140000 57.505000  93.315000 ;
      RECT 14.400000  93.160000 57.450000  93.175000 ;
      RECT 14.400000  93.160000 57.450000  93.175000 ;
      RECT 14.400000  93.175000 24.540000 100.125000 ;
      RECT 14.400000  93.315000 24.680000 100.125000 ;
      RECT 14.400000 100.125000 24.680000 102.295000 ;
      RECT 14.400000 116.180000 24.540000 123.030000 ;
      RECT 14.400000 116.180000 57.415000 116.315000 ;
      RECT 14.400000 116.315000 24.680000 123.030000 ;
      RECT 14.400000 123.030000 24.680000 125.295000 ;
      RECT 14.400000 139.285000 16.525000 146.100000 ;
      RECT 14.400000 139.285000 57.450000 139.315000 ;
      RECT 14.400000 139.315000 16.665000 146.100000 ;
      RECT 14.400000 146.100000 16.665000 146.770000 ;
      RECT 14.400000 162.195000 16.525000 169.105000 ;
      RECT 14.400000 162.195000 57.465000 162.315000 ;
      RECT 14.400000 162.315000 16.665000 169.105000 ;
      RECT 14.400000 169.105000 16.665000 171.295000 ;
      RECT 14.400000 185.170000 15.340000 189.470000 ;
      RECT 14.400000 185.170000 15.480000 189.470000 ;
      RECT 14.400000 189.470000 15.480000 190.155000 ;
      RECT 14.405000 116.175000 24.540000 116.180000 ;
      RECT 14.405000 116.175000 24.540000 116.180000 ;
      RECT 14.410000 162.185000 16.525000 162.195000 ;
      RECT 14.415000 185.155000 15.340000 185.170000 ;
      RECT 14.415000 185.155000 15.480000 185.170000 ;
      RECT 14.420000  70.120000 57.425000  70.140000 ;
      RECT 14.420000  70.120000 57.425000  70.140000 ;
      RECT 14.420000 162.175000 16.525000 162.185000 ;
      RECT 14.445000  45.385000 59.105000  45.430000 ;
      RECT 14.445000  45.385000 59.105000  45.430000 ;
      RECT 14.455000  93.085000 57.485000  93.140000 ;
      RECT 14.455000  93.085000 57.485000  93.140000 ;
      RECT 14.455000 139.230000 16.525000 139.285000 ;
      RECT 14.460000 116.120000 57.360000 116.175000 ;
      RECT 14.460000 116.120000 57.360000 116.175000 ;
      RECT 14.470000  54.100000 16.525000  54.170000 ;
      RECT 14.470000  77.125000 24.540000  77.195000 ;
      RECT 14.470000  77.125000 24.540000  77.195000 ;
      RECT 14.470000 100.125000 24.540000 100.195000 ;
      RECT 14.470000 100.125000 24.540000 100.195000 ;
      RECT 14.470000 123.030000 24.540000 123.100000 ;
      RECT 14.470000 123.030000 24.540000 123.100000 ;
      RECT 14.470000 146.100000 16.525000 146.170000 ;
      RECT 14.470000 169.105000 16.525000 169.175000 ;
      RECT 14.470000 189.470000 15.340000 189.540000 ;
      RECT 14.475000 162.120000 57.410000 162.175000 ;
      RECT 14.475000 162.120000 57.410000 162.175000 ;
      RECT 14.485000 185.085000 15.340000 185.155000 ;
      RECT 14.490000  70.050000 57.445000  70.120000 ;
      RECT 14.490000  70.050000 57.445000  70.120000 ;
      RECT 14.510000 139.175000 16.525000 139.230000 ;
      RECT 14.515000  45.315000 59.150000  45.385000 ;
      RECT 14.515000  45.315000 59.150000  45.385000 ;
      RECT 14.525000  93.015000 57.540000  93.085000 ;
      RECT 14.525000  93.015000 57.540000  93.085000 ;
      RECT 14.530000 116.050000 57.415000 116.120000 ;
      RECT 14.530000 116.050000 57.415000 116.120000 ;
      RECT 14.540000  54.170000 16.525000  54.240000 ;
      RECT 14.540000  77.195000 24.540000  77.265000 ;
      RECT 14.540000  77.195000 24.540000  77.265000 ;
      RECT 14.540000 100.195000 24.540000 100.265000 ;
      RECT 14.540000 100.195000 24.540000 100.265000 ;
      RECT 14.540000 123.100000 24.540000 123.170000 ;
      RECT 14.540000 123.100000 24.540000 123.170000 ;
      RECT 14.540000 146.170000 16.525000 146.240000 ;
      RECT 14.540000 169.175000 16.525000 169.245000 ;
      RECT 14.540000 189.540000 15.340000 189.610000 ;
      RECT 14.545000 162.050000 57.465000 162.120000 ;
      RECT 14.545000 162.050000 57.465000 162.120000 ;
      RECT 14.555000 185.015000 15.340000 185.085000 ;
      RECT 14.560000  69.980000 57.515000  70.050000 ;
      RECT 14.560000  69.980000 57.515000  70.050000 ;
      RECT 14.565000 139.120000 57.395000 139.175000 ;
      RECT 14.565000 139.120000 57.395000 139.175000 ;
      RECT 14.565000 185.005000 58.580000 185.015000 ;
      RECT 14.585000  45.245000 59.220000  45.315000 ;
      RECT 14.585000  45.245000 59.220000  45.315000 ;
      RECT 14.595000  92.945000 57.610000  93.015000 ;
      RECT 14.595000  92.945000 57.610000  93.015000 ;
      RECT 14.600000 115.980000 57.485000 116.050000 ;
      RECT 14.600000 115.980000 57.485000 116.050000 ;
      RECT 14.610000  54.240000 16.525000  54.310000 ;
      RECT 14.610000  77.265000 24.540000  77.335000 ;
      RECT 14.610000  77.265000 24.540000  77.335000 ;
      RECT 14.610000 100.265000 24.540000 100.335000 ;
      RECT 14.610000 100.265000 24.540000 100.335000 ;
      RECT 14.610000 123.170000 24.540000 123.240000 ;
      RECT 14.610000 123.170000 24.540000 123.240000 ;
      RECT 14.610000 146.240000 16.525000 146.310000 ;
      RECT 14.610000 169.245000 16.525000 169.315000 ;
      RECT 14.610000 189.610000 15.340000 189.680000 ;
      RECT 14.615000 161.980000 57.535000 162.050000 ;
      RECT 14.615000 161.980000 57.535000 162.050000 ;
      RECT 14.630000  69.910000 57.585000  69.980000 ;
      RECT 14.630000  69.910000 57.585000  69.980000 ;
      RECT 14.635000 139.050000 57.450000 139.120000 ;
      RECT 14.635000 139.050000 57.450000 139.120000 ;
      RECT 14.635000 184.935000 58.590000 185.005000 ;
      RECT 14.655000  45.175000 59.290000  45.245000 ;
      RECT 14.655000  45.175000 59.290000  45.245000 ;
      RECT 14.665000  92.875000 57.680000  92.945000 ;
      RECT 14.665000  92.875000 57.680000  92.945000 ;
      RECT 14.670000 115.910000 57.555000 115.980000 ;
      RECT 14.670000 115.910000 57.555000 115.980000 ;
      RECT 14.680000  54.310000 16.525000  54.380000 ;
      RECT 14.680000  77.335000 24.540000  77.405000 ;
      RECT 14.680000  77.335000 24.540000  77.405000 ;
      RECT 14.680000 100.335000 24.540000 100.405000 ;
      RECT 14.680000 100.335000 24.540000 100.405000 ;
      RECT 14.680000 123.240000 24.540000 123.310000 ;
      RECT 14.680000 123.240000 24.540000 123.310000 ;
      RECT 14.680000 146.310000 16.525000 146.380000 ;
      RECT 14.680000 169.315000 16.525000 169.385000 ;
      RECT 14.680000 189.680000 15.340000 189.750000 ;
      RECT 14.685000 161.910000 57.605000 161.980000 ;
      RECT 14.685000 161.910000 57.605000 161.980000 ;
      RECT 14.700000  69.840000 57.655000  69.910000 ;
      RECT 14.700000  69.840000 57.655000  69.910000 ;
      RECT 14.705000 138.980000 57.520000 139.050000 ;
      RECT 14.705000 138.980000 57.520000 139.050000 ;
      RECT 14.705000 184.865000 58.660000 184.935000 ;
      RECT 14.725000  45.105000 59.360000  45.175000 ;
      RECT 14.725000  45.105000 59.360000  45.175000 ;
      RECT 14.735000  92.805000 57.750000  92.875000 ;
      RECT 14.735000  92.805000 57.750000  92.875000 ;
      RECT 14.740000 115.840000 57.625000 115.910000 ;
      RECT 14.740000 115.840000 57.625000 115.910000 ;
      RECT 14.750000  54.380000 16.525000  54.450000 ;
      RECT 14.750000  77.405000 24.540000  77.475000 ;
      RECT 14.750000  77.405000 24.540000  77.475000 ;
      RECT 14.750000 100.405000 24.540000 100.475000 ;
      RECT 14.750000 100.405000 24.540000 100.475000 ;
      RECT 14.750000 123.310000 24.540000 123.380000 ;
      RECT 14.750000 123.310000 24.540000 123.380000 ;
      RECT 14.750000 146.380000 16.525000 146.450000 ;
      RECT 14.750000 169.385000 16.525000 169.455000 ;
      RECT 14.750000 189.750000 15.340000 189.820000 ;
      RECT 14.755000 161.840000 57.675000 161.910000 ;
      RECT 14.755000 161.840000 57.675000 161.910000 ;
      RECT 14.770000  69.770000 57.725000  69.840000 ;
      RECT 14.770000  69.770000 57.725000  69.840000 ;
      RECT 14.775000 138.910000 57.590000 138.980000 ;
      RECT 14.775000 138.910000 57.590000 138.980000 ;
      RECT 14.775000 184.795000 58.730000 184.865000 ;
      RECT 14.795000  45.035000 59.430000  45.105000 ;
      RECT 14.795000  45.035000 59.430000  45.105000 ;
      RECT 14.805000  92.735000 57.820000  92.805000 ;
      RECT 14.805000  92.735000 57.820000  92.805000 ;
      RECT 14.810000 115.770000 57.695000 115.840000 ;
      RECT 14.810000 115.770000 57.695000 115.840000 ;
      RECT 14.820000  54.450000 16.525000  54.520000 ;
      RECT 14.820000  77.475000 24.540000  77.545000 ;
      RECT 14.820000  77.475000 24.540000  77.545000 ;
      RECT 14.820000 100.475000 24.540000 100.545000 ;
      RECT 14.820000 100.475000 24.540000 100.545000 ;
      RECT 14.820000 123.380000 24.540000 123.450000 ;
      RECT 14.820000 123.380000 24.540000 123.450000 ;
      RECT 14.820000 146.450000 16.525000 146.520000 ;
      RECT 14.820000 169.455000 16.525000 169.525000 ;
      RECT 14.820000 189.820000 15.340000 189.890000 ;
      RECT 14.825000 161.770000 57.745000 161.840000 ;
      RECT 14.825000 161.770000 57.745000 161.840000 ;
      RECT 14.840000  69.700000 57.795000  69.770000 ;
      RECT 14.840000  69.700000 57.795000  69.770000 ;
      RECT 14.845000 138.840000 57.660000 138.910000 ;
      RECT 14.845000 138.840000 57.660000 138.910000 ;
      RECT 14.845000 184.725000 58.800000 184.795000 ;
      RECT 14.865000  44.965000 59.500000  45.035000 ;
      RECT 14.865000  44.965000 59.500000  45.035000 ;
      RECT 14.875000  92.665000 57.890000  92.735000 ;
      RECT 14.875000  92.665000 57.890000  92.735000 ;
      RECT 14.880000 115.700000 57.765000 115.770000 ;
      RECT 14.880000 115.700000 57.765000 115.770000 ;
      RECT 14.890000  54.520000 16.525000  54.590000 ;
      RECT 14.890000  77.545000 24.540000  77.615000 ;
      RECT 14.890000  77.545000 24.540000  77.615000 ;
      RECT 14.890000 100.545000 24.540000 100.615000 ;
      RECT 14.890000 100.545000 24.540000 100.615000 ;
      RECT 14.890000 123.450000 24.540000 123.520000 ;
      RECT 14.890000 123.450000 24.540000 123.520000 ;
      RECT 14.890000 146.520000 16.525000 146.590000 ;
      RECT 14.890000 169.525000 16.525000 169.595000 ;
      RECT 14.890000 189.890000 15.340000 189.960000 ;
      RECT 14.895000 161.700000 57.815000 161.770000 ;
      RECT 14.895000 161.700000 57.815000 161.770000 ;
      RECT 14.910000  69.630000 57.865000  69.700000 ;
      RECT 14.910000  69.630000 57.865000  69.700000 ;
      RECT 14.915000 138.770000 57.730000 138.840000 ;
      RECT 14.915000 138.770000 57.730000 138.840000 ;
      RECT 14.915000 184.655000 58.870000 184.725000 ;
      RECT 14.935000  44.895000 59.570000  44.965000 ;
      RECT 14.935000  44.895000 59.570000  44.965000 ;
      RECT 14.945000  92.595000 57.960000  92.665000 ;
      RECT 14.945000  92.595000 57.960000  92.665000 ;
      RECT 14.950000 115.630000 57.835000 115.700000 ;
      RECT 14.950000 115.630000 57.835000 115.700000 ;
      RECT 14.960000  54.590000 16.525000  54.660000 ;
      RECT 14.960000  77.615000 24.540000  77.685000 ;
      RECT 14.960000  77.615000 24.540000  77.685000 ;
      RECT 14.960000 100.615000 24.540000 100.685000 ;
      RECT 14.960000 100.615000 24.540000 100.685000 ;
      RECT 14.960000 123.520000 24.540000 123.590000 ;
      RECT 14.960000 123.520000 24.540000 123.590000 ;
      RECT 14.960000 146.590000 16.525000 146.660000 ;
      RECT 14.960000 169.595000 16.525000 169.665000 ;
      RECT 14.960000 189.960000 15.340000 190.030000 ;
      RECT 14.965000 161.630000 57.885000 161.700000 ;
      RECT 14.965000 161.630000 57.885000 161.700000 ;
      RECT 14.980000  69.560000 57.935000  69.630000 ;
      RECT 14.980000  69.560000 57.935000  69.630000 ;
      RECT 14.985000 138.700000 57.800000 138.770000 ;
      RECT 14.985000 138.700000 57.800000 138.770000 ;
      RECT 14.985000 184.585000 58.940000 184.655000 ;
      RECT 15.005000  44.825000 59.640000  44.895000 ;
      RECT 15.005000  44.825000 59.640000  44.895000 ;
      RECT 15.015000  92.525000 58.030000  92.595000 ;
      RECT 15.015000  92.525000 58.030000  92.595000 ;
      RECT 15.020000 115.560000 57.905000 115.630000 ;
      RECT 15.020000 115.560000 57.905000 115.630000 ;
      RECT 15.030000  54.660000 16.525000  54.730000 ;
      RECT 15.030000  77.685000 24.540000  77.755000 ;
      RECT 15.030000  77.685000 24.540000  77.755000 ;
      RECT 15.030000 100.685000 24.540000 100.755000 ;
      RECT 15.030000 100.685000 24.540000 100.755000 ;
      RECT 15.030000 123.590000 24.540000 123.660000 ;
      RECT 15.030000 123.590000 24.540000 123.660000 ;
      RECT 15.030000 146.660000 16.525000 146.730000 ;
      RECT 15.030000 169.665000 16.525000 169.735000 ;
      RECT 15.030000 190.030000 15.340000 190.100000 ;
      RECT 15.035000 161.560000 57.955000 161.630000 ;
      RECT 15.035000 161.560000 57.955000 161.630000 ;
      RECT 15.050000  69.490000 58.005000  69.560000 ;
      RECT 15.050000  69.490000 58.005000  69.560000 ;
      RECT 15.055000 138.630000 57.870000 138.700000 ;
      RECT 15.055000 138.630000 57.870000 138.700000 ;
      RECT 15.055000 184.515000 59.010000 184.585000 ;
      RECT 15.070000 146.770000 18.190000 148.295000 ;
      RECT 15.075000  44.755000 59.710000  44.825000 ;
      RECT 15.075000  44.755000 59.710000  44.825000 ;
      RECT 15.085000  92.455000 58.100000  92.525000 ;
      RECT 15.085000  92.455000 58.100000  92.525000 ;
      RECT 15.085000 190.155000 75.000000 190.280000 ;
      RECT 15.090000 115.490000 57.975000 115.560000 ;
      RECT 15.090000 115.490000 57.975000 115.560000 ;
      RECT 15.100000  54.730000 16.525000  54.800000 ;
      RECT 15.100000  77.755000 24.540000  77.825000 ;
      RECT 15.100000  77.755000 24.540000  77.825000 ;
      RECT 15.100000 100.755000 24.540000 100.825000 ;
      RECT 15.100000 100.755000 24.540000 100.825000 ;
      RECT 15.100000 123.660000 24.540000 123.730000 ;
      RECT 15.100000 123.660000 24.540000 123.730000 ;
      RECT 15.100000 146.730000 16.525000 146.800000 ;
      RECT 15.100000 169.735000 16.525000 169.805000 ;
      RECT 15.100000 190.100000 15.340000 190.170000 ;
      RECT 15.105000 161.490000 58.025000 161.560000 ;
      RECT 15.105000 161.490000 58.025000 161.560000 ;
      RECT 15.120000  69.420000 58.075000  69.490000 ;
      RECT 15.120000  69.420000 58.075000  69.490000 ;
      RECT 15.125000 138.560000 57.940000 138.630000 ;
      RECT 15.125000 138.560000 57.940000 138.630000 ;
      RECT 15.125000 146.800000 16.525000 146.825000 ;
      RECT 15.125000 184.445000 59.080000 184.515000 ;
      RECT 15.145000  44.685000 59.780000  44.755000 ;
      RECT 15.145000  44.685000 59.780000  44.755000 ;
      RECT 15.155000  92.385000 58.170000  92.455000 ;
      RECT 15.155000  92.385000 58.170000  92.455000 ;
      RECT 15.160000 115.420000 58.045000 115.490000 ;
      RECT 15.160000 115.420000 58.045000 115.490000 ;
      RECT 15.170000  54.800000 16.525000  54.870000 ;
      RECT 15.170000  77.825000 24.540000  77.895000 ;
      RECT 15.170000  77.825000 24.540000  77.895000 ;
      RECT 15.170000 100.825000 24.540000 100.895000 ;
      RECT 15.170000 100.825000 24.540000 100.895000 ;
      RECT 15.170000 123.730000 24.540000 123.800000 ;
      RECT 15.170000 123.730000 24.540000 123.800000 ;
      RECT 15.170000 169.805000 16.525000 169.875000 ;
      RECT 15.170000 190.170000 15.340000 190.240000 ;
      RECT 15.175000 161.420000 58.095000 161.490000 ;
      RECT 15.175000 161.420000 58.095000 161.490000 ;
      RECT 15.190000  69.350000 58.145000  69.420000 ;
      RECT 15.190000  69.350000 58.145000  69.420000 ;
      RECT 15.195000 138.490000 58.010000 138.560000 ;
      RECT 15.195000 138.490000 58.010000 138.560000 ;
      RECT 15.195000 146.825000 16.525000 146.895000 ;
      RECT 15.195000 184.375000 59.150000 184.445000 ;
      RECT 15.205000  54.905000 18.790000  56.295000 ;
      RECT 15.210000 190.240000 15.340000 190.280000 ;
      RECT 15.215000  44.615000 59.850000  44.685000 ;
      RECT 15.215000  44.615000 59.850000  44.685000 ;
      RECT 15.225000  92.315000 58.240000  92.385000 ;
      RECT 15.225000  92.315000 58.240000  92.385000 ;
      RECT 15.230000 115.350000 58.115000 115.420000 ;
      RECT 15.230000 115.350000 58.115000 115.420000 ;
      RECT 15.240000  54.870000 16.525000  54.940000 ;
      RECT 15.240000  77.895000 24.540000  77.965000 ;
      RECT 15.240000  77.895000 24.540000  77.965000 ;
      RECT 15.240000 100.895000 24.540000 100.965000 ;
      RECT 15.240000 100.895000 24.540000 100.965000 ;
      RECT 15.240000 123.800000 24.540000 123.870000 ;
      RECT 15.240000 123.800000 24.540000 123.870000 ;
      RECT 15.240000 169.875000 16.525000 169.945000 ;
      RECT 15.245000 161.350000 58.165000 161.420000 ;
      RECT 15.245000 161.350000 58.165000 161.420000 ;
      RECT 15.260000  69.280000 58.215000  69.350000 ;
      RECT 15.260000  69.280000 58.215000  69.350000 ;
      RECT 15.265000 138.420000 58.080000 138.490000 ;
      RECT 15.265000 138.420000 58.080000 138.490000 ;
      RECT 15.265000 146.895000 16.595000 146.965000 ;
      RECT 15.265000 184.305000 59.220000 184.375000 ;
      RECT 15.285000  44.545000 59.920000  44.615000 ;
      RECT 15.285000  44.545000 59.920000  44.615000 ;
      RECT 15.295000  92.245000 58.310000  92.315000 ;
      RECT 15.295000  92.245000 58.310000  92.315000 ;
      RECT 15.300000 115.280000 58.185000 115.350000 ;
      RECT 15.300000 115.280000 58.185000 115.350000 ;
      RECT 15.310000  54.940000 16.525000  55.010000 ;
      RECT 15.310000  77.965000 24.540000  78.035000 ;
      RECT 15.310000  77.965000 24.540000  78.035000 ;
      RECT 15.310000 100.965000 24.540000 101.035000 ;
      RECT 15.310000 100.965000 24.540000 101.035000 ;
      RECT 15.310000 123.870000 24.540000 123.940000 ;
      RECT 15.310000 123.870000 24.540000 123.940000 ;
      RECT 15.310000 169.945000 16.525000 170.015000 ;
      RECT 15.315000 161.280000 58.235000 161.350000 ;
      RECT 15.315000 161.280000 58.235000 161.350000 ;
      RECT 15.330000  69.210000 58.285000  69.280000 ;
      RECT 15.330000  69.210000 58.285000  69.280000 ;
      RECT 15.335000 138.350000 58.150000 138.420000 ;
      RECT 15.335000 138.350000 58.150000 138.420000 ;
      RECT 15.335000 146.965000 16.665000 147.035000 ;
      RECT 15.335000 184.235000 59.290000 184.305000 ;
      RECT 15.345000  55.010000 16.525000  55.045000 ;
      RECT 15.355000  44.475000 59.990000  44.545000 ;
      RECT 15.355000  44.475000 59.990000  44.545000 ;
      RECT 15.365000  92.175000 58.380000  92.245000 ;
      RECT 15.365000  92.175000 58.380000  92.245000 ;
      RECT 15.370000 115.210000 58.255000 115.280000 ;
      RECT 15.370000 115.210000 58.255000 115.280000 ;
      RECT 15.380000  78.035000 24.540000  78.105000 ;
      RECT 15.380000  78.035000 24.540000  78.105000 ;
      RECT 15.380000 101.035000 24.540000 101.105000 ;
      RECT 15.380000 101.035000 24.540000 101.105000 ;
      RECT 15.380000 123.940000 24.540000 124.010000 ;
      RECT 15.380000 123.940000 24.540000 124.010000 ;
      RECT 15.380000 170.015000 16.525000 170.085000 ;
      RECT 15.385000 161.210000 58.305000 161.280000 ;
      RECT 15.385000 161.210000 58.305000 161.280000 ;
      RECT 15.400000  69.140000 58.355000  69.210000 ;
      RECT 15.400000  69.140000 58.355000  69.210000 ;
      RECT 15.405000 138.280000 58.220000 138.350000 ;
      RECT 15.405000 138.280000 58.220000 138.350000 ;
      RECT 15.405000 147.035000 16.735000 147.105000 ;
      RECT 15.405000 184.165000 59.360000 184.235000 ;
      RECT 15.415000  55.045000 17.345000  55.115000 ;
      RECT 15.425000  44.405000 60.060000  44.475000 ;
      RECT 15.425000  44.405000 60.060000  44.475000 ;
      RECT 15.435000  92.105000 58.450000  92.175000 ;
      RECT 15.435000  92.105000 58.450000  92.175000 ;
      RECT 15.440000 115.140000 58.325000 115.210000 ;
      RECT 15.440000 115.140000 58.325000 115.210000 ;
      RECT 15.450000  78.105000 24.540000  78.175000 ;
      RECT 15.450000  78.105000 24.540000  78.175000 ;
      RECT 15.450000 101.105000 24.540000 101.175000 ;
      RECT 15.450000 101.105000 24.540000 101.175000 ;
      RECT 15.450000 124.010000 24.540000 124.080000 ;
      RECT 15.450000 124.010000 24.540000 124.080000 ;
      RECT 15.450000 170.085000 16.525000 170.155000 ;
      RECT 15.455000 161.140000 58.375000 161.210000 ;
      RECT 15.455000 161.140000 58.375000 161.210000 ;
      RECT 15.470000  69.070000 58.425000  69.140000 ;
      RECT 15.470000  69.070000 58.425000  69.140000 ;
      RECT 15.475000 138.210000 58.290000 138.280000 ;
      RECT 15.475000 138.210000 58.290000 138.280000 ;
      RECT 15.475000 147.105000 16.805000 147.175000 ;
      RECT 15.475000 184.095000 59.430000 184.165000 ;
      RECT 15.485000  29.430000 59.190000  29.500000 ;
      RECT 15.485000  29.430000 59.190000  29.500000 ;
      RECT 15.485000  29.430000 60.970000  31.015000 ;
      RECT 15.485000  29.500000 59.260000  29.570000 ;
      RECT 15.485000  29.500000 59.260000  29.570000 ;
      RECT 15.485000  29.570000 59.330000  29.640000 ;
      RECT 15.485000  29.570000 59.330000  29.640000 ;
      RECT 15.485000  29.640000 59.400000  29.710000 ;
      RECT 15.485000  29.640000 59.400000  29.710000 ;
      RECT 15.485000  29.710000 59.470000  29.780000 ;
      RECT 15.485000  29.710000 59.470000  29.780000 ;
      RECT 15.485000  29.780000 59.540000  29.850000 ;
      RECT 15.485000  29.780000 59.540000  29.850000 ;
      RECT 15.485000  29.850000 59.610000  29.920000 ;
      RECT 15.485000  29.850000 59.610000  29.920000 ;
      RECT 15.485000  29.920000 59.680000  29.990000 ;
      RECT 15.485000  29.920000 59.680000  29.990000 ;
      RECT 15.485000  29.990000 59.750000  30.060000 ;
      RECT 15.485000  29.990000 59.750000  30.060000 ;
      RECT 15.485000  30.060000 59.820000  30.130000 ;
      RECT 15.485000  30.060000 59.820000  30.130000 ;
      RECT 15.485000  30.130000 59.890000  30.200000 ;
      RECT 15.485000  30.130000 59.890000  30.200000 ;
      RECT 15.485000  30.200000 59.960000  30.270000 ;
      RECT 15.485000  30.200000 59.960000  30.270000 ;
      RECT 15.485000  30.270000 60.030000  30.340000 ;
      RECT 15.485000  30.270000 60.030000  30.340000 ;
      RECT 15.485000  30.340000 60.100000  30.410000 ;
      RECT 15.485000  30.340000 60.100000  30.410000 ;
      RECT 15.485000  30.410000 60.170000  30.480000 ;
      RECT 15.485000  30.410000 60.170000  30.480000 ;
      RECT 15.485000  30.480000 60.240000  30.550000 ;
      RECT 15.485000  30.480000 60.240000  30.550000 ;
      RECT 15.485000  30.550000 60.310000  30.620000 ;
      RECT 15.485000  30.550000 60.310000  30.620000 ;
      RECT 15.485000  30.620000 60.380000  30.690000 ;
      RECT 15.485000  30.620000 60.380000  30.690000 ;
      RECT 15.485000  30.690000 60.450000  30.760000 ;
      RECT 15.485000  30.690000 60.450000  30.760000 ;
      RECT 15.485000  30.760000 60.520000  30.830000 ;
      RECT 15.485000  30.760000 60.520000  30.830000 ;
      RECT 15.485000  30.830000 60.590000  30.900000 ;
      RECT 15.485000  30.830000 60.590000  30.900000 ;
      RECT 15.485000  30.900000 60.660000  30.970000 ;
      RECT 15.485000  30.900000 60.660000  30.970000 ;
      RECT 15.485000  30.970000 60.730000  31.040000 ;
      RECT 15.485000  30.970000 60.730000  31.040000 ;
      RECT 15.485000  31.015000 60.970000  35.550000 ;
      RECT 15.485000  31.040000 60.800000  31.070000 ;
      RECT 15.485000  31.040000 60.800000  31.070000 ;
      RECT 15.485000  31.070000 60.830000  35.550000 ;
      RECT 15.485000  35.550000 60.970000  35.975000 ;
      RECT 15.485000  55.115000 17.415000  55.185000 ;
      RECT 15.495000  44.335000 60.130000  44.405000 ;
      RECT 15.495000  44.335000 60.130000  44.405000 ;
      RECT 15.505000  29.410000 59.170000  29.430000 ;
      RECT 15.505000  29.410000 59.170000  29.430000 ;
      RECT 15.505000  92.035000 58.520000  92.105000 ;
      RECT 15.505000  92.035000 58.520000  92.105000 ;
      RECT 15.510000 115.070000 58.395000 115.140000 ;
      RECT 15.510000 115.070000 58.395000 115.140000 ;
      RECT 15.520000  78.175000 24.540000  78.245000 ;
      RECT 15.520000  78.175000 24.540000  78.245000 ;
      RECT 15.520000 101.175000 24.540000 101.245000 ;
      RECT 15.520000 101.175000 24.540000 101.245000 ;
      RECT 15.520000 124.080000 24.540000 124.150000 ;
      RECT 15.520000 124.080000 24.540000 124.150000 ;
      RECT 15.520000 170.155000 16.525000 170.225000 ;
      RECT 15.525000 161.070000 58.445000 161.140000 ;
      RECT 15.525000 161.070000 58.445000 161.140000 ;
      RECT 15.540000  69.000000 58.495000  69.070000 ;
      RECT 15.540000  69.000000 58.495000  69.070000 ;
      RECT 15.545000 138.140000 58.360000 138.210000 ;
      RECT 15.545000 138.140000 58.360000 138.210000 ;
      RECT 15.545000 147.175000 16.875000 147.245000 ;
      RECT 15.545000 184.025000 59.500000 184.095000 ;
      RECT 15.555000  35.550000 60.830000  35.620000 ;
      RECT 15.555000  35.550000 60.830000  35.620000 ;
      RECT 15.555000  55.185000 17.485000  55.255000 ;
      RECT 15.565000  44.265000 60.200000  44.335000 ;
      RECT 15.565000  44.265000 60.200000  44.335000 ;
      RECT 15.575000  29.340000 59.100000  29.410000 ;
      RECT 15.575000  29.340000 59.100000  29.410000 ;
      RECT 15.575000  91.965000 58.590000  92.035000 ;
      RECT 15.575000  91.965000 58.590000  92.035000 ;
      RECT 15.580000 115.000000 58.465000 115.070000 ;
      RECT 15.580000 115.000000 58.465000 115.070000 ;
      RECT 15.590000  78.245000 24.540000  78.315000 ;
      RECT 15.590000  78.245000 24.540000  78.315000 ;
      RECT 15.590000 101.245000 24.540000 101.315000 ;
      RECT 15.590000 101.245000 24.540000 101.315000 ;
      RECT 15.590000 124.150000 24.540000 124.220000 ;
      RECT 15.590000 124.150000 24.540000 124.220000 ;
      RECT 15.590000 170.225000 16.525000 170.295000 ;
      RECT 15.595000 161.000000 58.515000 161.070000 ;
      RECT 15.595000 161.000000 58.515000 161.070000 ;
      RECT 15.610000  68.930000 58.565000  69.000000 ;
      RECT 15.610000  68.930000 58.565000  69.000000 ;
      RECT 15.615000 138.070000 58.430000 138.140000 ;
      RECT 15.615000 138.070000 58.430000 138.140000 ;
      RECT 15.615000 147.245000 16.945000 147.315000 ;
      RECT 15.615000 183.955000 59.570000 184.025000 ;
      RECT 15.625000  35.620000 60.830000  35.690000 ;
      RECT 15.625000  35.620000 60.830000  35.690000 ;
      RECT 15.625000  55.255000 17.555000  55.325000 ;
      RECT 15.635000  44.195000 60.270000  44.265000 ;
      RECT 15.635000  44.195000 60.270000  44.265000 ;
      RECT 15.645000  29.270000 59.030000  29.340000 ;
      RECT 15.645000  29.270000 59.030000  29.340000 ;
      RECT 15.645000  91.895000 58.660000  91.965000 ;
      RECT 15.645000  91.895000 58.660000  91.965000 ;
      RECT 15.650000 114.930000 58.535000 115.000000 ;
      RECT 15.650000 114.930000 58.535000 115.000000 ;
      RECT 15.660000  78.315000 24.540000  78.385000 ;
      RECT 15.660000  78.315000 24.540000  78.385000 ;
      RECT 15.660000 101.315000 24.540000 101.385000 ;
      RECT 15.660000 101.315000 24.540000 101.385000 ;
      RECT 15.660000 124.220000 24.540000 124.290000 ;
      RECT 15.660000 124.220000 24.540000 124.290000 ;
      RECT 15.660000 170.295000 16.525000 170.365000 ;
      RECT 15.665000 160.930000 58.585000 161.000000 ;
      RECT 15.665000 160.930000 58.585000 161.000000 ;
      RECT 15.680000  68.860000 58.635000  68.930000 ;
      RECT 15.680000  68.860000 58.635000  68.930000 ;
      RECT 15.685000 138.000000 58.500000 138.070000 ;
      RECT 15.685000 138.000000 58.500000 138.070000 ;
      RECT 15.685000 147.315000 17.015000 147.385000 ;
      RECT 15.685000 183.885000 59.640000 183.955000 ;
      RECT 15.695000  35.690000 60.830000  35.760000 ;
      RECT 15.695000  35.690000 60.830000  35.760000 ;
      RECT 15.695000  55.325000 17.625000  55.395000 ;
      RECT 15.705000  44.125000 60.340000  44.195000 ;
      RECT 15.705000  44.125000 60.340000  44.195000 ;
      RECT 15.715000  29.200000 58.960000  29.270000 ;
      RECT 15.715000  29.200000 58.960000  29.270000 ;
      RECT 15.715000  91.825000 58.730000  91.895000 ;
      RECT 15.715000  91.825000 58.730000  91.895000 ;
      RECT 15.720000 114.860000 58.605000 114.930000 ;
      RECT 15.720000 114.860000 58.605000 114.930000 ;
      RECT 15.730000  78.385000 24.540000  78.455000 ;
      RECT 15.730000  78.385000 24.540000  78.455000 ;
      RECT 15.730000 101.385000 24.540000 101.455000 ;
      RECT 15.730000 101.385000 24.540000 101.455000 ;
      RECT 15.730000 124.290000 24.540000 124.360000 ;
      RECT 15.730000 124.290000 24.540000 124.360000 ;
      RECT 15.730000 170.365000 16.525000 170.435000 ;
      RECT 15.735000 160.860000 58.655000 160.930000 ;
      RECT 15.735000 160.860000 58.655000 160.930000 ;
      RECT 15.750000  68.790000 58.705000  68.860000 ;
      RECT 15.750000  68.790000 58.705000  68.860000 ;
      RECT 15.755000 137.930000 58.570000 138.000000 ;
      RECT 15.755000 137.930000 58.570000 138.000000 ;
      RECT 15.755000 147.385000 17.085000 147.455000 ;
      RECT 15.755000 183.815000 59.710000 183.885000 ;
      RECT 15.765000  35.760000 60.830000  35.830000 ;
      RECT 15.765000  35.760000 60.830000  35.830000 ;
      RECT 15.765000  55.395000 17.695000  55.465000 ;
      RECT 15.770000  35.830000 60.830000  35.835000 ;
      RECT 15.770000  35.830000 60.830000  35.835000 ;
      RECT 15.775000  44.055000 60.410000  44.125000 ;
      RECT 15.775000  44.055000 60.410000  44.125000 ;
      RECT 15.785000  29.130000 58.890000  29.200000 ;
      RECT 15.785000  29.130000 58.890000  29.200000 ;
      RECT 15.785000  91.755000 58.800000  91.825000 ;
      RECT 15.785000  91.755000 58.800000  91.825000 ;
      RECT 15.790000 114.790000 58.675000 114.860000 ;
      RECT 15.790000 114.790000 58.675000 114.860000 ;
      RECT 15.800000  78.455000 24.540000  78.525000 ;
      RECT 15.800000  78.455000 24.540000  78.525000 ;
      RECT 15.800000 101.455000 24.540000 101.525000 ;
      RECT 15.800000 101.455000 24.540000 101.525000 ;
      RECT 15.800000 124.360000 24.540000 124.430000 ;
      RECT 15.800000 124.360000 24.540000 124.430000 ;
      RECT 15.800000 170.435000 16.525000 170.505000 ;
      RECT 15.805000 160.790000 58.725000 160.860000 ;
      RECT 15.805000 160.790000 58.725000 160.860000 ;
      RECT 15.820000  68.720000 58.775000  68.790000 ;
      RECT 15.820000  68.720000 58.775000  68.790000 ;
      RECT 15.825000 137.860000 58.640000 137.930000 ;
      RECT 15.825000 137.860000 58.640000 137.930000 ;
      RECT 15.825000 147.455000 17.155000 147.525000 ;
      RECT 15.825000 183.745000 59.780000 183.815000 ;
      RECT 15.835000  55.465000 17.765000  55.535000 ;
      RECT 15.840000  35.835000 54.390000  35.905000 ;
      RECT 15.840000  35.835000 54.390000  35.905000 ;
      RECT 15.845000  43.985000 60.480000  44.055000 ;
      RECT 15.845000  43.985000 60.480000  44.055000 ;
      RECT 15.855000  29.060000 58.820000  29.130000 ;
      RECT 15.855000  29.060000 58.820000  29.130000 ;
      RECT 15.855000  91.685000 58.870000  91.755000 ;
      RECT 15.855000  91.685000 58.870000  91.755000 ;
      RECT 15.860000 114.720000 58.745000 114.790000 ;
      RECT 15.860000 114.720000 58.745000 114.790000 ;
      RECT 15.870000  78.525000 24.540000  78.595000 ;
      RECT 15.870000  78.525000 24.540000  78.595000 ;
      RECT 15.870000 101.525000 24.540000 101.595000 ;
      RECT 15.870000 101.525000 24.540000 101.595000 ;
      RECT 15.870000 124.430000 24.540000 124.500000 ;
      RECT 15.870000 124.430000 24.540000 124.500000 ;
      RECT 15.870000 170.505000 16.525000 170.575000 ;
      RECT 15.875000 160.720000 58.795000 160.790000 ;
      RECT 15.875000 160.720000 58.795000 160.790000 ;
      RECT 15.890000  68.650000 58.845000  68.720000 ;
      RECT 15.890000  68.650000 58.845000  68.720000 ;
      RECT 15.895000 137.790000 58.710000 137.860000 ;
      RECT 15.895000 137.790000 58.710000 137.860000 ;
      RECT 15.895000 147.525000 17.225000 147.595000 ;
      RECT 15.895000 183.675000 59.850000 183.745000 ;
      RECT 15.905000  55.535000 17.835000  55.605000 ;
      RECT 15.910000  35.905000 54.390000  35.975000 ;
      RECT 15.910000  35.905000 54.390000  35.975000 ;
      RECT 15.910000  35.975000 54.530000  38.195000 ;
      RECT 15.915000  43.915000 60.550000  43.985000 ;
      RECT 15.915000  43.915000 60.550000  43.985000 ;
      RECT 15.925000  28.990000 58.750000  29.060000 ;
      RECT 15.925000  28.990000 58.750000  29.060000 ;
      RECT 15.925000  91.615000 58.940000  91.685000 ;
      RECT 15.925000  91.615000 58.940000  91.685000 ;
      RECT 15.930000 114.650000 58.815000 114.720000 ;
      RECT 15.930000 114.650000 58.815000 114.720000 ;
      RECT 15.940000  78.595000 24.540000  78.665000 ;
      RECT 15.940000  78.595000 24.540000  78.665000 ;
      RECT 15.940000 101.595000 24.540000 101.665000 ;
      RECT 15.940000 101.595000 24.540000 101.665000 ;
      RECT 15.940000 124.500000 24.540000 124.570000 ;
      RECT 15.940000 124.500000 24.540000 124.570000 ;
      RECT 15.940000 170.575000 16.525000 170.645000 ;
      RECT 15.945000 160.650000 58.865000 160.720000 ;
      RECT 15.945000 160.650000 58.865000 160.720000 ;
      RECT 15.960000  68.580000 58.915000  68.650000 ;
      RECT 15.960000  68.580000 58.915000  68.650000 ;
      RECT 15.965000 137.720000 58.780000 137.790000 ;
      RECT 15.965000 137.720000 58.780000 137.790000 ;
      RECT 15.965000 147.595000 17.295000 147.665000 ;
      RECT 15.965000 183.605000 59.920000 183.675000 ;
      RECT 15.975000  55.605000 17.905000  55.675000 ;
      RECT 15.980000  35.975000 54.390000  36.045000 ;
      RECT 15.980000  35.975000 54.390000  36.045000 ;
      RECT 15.985000  43.845000 60.620000  43.915000 ;
      RECT 15.985000  43.845000 60.620000  43.915000 ;
      RECT 15.995000  28.920000 58.680000  28.990000 ;
      RECT 15.995000  28.920000 58.680000  28.990000 ;
      RECT 15.995000  91.545000 59.010000  91.615000 ;
      RECT 15.995000  91.545000 59.010000  91.615000 ;
      RECT 16.000000 114.580000 58.885000 114.650000 ;
      RECT 16.000000 114.580000 58.885000 114.650000 ;
      RECT 16.010000  78.665000 24.540000  78.735000 ;
      RECT 16.010000  78.665000 24.540000  78.735000 ;
      RECT 16.010000 101.665000 24.540000 101.735000 ;
      RECT 16.010000 101.665000 24.540000 101.735000 ;
      RECT 16.010000 124.570000 24.540000 124.640000 ;
      RECT 16.010000 124.570000 24.540000 124.640000 ;
      RECT 16.010000 170.645000 16.525000 170.715000 ;
      RECT 16.015000 160.580000 58.935000 160.650000 ;
      RECT 16.015000 160.580000 58.935000 160.650000 ;
      RECT 16.030000  68.510000 58.985000  68.580000 ;
      RECT 16.030000  68.510000 58.985000  68.580000 ;
      RECT 16.035000 137.650000 58.850000 137.720000 ;
      RECT 16.035000 137.650000 58.850000 137.720000 ;
      RECT 16.035000 147.665000 17.365000 147.735000 ;
      RECT 16.035000 183.535000 59.990000 183.605000 ;
      RECT 16.045000  55.675000 17.975000  55.745000 ;
      RECT 16.050000  36.045000 54.390000  36.115000 ;
      RECT 16.050000  36.045000 54.390000  36.115000 ;
      RECT 16.055000  43.775000 60.690000  43.845000 ;
      RECT 16.055000  43.775000 60.690000  43.845000 ;
      RECT 16.065000  28.850000 58.610000  28.920000 ;
      RECT 16.065000  28.850000 58.610000  28.920000 ;
      RECT 16.065000  91.475000 59.080000  91.545000 ;
      RECT 16.065000  91.475000 59.080000  91.545000 ;
      RECT 16.070000  43.760000 59.300000  45.430000 ;
      RECT 16.070000 114.510000 58.955000 114.580000 ;
      RECT 16.070000 114.510000 58.955000 114.580000 ;
      RECT 16.080000  78.735000 24.540000  78.805000 ;
      RECT 16.080000  78.735000 24.540000  78.805000 ;
      RECT 16.080000 101.735000 24.540000 101.805000 ;
      RECT 16.080000 101.735000 24.540000 101.805000 ;
      RECT 16.080000 124.640000 24.540000 124.710000 ;
      RECT 16.080000 124.640000 24.540000 124.710000 ;
      RECT 16.080000 170.715000 16.525000 170.785000 ;
      RECT 16.085000 160.510000 59.005000 160.580000 ;
      RECT 16.085000 160.510000 59.005000 160.580000 ;
      RECT 16.100000  68.440000 59.055000  68.510000 ;
      RECT 16.100000  68.440000 59.055000  68.510000 ;
      RECT 16.105000 137.580000 58.920000 137.650000 ;
      RECT 16.105000 137.580000 58.920000 137.650000 ;
      RECT 16.105000 147.735000 17.435000 147.805000 ;
      RECT 16.105000 183.465000 60.060000 183.535000 ;
      RECT 16.115000  55.745000 18.045000  55.815000 ;
      RECT 16.120000  36.115000 54.390000  36.185000 ;
      RECT 16.120000  36.115000 54.390000  36.185000 ;
      RECT 16.125000  43.705000 60.760000  43.775000 ;
      RECT 16.125000  43.705000 60.760000  43.775000 ;
      RECT 16.135000  28.780000 58.540000  28.850000 ;
      RECT 16.135000  28.780000 58.540000  28.850000 ;
      RECT 16.135000  91.405000 59.150000  91.475000 ;
      RECT 16.135000  91.405000 59.150000  91.475000 ;
      RECT 16.140000 114.440000 59.025000 114.510000 ;
      RECT 16.140000 114.440000 59.025000 114.510000 ;
      RECT 16.150000  78.805000 24.540000  78.875000 ;
      RECT 16.150000  78.805000 24.540000  78.875000 ;
      RECT 16.150000 101.805000 24.540000 101.875000 ;
      RECT 16.150000 101.805000 24.540000 101.875000 ;
      RECT 16.150000 124.710000 24.540000 124.780000 ;
      RECT 16.150000 124.710000 24.540000 124.780000 ;
      RECT 16.150000 170.785000 16.525000 170.855000 ;
      RECT 16.155000 160.440000 59.075000 160.510000 ;
      RECT 16.155000 160.440000 59.075000 160.510000 ;
      RECT 16.170000  68.370000 59.125000  68.440000 ;
      RECT 16.170000  68.370000 59.125000  68.440000 ;
      RECT 16.175000 137.510000 58.990000 137.580000 ;
      RECT 16.175000 137.510000 58.990000 137.580000 ;
      RECT 16.175000 147.805000 17.505000 147.875000 ;
      RECT 16.175000 183.395000 60.130000 183.465000 ;
      RECT 16.185000  55.815000 18.115000  55.885000 ;
      RECT 16.190000  36.185000 54.390000  36.255000 ;
      RECT 16.190000  36.185000 54.390000  36.255000 ;
      RECT 16.190000  43.640000 60.830000  43.705000 ;
      RECT 16.190000  43.640000 60.830000  43.705000 ;
      RECT 16.205000  28.710000 58.470000  28.780000 ;
      RECT 16.205000  28.710000 58.470000  28.780000 ;
      RECT 16.205000  91.335000 59.220000  91.405000 ;
      RECT 16.205000  91.335000 59.220000  91.405000 ;
      RECT 16.210000 114.370000 59.095000 114.440000 ;
      RECT 16.210000 114.370000 59.095000 114.440000 ;
      RECT 16.220000  78.875000 24.540000  78.945000 ;
      RECT 16.220000  78.875000 24.540000  78.945000 ;
      RECT 16.220000 101.875000 24.540000 101.945000 ;
      RECT 16.220000 101.875000 24.540000 101.945000 ;
      RECT 16.220000 124.780000 24.540000 124.850000 ;
      RECT 16.220000 124.780000 24.540000 124.850000 ;
      RECT 16.220000 170.855000 16.525000 170.925000 ;
      RECT 16.225000 160.370000 59.145000 160.440000 ;
      RECT 16.225000 160.370000 59.145000 160.440000 ;
      RECT 16.240000  68.300000 59.195000  68.370000 ;
      RECT 16.240000  68.300000 59.195000  68.370000 ;
      RECT 16.245000 137.440000 59.060000 137.510000 ;
      RECT 16.245000 137.440000 59.060000 137.510000 ;
      RECT 16.245000 147.875000 17.575000 147.945000 ;
      RECT 16.245000 183.325000 60.200000 183.395000 ;
      RECT 16.255000  55.885000 18.185000  55.955000 ;
      RECT 16.260000  36.255000 54.390000  36.325000 ;
      RECT 16.260000  36.255000 54.390000  36.325000 ;
      RECT 16.260000  43.570000 60.830000  43.640000 ;
      RECT 16.260000  43.570000 60.830000  43.640000 ;
      RECT 16.275000  28.640000 58.400000  28.710000 ;
      RECT 16.275000  28.640000 58.400000  28.710000 ;
      RECT 16.275000  91.265000 59.290000  91.335000 ;
      RECT 16.275000  91.265000 59.290000  91.335000 ;
      RECT 16.280000 114.300000 59.165000 114.370000 ;
      RECT 16.280000 114.300000 59.165000 114.370000 ;
      RECT 16.290000  78.945000 24.540000  79.015000 ;
      RECT 16.290000  78.945000 24.540000  79.015000 ;
      RECT 16.290000 101.945000 24.540000 102.015000 ;
      RECT 16.290000 101.945000 24.540000 102.015000 ;
      RECT 16.290000 124.850000 24.540000 124.920000 ;
      RECT 16.290000 124.850000 24.540000 124.920000 ;
      RECT 16.290000 170.925000 16.525000 170.995000 ;
      RECT 16.295000 160.300000 59.215000 160.370000 ;
      RECT 16.295000 160.300000 59.215000 160.370000 ;
      RECT 16.310000  68.230000 59.265000  68.300000 ;
      RECT 16.310000  68.230000 59.265000  68.300000 ;
      RECT 16.315000 137.370000 59.130000 137.440000 ;
      RECT 16.315000 137.370000 59.130000 137.440000 ;
      RECT 16.315000 147.945000 17.645000 148.015000 ;
      RECT 16.315000 183.255000 60.270000 183.325000 ;
      RECT 16.325000  55.955000 18.255000  56.025000 ;
      RECT 16.330000  36.325000 54.390000  36.395000 ;
      RECT 16.330000  36.325000 54.390000  36.395000 ;
      RECT 16.330000  43.500000 60.830000  43.570000 ;
      RECT 16.330000  43.500000 60.830000  43.570000 ;
      RECT 16.345000  28.570000 58.330000  28.640000 ;
      RECT 16.345000  28.570000 58.330000  28.640000 ;
      RECT 16.345000  91.195000 59.360000  91.265000 ;
      RECT 16.345000  91.195000 59.360000  91.265000 ;
      RECT 16.350000 114.230000 59.235000 114.300000 ;
      RECT 16.350000 114.230000 59.235000 114.300000 ;
      RECT 16.360000  79.015000 24.540000  79.085000 ;
      RECT 16.360000  79.015000 24.540000  79.085000 ;
      RECT 16.360000 102.015000 24.540000 102.085000 ;
      RECT 16.360000 102.015000 24.540000 102.085000 ;
      RECT 16.360000 124.920000 24.540000 124.990000 ;
      RECT 16.360000 124.920000 24.540000 124.990000 ;
      RECT 16.360000 170.995000 16.525000 171.065000 ;
      RECT 16.365000 160.230000 59.285000 160.300000 ;
      RECT 16.365000 160.230000 59.285000 160.300000 ;
      RECT 16.380000  68.160000 59.335000  68.230000 ;
      RECT 16.380000  68.160000 59.335000  68.230000 ;
      RECT 16.385000 137.300000 59.200000 137.370000 ;
      RECT 16.385000 137.300000 59.200000 137.370000 ;
      RECT 16.385000 148.015000 17.715000 148.085000 ;
      RECT 16.385000 183.185000 60.340000 183.255000 ;
      RECT 16.395000  56.025000 18.325000  56.095000 ;
      RECT 16.400000  36.395000 54.390000  36.465000 ;
      RECT 16.400000  36.395000 54.390000  36.465000 ;
      RECT 16.400000  43.430000 60.830000  43.500000 ;
      RECT 16.400000  43.430000 60.830000  43.500000 ;
      RECT 16.415000  28.500000 58.260000  28.570000 ;
      RECT 16.415000  28.500000 58.260000  28.570000 ;
      RECT 16.415000  91.125000 59.430000  91.195000 ;
      RECT 16.415000  91.125000 59.430000  91.195000 ;
      RECT 16.420000 114.160000 59.305000 114.230000 ;
      RECT 16.420000 114.160000 59.305000 114.230000 ;
      RECT 16.430000  79.085000 24.540000  79.155000 ;
      RECT 16.430000  79.085000 24.540000  79.155000 ;
      RECT 16.430000 102.085000 24.540000 102.155000 ;
      RECT 16.430000 102.085000 24.540000 102.155000 ;
      RECT 16.430000 124.990000 24.540000 125.060000 ;
      RECT 16.430000 124.990000 24.540000 125.060000 ;
      RECT 16.430000 171.065000 16.525000 171.135000 ;
      RECT 16.435000 160.160000 59.355000 160.230000 ;
      RECT 16.435000 160.160000 59.355000 160.230000 ;
      RECT 16.450000  68.090000 59.405000  68.160000 ;
      RECT 16.450000  68.090000 59.405000  68.160000 ;
      RECT 16.455000 137.230000 59.270000 137.300000 ;
      RECT 16.455000 137.230000 59.270000 137.300000 ;
      RECT 16.455000 148.085000 17.785000 148.155000 ;
      RECT 16.455000 183.115000 60.410000 183.185000 ;
      RECT 16.465000  56.095000 18.395000  56.165000 ;
      RECT 16.470000  36.465000 54.390000  36.535000 ;
      RECT 16.470000  36.465000 54.390000  36.535000 ;
      RECT 16.470000  43.360000 60.830000  43.430000 ;
      RECT 16.470000  43.360000 60.830000  43.430000 ;
      RECT 16.485000  28.430000 58.190000  28.500000 ;
      RECT 16.485000  28.430000 58.190000  28.500000 ;
      RECT 16.485000  91.055000 59.500000  91.125000 ;
      RECT 16.485000  91.055000 59.500000  91.125000 ;
      RECT 16.490000 114.090000 59.375000 114.160000 ;
      RECT 16.490000 114.090000 59.375000 114.160000 ;
      RECT 16.500000  79.155000 24.540000  79.225000 ;
      RECT 16.500000  79.155000 24.540000  79.225000 ;
      RECT 16.500000 102.155000 24.540000 102.225000 ;
      RECT 16.500000 102.155000 24.540000 102.225000 ;
      RECT 16.500000 125.060000 24.540000 125.130000 ;
      RECT 16.500000 125.060000 24.540000 125.130000 ;
      RECT 16.500000 171.135000 16.525000 171.205000 ;
      RECT 16.505000 160.090000 59.425000 160.160000 ;
      RECT 16.505000 160.090000 59.425000 160.160000 ;
      RECT 16.520000  68.020000 59.475000  68.090000 ;
      RECT 16.520000  68.020000 59.475000  68.090000 ;
      RECT 16.525000 137.160000 59.340000 137.230000 ;
      RECT 16.525000 137.160000 59.340000 137.230000 ;
      RECT 16.525000 148.155000 17.855000 148.225000 ;
      RECT 16.525000 183.045000 60.480000 183.115000 ;
      RECT 16.535000  56.165000 18.465000  56.235000 ;
      RECT 16.540000  36.535000 54.390000  36.605000 ;
      RECT 16.540000  36.535000 54.390000  36.605000 ;
      RECT 16.540000  43.290000 60.830000  43.360000 ;
      RECT 16.540000  43.290000 60.830000  43.360000 ;
      RECT 16.555000  28.360000 58.120000  28.430000 ;
      RECT 16.555000  28.360000 58.120000  28.430000 ;
      RECT 16.555000  90.985000 59.570000  91.055000 ;
      RECT 16.555000  90.985000 59.570000  91.055000 ;
      RECT 16.560000 114.020000 59.445000 114.090000 ;
      RECT 16.560000 114.020000 59.445000 114.090000 ;
      RECT 16.570000  79.225000 24.540000  79.295000 ;
      RECT 16.570000  79.225000 24.540000  79.295000 ;
      RECT 16.570000  79.295000 58.700000  80.500000 ;
      RECT 16.570000 102.225000 24.540000 102.295000 ;
      RECT 16.570000 102.225000 24.540000 102.295000 ;
      RECT 16.570000 102.295000 58.700000 103.500000 ;
      RECT 16.570000 125.130000 24.540000 125.200000 ;
      RECT 16.570000 125.130000 24.540000 125.200000 ;
      RECT 16.575000 160.020000 59.495000 160.090000 ;
      RECT 16.575000 160.020000 59.495000 160.090000 ;
      RECT 16.590000  67.950000 59.545000  68.020000 ;
      RECT 16.590000  67.950000 59.545000  68.020000 ;
      RECT 16.590000 171.295000 58.710000 172.500000 ;
      RECT 16.595000  56.295000 58.670000  57.500000 ;
      RECT 16.595000 137.090000 59.410000 137.160000 ;
      RECT 16.595000 137.090000 59.410000 137.160000 ;
      RECT 16.595000 148.225000 17.925000 148.295000 ;
      RECT 16.595000 148.295000 58.630000 149.500000 ;
      RECT 16.595000 182.975000 60.550000 183.045000 ;
      RECT 16.605000  56.235000 18.535000  56.305000 ;
      RECT 16.610000  36.605000 54.390000  36.675000 ;
      RECT 16.610000  36.605000 54.390000  36.675000 ;
      RECT 16.610000  43.220000 60.830000  43.290000 ;
      RECT 16.610000  43.220000 60.830000  43.290000 ;
      RECT 16.625000  28.290000 58.050000  28.360000 ;
      RECT 16.625000  28.290000 58.050000  28.360000 ;
      RECT 16.625000  90.915000 59.640000  90.985000 ;
      RECT 16.625000  90.915000 59.640000  90.985000 ;
      RECT 16.630000 113.950000 59.515000 114.020000 ;
      RECT 16.630000 113.950000 59.515000 114.020000 ;
      RECT 16.640000  79.295000 24.540000  79.365000 ;
      RECT 16.640000  79.295000 24.540000  79.365000 ;
      RECT 16.640000 102.295000 24.540000 102.365000 ;
      RECT 16.640000 102.295000 24.540000 102.365000 ;
      RECT 16.640000 125.200000 24.540000 125.270000 ;
      RECT 16.640000 125.200000 24.540000 125.270000 ;
      RECT 16.645000 159.950000 59.565000 160.020000 ;
      RECT 16.645000 159.950000 59.565000 160.020000 ;
      RECT 16.660000  67.880000 59.615000  67.950000 ;
      RECT 16.660000  67.880000 59.615000  67.950000 ;
      RECT 16.665000 125.295000 58.700000 126.500000 ;
      RECT 16.665000 137.020000 59.480000 137.090000 ;
      RECT 16.665000 137.020000 59.480000 137.090000 ;
      RECT 16.665000 148.295000 17.995000 148.365000 ;
      RECT 16.665000 182.905000 60.620000 182.975000 ;
      RECT 16.675000  56.305000 18.605000  56.375000 ;
      RECT 16.680000  36.675000 54.390000  36.745000 ;
      RECT 16.680000  36.675000 54.390000  36.745000 ;
      RECT 16.680000  43.150000 60.830000  43.220000 ;
      RECT 16.680000  43.150000 60.830000  43.220000 ;
      RECT 16.695000  28.220000 57.980000  28.290000 ;
      RECT 16.695000  28.220000 57.980000  28.290000 ;
      RECT 16.695000  90.845000 59.710000  90.915000 ;
      RECT 16.695000  90.845000 59.710000  90.915000 ;
      RECT 16.700000 113.880000 59.585000 113.950000 ;
      RECT 16.700000 113.880000 59.585000 113.950000 ;
      RECT 16.710000  79.365000 24.540000  79.435000 ;
      RECT 16.710000  79.365000 24.540000  79.435000 ;
      RECT 16.710000 102.365000 24.540000 102.435000 ;
      RECT 16.710000 102.365000 24.540000 102.435000 ;
      RECT 16.710000 125.270000 24.540000 125.340000 ;
      RECT 16.710000 125.270000 24.540000 125.340000 ;
      RECT 16.715000 159.880000 59.635000 159.950000 ;
      RECT 16.715000 159.880000 59.635000 159.950000 ;
      RECT 16.730000  67.810000 59.685000  67.880000 ;
      RECT 16.730000  67.810000 59.685000  67.880000 ;
      RECT 16.735000  56.375000 18.675000  56.435000 ;
      RECT 16.735000 136.950000 59.550000 137.020000 ;
      RECT 16.735000 136.950000 59.550000 137.020000 ;
      RECT 16.735000 148.365000 18.065000 148.435000 ;
      RECT 16.735000 182.835000 60.690000 182.905000 ;
      RECT 16.750000  36.745000 54.390000  36.815000 ;
      RECT 16.750000  36.745000 54.390000  36.815000 ;
      RECT 16.750000  43.080000 60.830000  43.150000 ;
      RECT 16.750000  43.080000 60.830000  43.150000 ;
      RECT 16.750000 182.820000 58.635000 185.155000 ;
      RECT 16.765000  28.150000 57.910000  28.220000 ;
      RECT 16.765000  28.150000 57.910000  28.220000 ;
      RECT 16.765000  90.775000 59.780000  90.845000 ;
      RECT 16.765000  90.775000 59.780000  90.845000 ;
      RECT 16.770000 113.810000 59.655000 113.880000 ;
      RECT 16.770000 113.810000 59.655000 113.880000 ;
      RECT 16.780000  79.435000 24.540000  79.505000 ;
      RECT 16.780000  79.435000 24.540000  79.505000 ;
      RECT 16.780000  79.435000 57.440000  79.505000 ;
      RECT 16.780000 102.435000 24.540000 102.505000 ;
      RECT 16.780000 102.435000 24.540000 102.505000 ;
      RECT 16.780000 102.435000 57.440000 102.505000 ;
      RECT 16.780000 125.340000 24.540000 125.410000 ;
      RECT 16.780000 125.340000 24.540000 125.410000 ;
      RECT 16.785000 159.810000 59.705000 159.880000 ;
      RECT 16.785000 159.810000 59.705000 159.880000 ;
      RECT 16.800000  67.740000 59.755000  67.810000 ;
      RECT 16.800000  67.740000 59.755000  67.810000 ;
      RECT 16.800000 171.435000 57.450000 171.505000 ;
      RECT 16.805000  56.435000 57.410000  56.505000 ;
      RECT 16.805000 125.410000 24.540000 125.435000 ;
      RECT 16.805000 125.410000 24.540000 125.435000 ;
      RECT 16.805000 136.880000 59.620000 136.950000 ;
      RECT 16.805000 136.880000 59.620000 136.950000 ;
      RECT 16.805000 148.435000 57.370000 148.505000 ;
      RECT 16.805000 182.765000 60.760000 182.835000 ;
      RECT 16.820000  36.815000 54.390000  36.885000 ;
      RECT 16.820000  36.815000 54.390000  36.885000 ;
      RECT 16.820000  43.010000 60.830000  43.080000 ;
      RECT 16.820000  43.010000 60.830000  43.080000 ;
      RECT 16.830000 182.740000 60.830000 182.765000 ;
      RECT 16.835000  28.080000 57.840000  28.150000 ;
      RECT 16.835000  28.080000 57.840000  28.150000 ;
      RECT 16.835000  90.705000 59.850000  90.775000 ;
      RECT 16.835000  90.705000 59.850000  90.775000 ;
      RECT 16.840000 113.740000 59.725000 113.810000 ;
      RECT 16.840000 113.740000 59.725000 113.810000 ;
      RECT 16.850000  79.505000 24.540000  79.575000 ;
      RECT 16.850000  79.505000 24.540000  79.575000 ;
      RECT 16.850000  79.505000 57.510000  79.575000 ;
      RECT 16.850000 102.505000 24.540000 102.575000 ;
      RECT 16.850000 102.505000 24.540000 102.575000 ;
      RECT 16.850000 102.505000 57.510000 102.575000 ;
      RECT 16.855000 159.740000 59.775000 159.810000 ;
      RECT 16.855000 159.740000 59.775000 159.810000 ;
      RECT 16.870000  67.670000 59.825000  67.740000 ;
      RECT 16.870000  67.670000 59.825000  67.740000 ;
      RECT 16.870000 171.505000 57.520000 171.575000 ;
      RECT 16.875000  56.505000 57.480000  56.575000 ;
      RECT 16.875000 125.435000 24.540000 125.505000 ;
      RECT 16.875000 125.435000 24.540000 125.505000 ;
      RECT 16.875000 125.435000 57.440000 125.505000 ;
      RECT 16.875000 136.810000 59.690000 136.880000 ;
      RECT 16.875000 136.810000 59.690000 136.880000 ;
      RECT 16.875000 148.505000 57.440000 148.575000 ;
      RECT 16.890000  36.885000 54.390000  36.955000 ;
      RECT 16.890000  36.885000 54.390000  36.955000 ;
      RECT 16.890000  42.940000 60.830000  43.010000 ;
      RECT 16.890000  42.940000 60.830000  43.010000 ;
      RECT 16.900000 182.670000 60.830000 182.740000 ;
      RECT 16.905000  28.010000 57.770000  28.080000 ;
      RECT 16.905000  28.010000 57.770000  28.080000 ;
      RECT 16.905000  90.635000 59.920000  90.705000 ;
      RECT 16.905000  90.635000 59.920000  90.705000 ;
      RECT 16.910000 113.670000 59.795000 113.740000 ;
      RECT 16.910000 113.670000 59.795000 113.740000 ;
      RECT 16.920000  79.575000 24.540000  79.645000 ;
      RECT 16.920000  79.575000 24.540000  79.645000 ;
      RECT 16.920000  79.575000 57.580000  79.645000 ;
      RECT 16.920000 102.575000 24.540000 102.645000 ;
      RECT 16.920000 102.575000 24.540000 102.645000 ;
      RECT 16.920000 102.575000 57.580000 102.645000 ;
      RECT 16.925000 159.670000 59.845000 159.740000 ;
      RECT 16.925000 159.670000 59.845000 159.740000 ;
      RECT 16.940000  67.600000 59.895000  67.670000 ;
      RECT 16.940000  67.600000 59.895000  67.670000 ;
      RECT 16.940000 171.575000 57.590000 171.645000 ;
      RECT 16.945000  56.575000 57.550000  56.645000 ;
      RECT 16.945000 125.505000 24.540000 125.575000 ;
      RECT 16.945000 125.505000 24.540000 125.575000 ;
      RECT 16.945000 125.505000 57.510000 125.575000 ;
      RECT 16.945000 136.740000 59.760000 136.810000 ;
      RECT 16.945000 136.740000 59.760000 136.810000 ;
      RECT 16.945000 148.575000 57.510000 148.645000 ;
      RECT 16.960000  36.955000 54.390000  37.025000 ;
      RECT 16.960000  36.955000 54.390000  37.025000 ;
      RECT 16.960000  42.870000 60.830000  42.940000 ;
      RECT 16.960000  42.870000 60.830000  42.940000 ;
      RECT 16.970000 182.600000 60.830000 182.670000 ;
      RECT 16.975000  27.940000 57.700000  28.010000 ;
      RECT 16.975000  27.940000 57.700000  28.010000 ;
      RECT 16.975000  90.565000 59.990000  90.635000 ;
      RECT 16.975000  90.565000 59.990000  90.635000 ;
      RECT 16.980000 113.600000 59.865000 113.670000 ;
      RECT 16.980000 113.600000 59.865000 113.670000 ;
      RECT 16.990000  79.645000 24.540000  79.715000 ;
      RECT 16.990000  79.645000 24.540000  79.715000 ;
      RECT 16.990000  79.645000 57.650000  79.715000 ;
      RECT 16.990000 102.645000 24.540000 102.715000 ;
      RECT 16.990000 102.645000 24.540000 102.715000 ;
      RECT 16.990000 102.645000 57.650000 102.715000 ;
      RECT 16.995000 159.600000 59.915000 159.670000 ;
      RECT 16.995000 159.600000 59.915000 159.670000 ;
      RECT 17.010000  67.530000 59.965000  67.600000 ;
      RECT 17.010000  67.530000 59.965000  67.600000 ;
      RECT 17.010000 171.645000 57.660000 171.715000 ;
      RECT 17.015000  56.645000 57.620000  56.715000 ;
      RECT 17.015000 125.575000 24.540000 125.645000 ;
      RECT 17.015000 125.575000 24.540000 125.645000 ;
      RECT 17.015000 125.575000 57.580000 125.645000 ;
      RECT 17.015000 136.670000 59.830000 136.740000 ;
      RECT 17.015000 136.670000 59.830000 136.740000 ;
      RECT 17.015000 148.645000 57.580000 148.715000 ;
      RECT 17.030000  37.025000 54.390000  37.095000 ;
      RECT 17.030000  37.025000 54.390000  37.095000 ;
      RECT 17.030000  42.800000 60.830000  42.870000 ;
      RECT 17.030000  42.800000 60.830000  42.870000 ;
      RECT 17.040000 182.530000 60.830000 182.600000 ;
      RECT 17.045000  27.870000 57.630000  27.940000 ;
      RECT 17.045000  27.870000 57.630000  27.940000 ;
      RECT 17.045000  90.495000 60.060000  90.565000 ;
      RECT 17.045000  90.495000 60.060000  90.565000 ;
      RECT 17.050000 113.530000 59.935000 113.600000 ;
      RECT 17.050000 113.530000 59.935000 113.600000 ;
      RECT 17.060000  79.715000 24.540000  79.785000 ;
      RECT 17.060000  79.715000 24.540000  79.785000 ;
      RECT 17.060000  79.715000 57.720000  79.785000 ;
      RECT 17.060000 102.715000 24.540000 102.785000 ;
      RECT 17.060000 102.715000 24.540000 102.785000 ;
      RECT 17.060000 102.715000 57.720000 102.785000 ;
      RECT 17.065000 159.530000 59.985000 159.600000 ;
      RECT 17.065000 159.530000 59.985000 159.600000 ;
      RECT 17.080000  67.460000 60.035000  67.530000 ;
      RECT 17.080000  67.460000 60.035000  67.530000 ;
      RECT 17.080000 171.715000 57.730000 171.785000 ;
      RECT 17.085000  56.715000 57.690000  56.785000 ;
      RECT 17.085000 125.645000 24.540000 125.715000 ;
      RECT 17.085000 125.645000 24.540000 125.715000 ;
      RECT 17.085000 125.645000 57.650000 125.715000 ;
      RECT 17.085000 136.600000 59.900000 136.670000 ;
      RECT 17.085000 136.600000 59.900000 136.670000 ;
      RECT 17.085000 148.715000 57.650000 148.785000 ;
      RECT 17.100000  37.095000 54.390000  37.165000 ;
      RECT 17.100000  37.095000 54.390000  37.165000 ;
      RECT 17.100000  42.730000 60.830000  42.800000 ;
      RECT 17.100000  42.730000 60.830000  42.800000 ;
      RECT 17.110000 182.460000 60.830000 182.530000 ;
      RECT 17.115000  27.800000 57.560000  27.870000 ;
      RECT 17.115000  27.800000 57.560000  27.870000 ;
      RECT 17.115000  90.425000 60.130000  90.495000 ;
      RECT 17.115000  90.425000 60.130000  90.495000 ;
      RECT 17.120000 113.460000 60.005000 113.530000 ;
      RECT 17.120000 113.460000 60.005000 113.530000 ;
      RECT 17.130000  79.785000 24.540000  79.855000 ;
      RECT 17.130000  79.785000 24.540000  79.855000 ;
      RECT 17.130000  79.785000 57.790000  79.855000 ;
      RECT 17.130000 102.785000 24.540000 102.855000 ;
      RECT 17.130000 102.785000 24.540000 102.855000 ;
      RECT 17.130000 102.785000 57.790000 102.855000 ;
      RECT 17.135000 159.460000 60.055000 159.530000 ;
      RECT 17.135000 159.460000 60.055000 159.530000 ;
      RECT 17.150000  67.390000 60.105000  67.460000 ;
      RECT 17.150000  67.390000 60.105000  67.460000 ;
      RECT 17.150000 171.785000 57.800000 171.855000 ;
      RECT 17.155000  56.785000 57.760000  56.855000 ;
      RECT 17.155000 125.715000 24.540000 125.785000 ;
      RECT 17.155000 125.715000 24.540000 125.785000 ;
      RECT 17.155000 125.715000 57.720000 125.785000 ;
      RECT 17.155000 136.530000 59.970000 136.600000 ;
      RECT 17.155000 136.530000 59.970000 136.600000 ;
      RECT 17.155000 148.785000 57.720000 148.855000 ;
      RECT 17.170000  37.165000 54.390000  37.235000 ;
      RECT 17.170000  37.165000 54.390000  37.235000 ;
      RECT 17.170000  42.660000 60.830000  42.730000 ;
      RECT 17.170000  42.660000 60.830000  42.730000 ;
      RECT 17.170000  42.660000 60.970000  43.760000 ;
      RECT 17.180000 182.390000 60.830000 182.460000 ;
      RECT 17.185000  27.730000 57.490000  27.800000 ;
      RECT 17.185000  27.730000 57.490000  27.800000 ;
      RECT 17.185000  90.355000 60.200000  90.425000 ;
      RECT 17.185000  90.355000 60.200000  90.425000 ;
      RECT 17.190000 113.390000 60.075000 113.460000 ;
      RECT 17.190000 113.390000 60.075000 113.460000 ;
      RECT 17.200000  79.855000 24.540000  79.925000 ;
      RECT 17.200000  79.855000 24.540000  79.925000 ;
      RECT 17.200000  79.855000 57.860000  79.925000 ;
      RECT 17.200000 102.855000 24.540000 102.925000 ;
      RECT 17.200000 102.855000 24.540000 102.925000 ;
      RECT 17.200000 102.855000 57.860000 102.925000 ;
      RECT 17.205000 159.390000 60.125000 159.460000 ;
      RECT 17.205000 159.390000 60.125000 159.460000 ;
      RECT 17.220000  67.320000 60.175000  67.390000 ;
      RECT 17.220000  67.320000 60.175000  67.390000 ;
      RECT 17.220000 171.855000 57.870000 171.925000 ;
      RECT 17.225000  56.855000 57.830000  56.925000 ;
      RECT 17.225000 125.785000 24.540000 125.855000 ;
      RECT 17.225000 125.785000 24.540000 125.855000 ;
      RECT 17.225000 125.785000 57.790000 125.855000 ;
      RECT 17.225000 136.460000 60.040000 136.530000 ;
      RECT 17.225000 136.460000 60.040000 136.530000 ;
      RECT 17.225000 148.855000 57.790000 148.925000 ;
      RECT 17.240000  37.235000 54.390000  37.305000 ;
      RECT 17.240000  37.235000 54.390000  37.305000 ;
      RECT 17.250000 182.320000 60.830000 182.390000 ;
      RECT 17.255000  27.660000 57.420000  27.730000 ;
      RECT 17.255000  27.660000 57.420000  27.730000 ;
      RECT 17.255000  90.285000 60.270000  90.355000 ;
      RECT 17.255000  90.285000 60.270000  90.355000 ;
      RECT 17.260000 113.320000 60.145000 113.390000 ;
      RECT 17.260000 113.320000 60.145000 113.390000 ;
      RECT 17.270000  79.925000 24.540000  79.995000 ;
      RECT 17.270000  79.925000 24.540000  79.995000 ;
      RECT 17.270000  79.925000 57.930000  79.995000 ;
      RECT 17.270000 102.925000 24.540000 102.995000 ;
      RECT 17.270000 102.925000 24.540000 102.995000 ;
      RECT 17.270000 102.925000 57.930000 102.995000 ;
      RECT 17.275000 159.320000 60.195000 159.390000 ;
      RECT 17.275000 159.320000 60.195000 159.390000 ;
      RECT 17.290000  67.250000 60.245000  67.320000 ;
      RECT 17.290000  67.250000 60.245000  67.320000 ;
      RECT 17.290000 171.925000 57.940000 171.995000 ;
      RECT 17.295000  56.925000 57.900000  56.995000 ;
      RECT 17.295000 125.855000 24.540000 125.925000 ;
      RECT 17.295000 125.855000 24.540000 125.925000 ;
      RECT 17.295000 125.855000 57.860000 125.925000 ;
      RECT 17.295000 136.390000 60.110000 136.460000 ;
      RECT 17.295000 136.390000 60.110000 136.460000 ;
      RECT 17.295000 148.925000 57.860000 148.995000 ;
      RECT 17.310000  37.305000 54.390000  37.375000 ;
      RECT 17.310000  37.305000 54.390000  37.375000 ;
      RECT 17.320000 182.250000 60.830000 182.320000 ;
      RECT 17.325000  27.590000 57.350000  27.660000 ;
      RECT 17.325000  27.590000 57.350000  27.660000 ;
      RECT 17.325000  90.215000 60.340000  90.285000 ;
      RECT 17.325000  90.215000 60.340000  90.285000 ;
      RECT 17.330000 113.250000 60.215000 113.320000 ;
      RECT 17.330000 113.250000 60.215000 113.320000 ;
      RECT 17.340000  79.995000 24.540000  80.065000 ;
      RECT 17.340000  79.995000 24.540000  80.065000 ;
      RECT 17.340000  79.995000 58.000000  80.065000 ;
      RECT 17.340000 102.995000 24.540000 103.065000 ;
      RECT 17.340000 102.995000 24.540000 103.065000 ;
      RECT 17.340000 102.995000 58.000000 103.065000 ;
      RECT 17.345000 159.250000 60.265000 159.320000 ;
      RECT 17.345000 159.250000 60.265000 159.320000 ;
      RECT 17.360000  67.180000 60.315000  67.250000 ;
      RECT 17.360000  67.180000 60.315000  67.250000 ;
      RECT 17.360000 171.995000 58.010000 172.065000 ;
      RECT 17.365000  56.995000 57.970000  57.065000 ;
      RECT 17.365000 125.925000 24.540000 125.995000 ;
      RECT 17.365000 125.925000 24.540000 125.995000 ;
      RECT 17.365000 125.925000 57.930000 125.995000 ;
      RECT 17.365000 136.320000 60.180000 136.390000 ;
      RECT 17.365000 136.320000 60.180000 136.390000 ;
      RECT 17.365000 148.995000 57.930000 149.065000 ;
      RECT 17.380000  37.375000 54.390000  37.445000 ;
      RECT 17.380000  37.375000 54.390000  37.445000 ;
      RECT 17.390000 182.180000 60.830000 182.250000 ;
      RECT 17.395000  27.520000 57.280000  27.590000 ;
      RECT 17.395000  27.520000 57.280000  27.590000 ;
      RECT 17.395000  90.145000 60.410000  90.215000 ;
      RECT 17.395000  90.145000 60.410000  90.215000 ;
      RECT 17.400000 113.180000 60.285000 113.250000 ;
      RECT 17.400000 113.180000 60.285000 113.250000 ;
      RECT 17.410000  80.065000 24.540000  80.135000 ;
      RECT 17.410000  80.065000 24.540000  80.135000 ;
      RECT 17.410000  80.065000 58.070000  80.135000 ;
      RECT 17.410000 103.065000 24.540000 103.135000 ;
      RECT 17.410000 103.065000 24.540000 103.135000 ;
      RECT 17.410000 103.065000 58.070000 103.135000 ;
      RECT 17.415000 159.180000 60.335000 159.250000 ;
      RECT 17.415000 159.180000 60.335000 159.250000 ;
      RECT 17.430000  67.110000 60.385000  67.180000 ;
      RECT 17.430000  67.110000 60.385000  67.180000 ;
      RECT 17.430000 172.065000 58.080000 172.135000 ;
      RECT 17.435000  57.065000 58.040000  57.135000 ;
      RECT 17.435000 125.995000 24.540000 126.065000 ;
      RECT 17.435000 125.995000 24.540000 126.065000 ;
      RECT 17.435000 125.995000 58.000000 126.065000 ;
      RECT 17.435000 136.250000 60.250000 136.320000 ;
      RECT 17.435000 136.250000 60.250000 136.320000 ;
      RECT 17.435000 149.065000 58.000000 149.135000 ;
      RECT 17.450000  37.445000 54.390000  37.515000 ;
      RECT 17.450000  37.445000 54.390000  37.515000 ;
      RECT 17.460000 182.110000 60.830000 182.180000 ;
      RECT 17.465000  27.450000 57.210000  27.520000 ;
      RECT 17.465000  27.450000 57.210000  27.520000 ;
      RECT 17.465000  90.075000 60.480000  90.145000 ;
      RECT 17.465000  90.075000 60.480000  90.145000 ;
      RECT 17.470000 113.110000 60.355000 113.180000 ;
      RECT 17.470000 113.110000 60.355000 113.180000 ;
      RECT 17.480000  80.135000 24.540000  80.205000 ;
      RECT 17.480000  80.135000 24.540000  80.205000 ;
      RECT 17.480000  80.135000 58.140000  80.205000 ;
      RECT 17.480000 103.135000 24.540000 103.205000 ;
      RECT 17.480000 103.135000 24.540000 103.205000 ;
      RECT 17.480000 103.135000 58.140000 103.205000 ;
      RECT 17.485000 159.110000 60.405000 159.180000 ;
      RECT 17.485000 159.110000 60.405000 159.180000 ;
      RECT 17.500000  67.040000 60.455000  67.110000 ;
      RECT 17.500000  67.040000 60.455000  67.110000 ;
      RECT 17.500000 172.135000 58.150000 172.205000 ;
      RECT 17.505000  57.135000 58.110000  57.205000 ;
      RECT 17.505000 126.065000 24.540000 126.135000 ;
      RECT 17.505000 126.065000 24.540000 126.135000 ;
      RECT 17.505000 126.065000 58.070000 126.135000 ;
      RECT 17.505000 136.180000 60.320000 136.250000 ;
      RECT 17.505000 136.180000 60.320000 136.250000 ;
      RECT 17.505000 149.135000 58.070000 149.205000 ;
      RECT 17.520000  37.515000 54.390000  37.585000 ;
      RECT 17.520000  37.515000 54.390000  37.585000 ;
      RECT 17.530000 182.040000 60.830000 182.110000 ;
      RECT 17.535000  27.380000 57.140000  27.450000 ;
      RECT 17.535000  27.380000 57.140000  27.450000 ;
      RECT 17.535000  90.005000 60.550000  90.075000 ;
      RECT 17.535000  90.005000 60.550000  90.075000 ;
      RECT 17.540000 113.040000 60.425000 113.110000 ;
      RECT 17.540000 113.040000 60.425000 113.110000 ;
      RECT 17.550000  80.205000 24.540000  80.275000 ;
      RECT 17.550000  80.205000 24.540000  80.275000 ;
      RECT 17.550000  80.205000 58.210000  80.275000 ;
      RECT 17.550000 103.205000 24.540000 103.275000 ;
      RECT 17.550000 103.205000 24.540000 103.275000 ;
      RECT 17.550000 103.205000 58.210000 103.275000 ;
      RECT 17.555000 159.040000 60.475000 159.110000 ;
      RECT 17.555000 159.040000 60.475000 159.110000 ;
      RECT 17.570000  66.970000 60.525000  67.040000 ;
      RECT 17.570000  66.970000 60.525000  67.040000 ;
      RECT 17.570000 172.205000 58.220000 172.275000 ;
      RECT 17.575000  57.205000 58.180000  57.275000 ;
      RECT 17.575000 126.135000 24.540000 126.205000 ;
      RECT 17.575000 126.135000 24.540000 126.205000 ;
      RECT 17.575000 126.135000 58.140000 126.205000 ;
      RECT 17.575000 136.110000 60.390000 136.180000 ;
      RECT 17.575000 136.110000 60.390000 136.180000 ;
      RECT 17.575000 149.205000 58.140000 149.275000 ;
      RECT 17.590000  37.585000 54.390000  37.655000 ;
      RECT 17.590000  37.585000 54.390000  37.655000 ;
      RECT 17.600000 181.970000 60.830000 182.040000 ;
      RECT 17.605000  27.310000 57.070000  27.380000 ;
      RECT 17.605000  27.310000 57.070000  27.380000 ;
      RECT 17.605000  89.935000 60.620000  90.005000 ;
      RECT 17.605000  89.935000 60.620000  90.005000 ;
      RECT 17.610000 112.970000 60.495000 113.040000 ;
      RECT 17.610000 112.970000 60.495000 113.040000 ;
      RECT 17.620000  80.275000 24.540000  80.345000 ;
      RECT 17.620000  80.275000 24.540000  80.345000 ;
      RECT 17.620000  80.275000 58.280000  80.345000 ;
      RECT 17.620000 103.275000 24.540000 103.345000 ;
      RECT 17.620000 103.275000 24.540000 103.345000 ;
      RECT 17.620000 103.275000 58.280000 103.345000 ;
      RECT 17.625000 158.970000 60.545000 159.040000 ;
      RECT 17.625000 158.970000 60.545000 159.040000 ;
      RECT 17.640000  66.900000 60.595000  66.970000 ;
      RECT 17.640000  66.900000 60.595000  66.970000 ;
      RECT 17.640000 172.275000 58.290000 172.345000 ;
      RECT 17.645000  57.275000 58.250000  57.345000 ;
      RECT 17.645000 126.205000 24.540000 126.275000 ;
      RECT 17.645000 126.205000 24.540000 126.275000 ;
      RECT 17.645000 126.205000 58.210000 126.275000 ;
      RECT 17.645000 136.040000 60.460000 136.110000 ;
      RECT 17.645000 136.040000 60.460000 136.110000 ;
      RECT 17.645000 149.275000 58.210000 149.345000 ;
      RECT 17.660000  37.655000 54.390000  37.725000 ;
      RECT 17.660000  37.655000 54.390000  37.725000 ;
      RECT 17.670000 181.900000 60.830000 181.970000 ;
      RECT 17.675000  27.240000 57.000000  27.310000 ;
      RECT 17.675000  27.240000 57.000000  27.310000 ;
      RECT 17.675000  89.865000 60.690000  89.935000 ;
      RECT 17.675000  89.865000 60.690000  89.935000 ;
      RECT 17.680000 112.900000 60.565000 112.970000 ;
      RECT 17.680000 112.900000 60.565000 112.970000 ;
      RECT 17.690000  80.345000 24.540000  80.415000 ;
      RECT 17.690000  80.345000 24.540000  80.415000 ;
      RECT 17.690000  80.345000 58.350000  80.415000 ;
      RECT 17.690000  89.850000 57.680000  93.140000 ;
      RECT 17.690000 103.345000 24.540000 103.415000 ;
      RECT 17.690000 103.345000 24.540000 103.415000 ;
      RECT 17.690000 103.345000 58.350000 103.415000 ;
      RECT 17.695000 158.900000 60.615000 158.970000 ;
      RECT 17.695000 158.900000 60.615000 158.970000 ;
      RECT 17.710000  66.830000 60.665000  66.900000 ;
      RECT 17.710000  66.830000 60.665000  66.900000 ;
      RECT 17.710000 172.345000 58.360000 172.415000 ;
      RECT 17.715000  57.345000 58.320000  57.415000 ;
      RECT 17.715000 126.275000 24.540000 126.345000 ;
      RECT 17.715000 126.275000 24.540000 126.345000 ;
      RECT 17.715000 126.275000 58.280000 126.345000 ;
      RECT 17.715000 135.970000 60.530000 136.040000 ;
      RECT 17.715000 135.970000 60.530000 136.040000 ;
      RECT 17.715000 149.345000 58.280000 149.415000 ;
      RECT 17.730000  37.725000 54.390000  37.795000 ;
      RECT 17.730000  37.725000 54.390000  37.795000 ;
      RECT 17.740000 181.830000 60.830000 181.900000 ;
      RECT 17.745000  27.170000 56.930000  27.240000 ;
      RECT 17.745000  27.170000 56.930000  27.240000 ;
      RECT 17.745000  89.795000 60.760000  89.865000 ;
      RECT 17.745000  89.795000 60.760000  89.865000 ;
      RECT 17.750000  66.790000 57.620000  70.140000 ;
      RECT 17.750000  89.790000 60.830000  89.795000 ;
      RECT 17.750000  89.790000 60.830000  89.795000 ;
      RECT 17.750000 112.830000 60.635000 112.900000 ;
      RECT 17.750000 112.830000 60.635000 112.900000 ;
      RECT 17.760000  80.415000 24.540000  80.485000 ;
      RECT 17.760000  80.415000 24.540000  80.485000 ;
      RECT 17.760000  80.415000 58.420000  80.485000 ;
      RECT 17.760000 103.415000 24.540000 103.485000 ;
      RECT 17.760000 103.415000 24.540000 103.485000 ;
      RECT 17.760000 103.415000 58.420000 103.485000 ;
      RECT 17.765000  89.775000 60.830000  89.790000 ;
      RECT 17.765000  89.775000 60.830000  89.790000 ;
      RECT 17.765000 158.830000 60.685000 158.900000 ;
      RECT 17.765000 158.830000 60.685000 158.900000 ;
      RECT 17.775000  80.485000 24.540000  80.500000 ;
      RECT 17.775000  80.485000 24.540000  80.500000 ;
      RECT 17.775000  80.485000 58.490000  80.500000 ;
      RECT 17.775000 103.485000 24.540000 103.500000 ;
      RECT 17.775000 103.485000 24.540000 103.500000 ;
      RECT 17.775000 103.485000 58.490000 103.500000 ;
      RECT 17.780000  66.760000 60.735000  66.830000 ;
      RECT 17.780000  66.760000 60.735000  66.830000 ;
      RECT 17.780000  66.760000 60.970000  66.790000 ;
      RECT 17.780000  89.760000 60.830000  89.775000 ;
      RECT 17.780000  89.760000 60.830000  89.775000 ;
      RECT 17.780000  89.760000 60.970000  89.850000 ;
      RECT 17.780000 172.415000 58.430000 172.485000 ;
      RECT 17.785000  57.415000 58.390000  57.485000 ;
      RECT 17.785000 126.345000 24.540000 126.415000 ;
      RECT 17.785000 126.345000 24.540000 126.415000 ;
      RECT 17.785000 126.345000 58.350000 126.415000 ;
      RECT 17.785000 135.900000 60.600000 135.970000 ;
      RECT 17.785000 135.900000 60.600000 135.970000 ;
      RECT 17.785000 149.415000 58.350000 149.485000 ;
      RECT 17.785000 158.810000 57.585000 162.195000 ;
      RECT 17.795000 172.485000 58.500000 172.500000 ;
      RECT 17.800000  37.795000 54.390000  37.865000 ;
      RECT 17.800000  37.795000 54.390000  37.865000 ;
      RECT 17.800000  57.485000 58.460000  57.500000 ;
      RECT 17.800000 149.485000 58.420000 149.500000 ;
      RECT 17.810000 181.760000 60.830000 181.830000 ;
      RECT 17.810000 181.760000 60.970000 182.820000 ;
      RECT 17.815000  27.100000 56.860000  27.170000 ;
      RECT 17.815000  27.100000 56.860000  27.170000 ;
      RECT 17.820000 112.760000 57.550000 116.180000 ;
      RECT 17.820000 112.760000 60.705000 112.830000 ;
      RECT 17.820000 112.760000 60.705000 112.830000 ;
      RECT 17.821000 112.760000 60.970000 112.762000 ;
      RECT 17.835000 158.760000 60.755000 158.830000 ;
      RECT 17.835000 158.760000 60.755000 158.830000 ;
      RECT 17.835000 158.760000 60.970000 158.810000 ;
      RECT 17.855000 126.415000 24.540000 126.485000 ;
      RECT 17.855000 126.415000 24.540000 126.485000 ;
      RECT 17.855000 126.415000 58.420000 126.485000 ;
      RECT 17.855000 135.830000 60.670000 135.900000 ;
      RECT 17.855000 135.830000 60.670000 135.900000 ;
      RECT 17.870000  37.865000 54.390000  37.935000 ;
      RECT 17.870000  37.865000 54.390000  37.935000 ;
      RECT 17.870000 126.485000 24.540000 126.500000 ;
      RECT 17.870000 126.485000 24.540000 126.500000 ;
      RECT 17.870000 126.485000 58.490000 126.500000 ;
      RECT 17.885000  27.030000 56.790000  27.100000 ;
      RECT 17.885000  27.030000 56.790000  27.100000 ;
      RECT 17.890000 135.795000 57.480000 139.285000 ;
      RECT 17.925000 135.760000 60.740000 135.830000 ;
      RECT 17.925000 135.760000 60.740000 135.830000 ;
      RECT 17.925000 135.760000 60.970000 135.795000 ;
      RECT 17.940000  37.935000 54.390000  38.005000 ;
      RECT 17.940000  37.935000 54.390000  38.005000 ;
      RECT 17.955000  26.960000 56.720000  27.030000 ;
      RECT 17.955000  26.960000 56.720000  27.030000 ;
      RECT 18.010000  38.005000 54.390000  38.075000 ;
      RECT 18.010000  38.005000 54.390000  38.075000 ;
      RECT 18.025000  26.890000 56.650000  26.960000 ;
      RECT 18.025000  26.890000 56.650000  26.960000 ;
      RECT 18.075000  38.075000 54.390000  38.140000 ;
      RECT 18.075000  38.075000 54.390000  38.140000 ;
      RECT 18.095000  26.820000 56.580000  26.890000 ;
      RECT 18.095000  26.820000 56.580000  26.890000 ;
      RECT 18.135000  38.195000 52.655000  40.070000 ;
      RECT 18.145000  38.140000 54.320000  38.210000 ;
      RECT 18.145000  38.140000 54.320000  38.210000 ;
      RECT 18.165000  26.750000 56.510000  26.820000 ;
      RECT 18.165000  26.750000 56.510000  26.820000 ;
      RECT 18.215000  38.210000 54.250000  38.280000 ;
      RECT 18.215000  38.210000 54.250000  38.280000 ;
      RECT 18.235000  26.680000 56.440000  26.750000 ;
      RECT 18.235000  26.680000 56.440000  26.750000 ;
      RECT 18.285000  38.280000 54.180000  38.350000 ;
      RECT 18.285000  38.280000 54.180000  38.350000 ;
      RECT 18.305000  26.610000 56.370000  26.680000 ;
      RECT 18.305000  26.610000 56.370000  26.680000 ;
      RECT 18.355000  38.350000 54.110000  38.420000 ;
      RECT 18.355000  38.350000 54.110000  38.420000 ;
      RECT 18.375000  26.540000 56.300000  26.610000 ;
      RECT 18.375000  26.540000 56.300000  26.610000 ;
      RECT 18.425000  38.420000 54.040000  38.490000 ;
      RECT 18.425000  38.420000 54.040000  38.490000 ;
      RECT 18.445000  26.470000 56.230000  26.540000 ;
      RECT 18.445000  26.470000 56.230000  26.540000 ;
      RECT 18.495000  38.490000 53.970000  38.560000 ;
      RECT 18.495000  38.490000 53.970000  38.560000 ;
      RECT 18.515000  26.400000 56.160000  26.470000 ;
      RECT 18.515000  26.400000 56.160000  26.470000 ;
      RECT 18.565000  38.560000 53.900000  38.630000 ;
      RECT 18.565000  38.560000 53.900000  38.630000 ;
      RECT 18.585000  26.330000 56.090000  26.400000 ;
      RECT 18.585000  26.330000 56.090000  26.400000 ;
      RECT 18.635000  38.630000 53.830000  38.700000 ;
      RECT 18.635000  38.630000 53.830000  38.700000 ;
      RECT 18.655000  26.260000 56.020000  26.330000 ;
      RECT 18.655000  26.260000 56.020000  26.330000 ;
      RECT 18.705000  38.700000 53.760000  38.770000 ;
      RECT 18.705000  38.700000 53.760000  38.770000 ;
      RECT 18.725000  26.190000 55.950000  26.260000 ;
      RECT 18.725000  26.190000 55.950000  26.260000 ;
      RECT 18.775000  38.770000 53.690000  38.840000 ;
      RECT 18.775000  38.770000 53.690000  38.840000 ;
      RECT 18.795000  26.120000 55.880000  26.190000 ;
      RECT 18.795000  26.120000 55.880000  26.190000 ;
      RECT 18.845000  38.840000 53.620000  38.910000 ;
      RECT 18.845000  38.840000 53.620000  38.910000 ;
      RECT 18.865000  26.050000 55.810000  26.120000 ;
      RECT 18.865000  26.050000 55.810000  26.120000 ;
      RECT 18.915000  38.910000 53.550000  38.980000 ;
      RECT 18.915000  38.910000 53.550000  38.980000 ;
      RECT 18.935000  25.980000 55.740000  26.050000 ;
      RECT 18.935000  25.980000 55.740000  26.050000 ;
      RECT 18.935000  25.980000 59.390000  29.430000 ;
      RECT 18.985000  38.980000 53.480000  39.050000 ;
      RECT 18.985000  38.980000 53.480000  39.050000 ;
      RECT 19.055000  39.050000 53.410000  39.120000 ;
      RECT 19.055000  39.050000 53.410000  39.120000 ;
      RECT 19.125000  39.120000 53.340000  39.190000 ;
      RECT 19.125000  39.120000 53.340000  39.190000 ;
      RECT 19.195000  39.190000 53.270000  39.260000 ;
      RECT 19.195000  39.190000 53.270000  39.260000 ;
      RECT 19.265000  39.260000 53.200000  39.330000 ;
      RECT 19.265000  39.260000 53.200000  39.330000 ;
      RECT 19.335000  39.330000 53.130000  39.400000 ;
      RECT 19.335000  39.330000 53.130000  39.400000 ;
      RECT 19.405000  39.400000 53.060000  39.470000 ;
      RECT 19.405000  39.400000 53.060000  39.470000 ;
      RECT 19.475000  39.470000 52.990000  39.540000 ;
      RECT 19.475000  39.470000 52.990000  39.540000 ;
      RECT 19.545000  39.540000 52.920000  39.610000 ;
      RECT 19.545000  39.540000 52.920000  39.610000 ;
      RECT 19.615000  39.610000 52.850000  39.680000 ;
      RECT 19.615000  39.610000 52.850000  39.680000 ;
      RECT 19.685000  39.680000 52.780000  39.750000 ;
      RECT 19.685000  39.680000 52.780000  39.750000 ;
      RECT 19.755000  39.750000 52.710000  39.820000 ;
      RECT 19.755000  39.750000 52.710000  39.820000 ;
      RECT 19.825000  39.820000 52.640000  39.890000 ;
      RECT 19.825000  39.820000 52.640000  39.890000 ;
      RECT 19.895000  39.890000 52.570000  39.960000 ;
      RECT 19.895000  39.890000 52.570000  39.960000 ;
      RECT 19.965000  39.960000 52.500000  40.030000 ;
      RECT 19.965000  39.960000 52.500000  40.030000 ;
      RECT 20.005000  40.030000 52.460000  40.070000 ;
      RECT 20.005000  40.030000 52.460000  40.070000 ;
      RECT 20.400000  40.070000 52.515000  40.210000 ;
      RECT 22.850000  42.520000 60.970000  42.660000 ;
      RECT 24.675000   0.000000 25.615000   0.815000 ;
      RECT 24.675000   0.000000 25.755000   0.675000 ;
      RECT 24.675000   0.675000 50.250000   8.480000 ;
      RECT 24.675000   0.815000 50.110000   8.480000 ;
      RECT 24.675000   8.480000 50.250000   8.565000 ;
      RECT 24.690000   8.480000 50.110000   8.495000 ;
      RECT 24.690000   8.480000 50.110000   8.495000 ;
      RECT 24.705000   8.495000 50.110000   8.510000 ;
      RECT 24.705000   8.495000 50.110000   8.510000 ;
      RECT 24.765000   8.565000 46.695000  12.120000 ;
      RECT 24.775000   8.510000 50.040000   8.580000 ;
      RECT 24.775000   8.510000 50.040000   8.580000 ;
      RECT 24.845000   8.580000 49.970000   8.650000 ;
      RECT 24.845000   8.580000 49.970000   8.650000 ;
      RECT 24.915000   8.650000 49.900000   8.720000 ;
      RECT 24.915000   8.650000 49.900000   8.720000 ;
      RECT 24.985000   8.720000 49.830000   8.790000 ;
      RECT 24.985000   8.720000 49.830000   8.790000 ;
      RECT 25.055000   8.790000 49.760000   8.860000 ;
      RECT 25.055000   8.790000 49.760000   8.860000 ;
      RECT 25.125000   8.860000 49.690000   8.930000 ;
      RECT 25.125000   8.860000 49.690000   8.930000 ;
      RECT 25.195000   8.930000 49.620000   9.000000 ;
      RECT 25.195000   8.930000 49.620000   9.000000 ;
      RECT 25.265000   9.000000 49.550000   9.070000 ;
      RECT 25.265000   9.000000 49.550000   9.070000 ;
      RECT 25.335000   9.070000 49.480000   9.140000 ;
      RECT 25.335000   9.070000 49.480000   9.140000 ;
      RECT 25.405000   9.140000 49.410000   9.210000 ;
      RECT 25.405000   9.140000 49.410000   9.210000 ;
      RECT 25.475000   9.210000 49.340000   9.280000 ;
      RECT 25.475000   9.210000 49.340000   9.280000 ;
      RECT 25.545000   9.280000 49.270000   9.350000 ;
      RECT 25.545000   9.280000 49.270000   9.350000 ;
      RECT 25.615000   9.350000 49.200000   9.420000 ;
      RECT 25.615000   9.350000 49.200000   9.420000 ;
      RECT 25.685000   9.420000 49.130000   9.490000 ;
      RECT 25.685000   9.420000 49.130000   9.490000 ;
      RECT 25.755000   9.490000 49.060000   9.560000 ;
      RECT 25.755000   9.490000 49.060000   9.560000 ;
      RECT 25.825000   9.560000 48.990000   9.630000 ;
      RECT 25.825000   9.560000 48.990000   9.630000 ;
      RECT 25.895000   9.630000 48.920000   9.700000 ;
      RECT 25.895000   9.630000 48.920000   9.700000 ;
      RECT 25.965000   9.700000 48.850000   9.770000 ;
      RECT 25.965000   9.700000 48.850000   9.770000 ;
      RECT 26.035000   9.770000 48.780000   9.840000 ;
      RECT 26.035000   9.770000 48.780000   9.840000 ;
      RECT 26.105000   9.840000 48.710000   9.910000 ;
      RECT 26.105000   9.840000 48.710000   9.910000 ;
      RECT 26.175000   9.910000 48.640000   9.980000 ;
      RECT 26.175000   9.910000 48.640000   9.980000 ;
      RECT 26.245000   9.980000 48.570000  10.050000 ;
      RECT 26.245000   9.980000 48.570000  10.050000 ;
      RECT 26.315000  10.050000 48.500000  10.120000 ;
      RECT 26.315000  10.050000 48.500000  10.120000 ;
      RECT 26.385000  10.120000 48.430000  10.190000 ;
      RECT 26.385000  10.120000 48.430000  10.190000 ;
      RECT 26.455000  10.190000 48.360000  10.260000 ;
      RECT 26.455000  10.190000 48.360000  10.260000 ;
      RECT 26.525000  10.260000 48.290000  10.330000 ;
      RECT 26.525000  10.260000 48.290000  10.330000 ;
      RECT 26.595000  10.330000 48.220000  10.400000 ;
      RECT 26.595000  10.330000 48.220000  10.400000 ;
      RECT 26.665000  10.400000 48.150000  10.470000 ;
      RECT 26.665000  10.400000 48.150000  10.470000 ;
      RECT 26.735000  10.470000 48.080000  10.540000 ;
      RECT 26.735000  10.470000 48.080000  10.540000 ;
      RECT 26.805000  10.540000 48.010000  10.610000 ;
      RECT 26.805000  10.540000 48.010000  10.610000 ;
      RECT 26.875000  10.610000 47.940000  10.680000 ;
      RECT 26.875000  10.610000 47.940000  10.680000 ;
      RECT 26.945000  10.680000 47.870000  10.750000 ;
      RECT 26.945000  10.680000 47.870000  10.750000 ;
      RECT 27.015000  10.750000 47.800000  10.820000 ;
      RECT 27.015000  10.750000 47.800000  10.820000 ;
      RECT 27.085000  10.820000 47.730000  10.890000 ;
      RECT 27.085000  10.820000 47.730000  10.890000 ;
      RECT 27.155000  10.890000 47.660000  10.960000 ;
      RECT 27.155000  10.890000 47.660000  10.960000 ;
      RECT 27.225000  10.960000 47.590000  11.030000 ;
      RECT 27.225000  10.960000 47.590000  11.030000 ;
      RECT 27.295000  11.030000 47.520000  11.100000 ;
      RECT 27.295000  11.030000 47.520000  11.100000 ;
      RECT 27.365000  11.100000 47.450000  11.170000 ;
      RECT 27.365000  11.100000 47.450000  11.170000 ;
      RECT 27.435000  11.170000 47.380000  11.240000 ;
      RECT 27.435000  11.170000 47.380000  11.240000 ;
      RECT 27.505000  11.240000 47.310000  11.310000 ;
      RECT 27.505000  11.240000 47.310000  11.310000 ;
      RECT 27.575000  11.310000 47.240000  11.380000 ;
      RECT 27.575000  11.310000 47.240000  11.380000 ;
      RECT 27.645000  11.380000 47.170000  11.450000 ;
      RECT 27.645000  11.380000 47.170000  11.450000 ;
      RECT 27.715000  11.450000 47.100000  11.520000 ;
      RECT 27.715000  11.450000 47.100000  11.520000 ;
      RECT 27.785000  11.520000 47.030000  11.590000 ;
      RECT 27.785000  11.520000 47.030000  11.590000 ;
      RECT 27.855000  11.590000 46.960000  11.660000 ;
      RECT 27.855000  11.590000 46.960000  11.660000 ;
      RECT 27.925000  11.660000 46.890000  11.730000 ;
      RECT 27.925000  11.660000 46.890000  11.730000 ;
      RECT 27.995000  11.730000 46.820000  11.800000 ;
      RECT 27.995000  11.730000 46.820000  11.800000 ;
      RECT 28.035000   0.000000 50.250000   0.675000 ;
      RECT 28.065000  11.800000 46.750000  11.870000 ;
      RECT 28.065000  11.800000 46.750000  11.870000 ;
      RECT 28.135000  11.870000 46.680000  11.940000 ;
      RECT 28.135000  11.870000 46.680000  11.940000 ;
      RECT 28.175000   0.000000 50.110000   0.815000 ;
      RECT 28.175000   0.000000 50.110000   8.480000 ;
      RECT 28.205000  11.940000 46.610000  12.010000 ;
      RECT 28.205000  11.940000 46.610000  12.010000 ;
      RECT 28.210000  12.010000 46.605000  12.015000 ;
      RECT 28.210000  12.010000 46.605000  12.015000 ;
      RECT 28.260000  12.015000 37.610000  12.065000 ;
      RECT 28.260000  12.015000 37.610000  12.065000 ;
      RECT 28.310000  12.065000 37.610000  12.115000 ;
      RECT 28.310000  12.065000 37.610000  12.115000 ;
      RECT 28.315000  12.115000 37.610000  12.120000 ;
      RECT 28.315000  12.115000 37.610000  12.120000 ;
      RECT 37.175000  12.120000 37.610000  25.940000 ;
      RECT 37.175000  12.120000 46.660000  12.155000 ;
      RECT 37.175000  12.155000 37.750000  25.800000 ;
      RECT 37.175000  25.800000 55.935000  25.980000 ;
      RECT 37.175000  25.940000 55.700000  25.960000 ;
      RECT 37.175000  25.940000 55.700000  25.960000 ;
      RECT 37.175000  25.960000 55.720000  25.980000 ;
      RECT 37.175000  25.960000 55.720000  25.980000 ;
      RECT 54.325000  42.650000 60.830000  42.660000 ;
      RECT 54.325000  42.650000 60.830000  42.660000 ;
      RECT 54.395000  42.580000 60.830000  42.650000 ;
      RECT 54.395000  42.580000 60.830000  42.650000 ;
      RECT 54.465000  42.510000 60.830000  42.580000 ;
      RECT 54.465000  42.510000 60.830000  42.580000 ;
      RECT 54.535000  42.440000 60.830000  42.510000 ;
      RECT 54.535000  42.440000 60.830000  42.510000 ;
      RECT 54.605000  42.370000 60.830000  42.440000 ;
      RECT 54.605000  42.370000 60.830000  42.440000 ;
      RECT 54.675000  42.300000 60.830000  42.370000 ;
      RECT 54.675000  42.300000 60.830000  42.370000 ;
      RECT 54.745000  42.230000 60.830000  42.300000 ;
      RECT 54.745000  42.230000 60.830000  42.300000 ;
      RECT 54.815000  42.160000 60.830000  42.230000 ;
      RECT 54.815000  42.160000 60.830000  42.230000 ;
      RECT 54.885000  42.090000 60.830000  42.160000 ;
      RECT 54.885000  42.090000 60.830000  42.160000 ;
      RECT 54.955000  42.020000 60.830000  42.090000 ;
      RECT 54.955000  42.020000 60.830000  42.090000 ;
      RECT 55.025000  41.950000 60.830000  42.020000 ;
      RECT 55.025000  41.950000 60.830000  42.020000 ;
      RECT 55.095000  41.880000 60.830000  41.950000 ;
      RECT 55.095000  41.880000 60.830000  41.950000 ;
      RECT 55.165000  41.810000 60.830000  41.880000 ;
      RECT 55.165000  41.810000 60.830000  41.880000 ;
      RECT 55.235000  41.740000 60.830000  41.810000 ;
      RECT 55.235000  41.740000 60.830000  41.810000 ;
      RECT 55.305000  41.670000 60.830000  41.740000 ;
      RECT 55.305000  41.670000 60.830000  41.740000 ;
      RECT 55.375000  41.600000 60.830000  41.670000 ;
      RECT 55.375000  41.600000 60.830000  41.670000 ;
      RECT 55.445000  41.530000 60.830000  41.600000 ;
      RECT 55.445000  41.530000 60.830000  41.600000 ;
      RECT 55.515000  41.460000 60.830000  41.530000 ;
      RECT 55.515000  41.460000 60.830000  41.530000 ;
      RECT 55.585000  41.390000 60.830000  41.460000 ;
      RECT 55.585000  41.390000 60.830000  41.460000 ;
      RECT 55.655000  41.320000 60.830000  41.390000 ;
      RECT 55.655000  41.320000 60.830000  41.390000 ;
      RECT 55.725000  41.250000 60.830000  41.320000 ;
      RECT 55.725000  41.250000 60.830000  41.320000 ;
      RECT 55.795000  41.180000 60.830000  41.250000 ;
      RECT 55.795000  41.180000 60.830000  41.250000 ;
      RECT 55.865000  41.110000 60.830000  41.180000 ;
      RECT 55.865000  41.110000 60.830000  41.180000 ;
      RECT 55.935000  41.040000 60.830000  41.110000 ;
      RECT 55.935000  41.040000 60.830000  41.110000 ;
      RECT 56.005000  40.970000 60.830000  41.040000 ;
      RECT 56.005000  40.970000 60.830000  41.040000 ;
      RECT 56.075000  40.900000 60.830000  40.970000 ;
      RECT 56.075000  40.900000 60.830000  40.970000 ;
      RECT 56.145000  40.830000 60.830000  40.900000 ;
      RECT 56.145000  40.830000 60.830000  40.900000 ;
      RECT 56.215000  40.760000 60.830000  40.830000 ;
      RECT 56.215000  40.760000 60.830000  40.830000 ;
      RECT 56.285000  40.690000 60.830000  40.760000 ;
      RECT 56.285000  40.690000 60.830000  40.760000 ;
      RECT 56.355000  40.620000 60.830000  40.690000 ;
      RECT 56.355000  40.620000 60.830000  40.690000 ;
      RECT 56.425000  40.550000 60.830000  40.620000 ;
      RECT 56.425000  40.550000 60.830000  40.620000 ;
      RECT 56.495000  40.480000 60.830000  40.550000 ;
      RECT 56.495000  40.480000 60.830000  40.550000 ;
      RECT 56.565000  40.410000 60.830000  40.480000 ;
      RECT 56.565000  40.410000 60.830000  40.480000 ;
      RECT 56.635000  40.340000 60.830000  40.410000 ;
      RECT 56.635000  40.340000 60.830000  40.410000 ;
      RECT 56.705000  40.270000 60.830000  40.340000 ;
      RECT 56.705000  40.270000 60.830000  40.340000 ;
      RECT 56.775000  40.200000 60.830000  40.270000 ;
      RECT 56.775000  40.200000 60.830000  40.270000 ;
      RECT 56.845000  40.130000 60.830000  40.200000 ;
      RECT 56.845000  40.130000 60.830000  40.200000 ;
      RECT 56.915000  40.060000 60.830000  40.130000 ;
      RECT 56.915000  40.060000 60.830000  40.130000 ;
      RECT 56.985000  39.990000 60.830000  40.060000 ;
      RECT 56.985000  39.990000 60.830000  40.060000 ;
      RECT 56.985000  79.435000 57.440000  79.505000 ;
      RECT 56.985000  79.435000 57.440000  79.505000 ;
      RECT 56.985000  79.505000 57.510000  79.575000 ;
      RECT 56.985000  79.505000 57.510000  79.575000 ;
      RECT 56.985000  79.575000 57.580000  79.645000 ;
      RECT 56.985000  79.575000 57.580000  79.645000 ;
      RECT 56.985000  79.645000 57.650000  79.715000 ;
      RECT 56.985000  79.645000 57.650000  79.715000 ;
      RECT 56.985000  79.715000 57.720000  79.785000 ;
      RECT 56.985000  79.715000 57.720000  79.785000 ;
      RECT 56.985000  79.785000 57.790000  79.855000 ;
      RECT 56.985000  79.785000 57.790000  79.855000 ;
      RECT 56.985000  79.855000 57.860000  79.925000 ;
      RECT 56.985000  79.855000 57.860000  79.925000 ;
      RECT 56.985000  79.925000 57.930000  79.995000 ;
      RECT 56.985000  79.925000 57.930000  79.995000 ;
      RECT 56.985000  79.995000 58.000000  80.065000 ;
      RECT 56.985000  79.995000 58.000000  80.065000 ;
      RECT 56.985000  80.065000 58.070000  80.135000 ;
      RECT 56.985000  80.065000 58.070000  80.135000 ;
      RECT 56.985000  80.135000 58.140000  80.205000 ;
      RECT 56.985000  80.135000 58.140000  80.205000 ;
      RECT 56.985000  80.205000 58.210000  80.275000 ;
      RECT 56.985000  80.205000 58.210000  80.275000 ;
      RECT 56.985000  80.275000 58.280000  80.345000 ;
      RECT 56.985000  80.275000 58.280000  80.345000 ;
      RECT 56.985000  80.345000 58.350000  80.415000 ;
      RECT 56.985000  80.345000 58.350000  80.415000 ;
      RECT 56.985000  80.415000 58.420000  80.485000 ;
      RECT 56.985000  80.415000 58.420000  80.485000 ;
      RECT 56.985000  80.485000 58.490000  80.500000 ;
      RECT 56.985000  80.485000 58.490000  80.500000 ;
      RECT 56.985000  80.500000 58.505000  80.570000 ;
      RECT 56.985000  80.500000 58.505000  80.570000 ;
      RECT 56.985000  80.500000 60.970000  82.770000 ;
      RECT 56.985000  80.570000 58.575000  80.640000 ;
      RECT 56.985000  80.570000 58.575000  80.640000 ;
      RECT 56.985000  80.640000 58.645000  80.710000 ;
      RECT 56.985000  80.640000 58.645000  80.710000 ;
      RECT 56.985000  80.710000 58.715000  80.780000 ;
      RECT 56.985000  80.710000 58.715000  80.780000 ;
      RECT 56.985000  80.780000 58.785000  80.850000 ;
      RECT 56.985000  80.780000 58.785000  80.850000 ;
      RECT 56.985000  80.850000 58.855000  80.920000 ;
      RECT 56.985000  80.850000 58.855000  80.920000 ;
      RECT 56.985000  80.920000 58.925000  80.990000 ;
      RECT 56.985000  80.920000 58.925000  80.990000 ;
      RECT 56.985000  80.990000 58.995000  81.060000 ;
      RECT 56.985000  80.990000 58.995000  81.060000 ;
      RECT 56.985000  81.060000 59.065000  81.130000 ;
      RECT 56.985000  81.060000 59.065000  81.130000 ;
      RECT 56.985000  81.130000 59.135000  81.200000 ;
      RECT 56.985000  81.130000 59.135000  81.200000 ;
      RECT 56.985000  81.200000 59.205000  81.270000 ;
      RECT 56.985000  81.200000 59.205000  81.270000 ;
      RECT 56.985000  81.270000 59.275000  81.340000 ;
      RECT 56.985000  81.270000 59.275000  81.340000 ;
      RECT 56.985000  81.340000 59.345000  81.410000 ;
      RECT 56.985000  81.340000 59.345000  81.410000 ;
      RECT 56.985000  81.410000 59.415000  81.480000 ;
      RECT 56.985000  81.410000 59.415000  81.480000 ;
      RECT 56.985000  81.480000 59.485000  81.550000 ;
      RECT 56.985000  81.480000 59.485000  81.550000 ;
      RECT 56.985000  81.550000 59.555000  81.620000 ;
      RECT 56.985000  81.550000 59.555000  81.620000 ;
      RECT 56.985000  81.620000 59.625000  81.690000 ;
      RECT 56.985000  81.620000 59.625000  81.690000 ;
      RECT 56.985000  81.690000 59.695000  81.760000 ;
      RECT 56.985000  81.690000 59.695000  81.760000 ;
      RECT 56.985000  81.760000 59.765000  81.830000 ;
      RECT 56.985000  81.760000 59.765000  81.830000 ;
      RECT 56.985000  81.830000 59.835000  81.900000 ;
      RECT 56.985000  81.830000 59.835000  81.900000 ;
      RECT 56.985000  81.900000 59.905000  81.970000 ;
      RECT 56.985000  81.900000 59.905000  81.970000 ;
      RECT 56.985000  81.970000 59.975000  82.040000 ;
      RECT 56.985000  81.970000 59.975000  82.040000 ;
      RECT 56.985000  82.040000 60.045000  82.110000 ;
      RECT 56.985000  82.040000 60.045000  82.110000 ;
      RECT 56.985000  82.110000 60.115000  82.180000 ;
      RECT 56.985000  82.110000 60.115000  82.180000 ;
      RECT 56.985000  82.180000 60.185000  82.250000 ;
      RECT 56.985000  82.180000 60.185000  82.250000 ;
      RECT 56.985000  82.250000 60.255000  82.320000 ;
      RECT 56.985000  82.250000 60.255000  82.320000 ;
      RECT 56.985000  82.320000 60.325000  82.390000 ;
      RECT 56.985000  82.320000 60.325000  82.390000 ;
      RECT 56.985000  82.390000 60.395000  82.460000 ;
      RECT 56.985000  82.390000 60.395000  82.460000 ;
      RECT 56.985000  82.460000 60.465000  82.530000 ;
      RECT 56.985000  82.460000 60.465000  82.530000 ;
      RECT 56.985000  82.530000 60.535000  82.600000 ;
      RECT 56.985000  82.530000 60.535000  82.600000 ;
      RECT 56.985000  82.600000 60.605000  82.670000 ;
      RECT 56.985000  82.600000 60.605000  82.670000 ;
      RECT 56.985000  82.670000 60.675000  82.740000 ;
      RECT 56.985000  82.670000 60.675000  82.740000 ;
      RECT 56.985000  82.740000 60.745000  82.810000 ;
      RECT 56.985000  82.740000 60.745000  82.810000 ;
      RECT 56.985000  82.770000 60.970000  89.760000 ;
      RECT 56.985000  82.810000 60.815000  82.825000 ;
      RECT 56.985000  82.810000 60.815000  82.825000 ;
      RECT 56.985000  82.825000 60.830000  89.760000 ;
      RECT 56.985000 102.435000 57.440000 102.505000 ;
      RECT 56.985000 102.435000 57.440000 102.505000 ;
      RECT 56.985000 102.505000 57.510000 102.575000 ;
      RECT 56.985000 102.505000 57.510000 102.575000 ;
      RECT 56.985000 102.575000 57.580000 102.645000 ;
      RECT 56.985000 102.575000 57.580000 102.645000 ;
      RECT 56.985000 102.645000 57.650000 102.715000 ;
      RECT 56.985000 102.645000 57.650000 102.715000 ;
      RECT 56.985000 102.715000 57.720000 102.785000 ;
      RECT 56.985000 102.715000 57.720000 102.785000 ;
      RECT 56.985000 102.785000 57.790000 102.855000 ;
      RECT 56.985000 102.785000 57.790000 102.855000 ;
      RECT 56.985000 102.855000 57.860000 102.925000 ;
      RECT 56.985000 102.855000 57.860000 102.925000 ;
      RECT 56.985000 102.925000 57.930000 102.995000 ;
      RECT 56.985000 102.925000 57.930000 102.995000 ;
      RECT 56.985000 102.995000 58.000000 103.065000 ;
      RECT 56.985000 102.995000 58.000000 103.065000 ;
      RECT 56.985000 103.065000 58.070000 103.135000 ;
      RECT 56.985000 103.065000 58.070000 103.135000 ;
      RECT 56.985000 103.135000 58.140000 103.205000 ;
      RECT 56.985000 103.135000 58.140000 103.205000 ;
      RECT 56.985000 103.205000 58.210000 103.275000 ;
      RECT 56.985000 103.205000 58.210000 103.275000 ;
      RECT 56.985000 103.275000 58.280000 103.345000 ;
      RECT 56.985000 103.275000 58.280000 103.345000 ;
      RECT 56.985000 103.345000 58.350000 103.415000 ;
      RECT 56.985000 103.345000 58.350000 103.415000 ;
      RECT 56.985000 103.415000 58.420000 103.485000 ;
      RECT 56.985000 103.415000 58.420000 103.485000 ;
      RECT 56.985000 103.485000 58.490000 103.500000 ;
      RECT 56.985000 103.485000 58.490000 103.500000 ;
      RECT 56.985000 103.500000 58.505000 103.570000 ;
      RECT 56.985000 103.500000 58.505000 103.570000 ;
      RECT 56.985000 103.500000 60.970000 105.770000 ;
      RECT 56.985000 103.570000 58.575000 103.640000 ;
      RECT 56.985000 103.570000 58.575000 103.640000 ;
      RECT 56.985000 103.640000 58.645000 103.710000 ;
      RECT 56.985000 103.640000 58.645000 103.710000 ;
      RECT 56.985000 103.710000 58.715000 103.780000 ;
      RECT 56.985000 103.710000 58.715000 103.780000 ;
      RECT 56.985000 103.780000 58.785000 103.850000 ;
      RECT 56.985000 103.780000 58.785000 103.850000 ;
      RECT 56.985000 103.850000 58.855000 103.920000 ;
      RECT 56.985000 103.850000 58.855000 103.920000 ;
      RECT 56.985000 103.920000 58.925000 103.990000 ;
      RECT 56.985000 103.920000 58.925000 103.990000 ;
      RECT 56.985000 103.990000 58.995000 104.060000 ;
      RECT 56.985000 103.990000 58.995000 104.060000 ;
      RECT 56.985000 104.060000 59.065000 104.130000 ;
      RECT 56.985000 104.060000 59.065000 104.130000 ;
      RECT 56.985000 104.130000 59.135000 104.200000 ;
      RECT 56.985000 104.130000 59.135000 104.200000 ;
      RECT 56.985000 104.200000 59.205000 104.270000 ;
      RECT 56.985000 104.200000 59.205000 104.270000 ;
      RECT 56.985000 104.270000 59.275000 104.340000 ;
      RECT 56.985000 104.270000 59.275000 104.340000 ;
      RECT 56.985000 104.340000 59.345000 104.410000 ;
      RECT 56.985000 104.340000 59.345000 104.410000 ;
      RECT 56.985000 104.410000 59.415000 104.480000 ;
      RECT 56.985000 104.410000 59.415000 104.480000 ;
      RECT 56.985000 104.480000 59.485000 104.550000 ;
      RECT 56.985000 104.480000 59.485000 104.550000 ;
      RECT 56.985000 104.550000 59.555000 104.620000 ;
      RECT 56.985000 104.550000 59.555000 104.620000 ;
      RECT 56.985000 104.620000 59.625000 104.690000 ;
      RECT 56.985000 104.620000 59.625000 104.690000 ;
      RECT 56.985000 104.690000 59.695000 104.760000 ;
      RECT 56.985000 104.690000 59.695000 104.760000 ;
      RECT 56.985000 104.760000 59.765000 104.830000 ;
      RECT 56.985000 104.760000 59.765000 104.830000 ;
      RECT 56.985000 104.830000 59.835000 104.900000 ;
      RECT 56.985000 104.830000 59.835000 104.900000 ;
      RECT 56.985000 104.900000 59.905000 104.970000 ;
      RECT 56.985000 104.900000 59.905000 104.970000 ;
      RECT 56.985000 104.970000 59.975000 105.040000 ;
      RECT 56.985000 104.970000 59.975000 105.040000 ;
      RECT 56.985000 105.040000 60.045000 105.110000 ;
      RECT 56.985000 105.040000 60.045000 105.110000 ;
      RECT 56.985000 105.110000 60.115000 105.180000 ;
      RECT 56.985000 105.110000 60.115000 105.180000 ;
      RECT 56.985000 105.180000 60.185000 105.250000 ;
      RECT 56.985000 105.180000 60.185000 105.250000 ;
      RECT 56.985000 105.250000 60.255000 105.320000 ;
      RECT 56.985000 105.250000 60.255000 105.320000 ;
      RECT 56.985000 105.320000 60.325000 105.390000 ;
      RECT 56.985000 105.320000 60.325000 105.390000 ;
      RECT 56.985000 105.390000 60.395000 105.460000 ;
      RECT 56.985000 105.390000 60.395000 105.460000 ;
      RECT 56.985000 105.460000 60.465000 105.530000 ;
      RECT 56.985000 105.460000 60.465000 105.530000 ;
      RECT 56.985000 105.530000 60.535000 105.600000 ;
      RECT 56.985000 105.530000 60.535000 105.600000 ;
      RECT 56.985000 105.600000 60.605000 105.670000 ;
      RECT 56.985000 105.600000 60.605000 105.670000 ;
      RECT 56.985000 105.670000 60.675000 105.740000 ;
      RECT 56.985000 105.670000 60.675000 105.740000 ;
      RECT 56.985000 105.740000 60.745000 105.810000 ;
      RECT 56.985000 105.740000 60.745000 105.810000 ;
      RECT 56.985000 105.770000 60.970000 112.760000 ;
      RECT 56.985000 105.810000 60.815000 105.825000 ;
      RECT 56.985000 105.810000 60.815000 105.825000 ;
      RECT 56.985000 105.825000 60.830000 112.705000 ;
      RECT 56.985000 112.705000 60.805000 112.730000 ;
      RECT 56.985000 112.705000 60.805000 112.730000 ;
      RECT 56.985000 112.730000 60.775000 112.760000 ;
      RECT 56.985000 112.730000 60.775000 112.760000 ;
      RECT 56.985000 125.435000 57.440000 125.505000 ;
      RECT 56.985000 125.435000 57.440000 125.505000 ;
      RECT 56.985000 125.505000 57.510000 125.575000 ;
      RECT 56.985000 125.505000 57.510000 125.575000 ;
      RECT 56.985000 125.575000 57.580000 125.645000 ;
      RECT 56.985000 125.575000 57.580000 125.645000 ;
      RECT 56.985000 125.645000 57.650000 125.715000 ;
      RECT 56.985000 125.645000 57.650000 125.715000 ;
      RECT 56.985000 125.715000 57.720000 125.785000 ;
      RECT 56.985000 125.715000 57.720000 125.785000 ;
      RECT 56.985000 125.785000 57.790000 125.855000 ;
      RECT 56.985000 125.785000 57.790000 125.855000 ;
      RECT 56.985000 125.855000 57.860000 125.925000 ;
      RECT 56.985000 125.855000 57.860000 125.925000 ;
      RECT 56.985000 125.925000 57.930000 125.995000 ;
      RECT 56.985000 125.925000 57.930000 125.995000 ;
      RECT 56.985000 125.995000 58.000000 126.065000 ;
      RECT 56.985000 125.995000 58.000000 126.065000 ;
      RECT 56.985000 126.065000 58.070000 126.135000 ;
      RECT 56.985000 126.065000 58.070000 126.135000 ;
      RECT 56.985000 126.135000 58.140000 126.205000 ;
      RECT 56.985000 126.135000 58.140000 126.205000 ;
      RECT 56.985000 126.205000 58.210000 126.275000 ;
      RECT 56.985000 126.205000 58.210000 126.275000 ;
      RECT 56.985000 126.275000 58.280000 126.345000 ;
      RECT 56.985000 126.275000 58.280000 126.345000 ;
      RECT 56.985000 126.345000 58.350000 126.415000 ;
      RECT 56.985000 126.345000 58.350000 126.415000 ;
      RECT 56.985000 126.415000 58.420000 126.485000 ;
      RECT 56.985000 126.415000 58.420000 126.485000 ;
      RECT 56.985000 126.485000 58.490000 126.500000 ;
      RECT 56.985000 126.485000 58.490000 126.500000 ;
      RECT 56.985000 126.500000 58.505000 126.570000 ;
      RECT 56.985000 126.500000 58.505000 126.570000 ;
      RECT 56.985000 126.500000 60.970000 128.770000 ;
      RECT 56.985000 126.570000 58.575000 126.640000 ;
      RECT 56.985000 126.570000 58.575000 126.640000 ;
      RECT 56.985000 126.640000 58.645000 126.710000 ;
      RECT 56.985000 126.640000 58.645000 126.710000 ;
      RECT 56.985000 126.710000 58.715000 126.780000 ;
      RECT 56.985000 126.710000 58.715000 126.780000 ;
      RECT 56.985000 126.780000 58.785000 126.850000 ;
      RECT 56.985000 126.780000 58.785000 126.850000 ;
      RECT 56.985000 126.850000 58.855000 126.920000 ;
      RECT 56.985000 126.850000 58.855000 126.920000 ;
      RECT 56.985000 126.920000 58.925000 126.990000 ;
      RECT 56.985000 126.920000 58.925000 126.990000 ;
      RECT 56.985000 126.990000 58.995000 127.060000 ;
      RECT 56.985000 126.990000 58.995000 127.060000 ;
      RECT 56.985000 127.060000 59.065000 127.130000 ;
      RECT 56.985000 127.060000 59.065000 127.130000 ;
      RECT 56.985000 127.130000 59.135000 127.200000 ;
      RECT 56.985000 127.130000 59.135000 127.200000 ;
      RECT 56.985000 127.200000 59.205000 127.270000 ;
      RECT 56.985000 127.200000 59.205000 127.270000 ;
      RECT 56.985000 127.270000 59.275000 127.340000 ;
      RECT 56.985000 127.270000 59.275000 127.340000 ;
      RECT 56.985000 127.340000 59.345000 127.410000 ;
      RECT 56.985000 127.340000 59.345000 127.410000 ;
      RECT 56.985000 127.410000 59.415000 127.480000 ;
      RECT 56.985000 127.410000 59.415000 127.480000 ;
      RECT 56.985000 127.480000 59.485000 127.550000 ;
      RECT 56.985000 127.480000 59.485000 127.550000 ;
      RECT 56.985000 127.550000 59.555000 127.620000 ;
      RECT 56.985000 127.550000 59.555000 127.620000 ;
      RECT 56.985000 127.620000 59.625000 127.690000 ;
      RECT 56.985000 127.620000 59.625000 127.690000 ;
      RECT 56.985000 127.690000 59.695000 127.760000 ;
      RECT 56.985000 127.690000 59.695000 127.760000 ;
      RECT 56.985000 127.760000 59.765000 127.830000 ;
      RECT 56.985000 127.760000 59.765000 127.830000 ;
      RECT 56.985000 127.830000 59.835000 127.900000 ;
      RECT 56.985000 127.830000 59.835000 127.900000 ;
      RECT 56.985000 127.900000 59.905000 127.970000 ;
      RECT 56.985000 127.900000 59.905000 127.970000 ;
      RECT 56.985000 127.970000 59.975000 128.040000 ;
      RECT 56.985000 127.970000 59.975000 128.040000 ;
      RECT 56.985000 128.040000 60.045000 128.110000 ;
      RECT 56.985000 128.040000 60.045000 128.110000 ;
      RECT 56.985000 128.110000 60.115000 128.180000 ;
      RECT 56.985000 128.110000 60.115000 128.180000 ;
      RECT 56.985000 128.180000 60.185000 128.250000 ;
      RECT 56.985000 128.180000 60.185000 128.250000 ;
      RECT 56.985000 128.250000 60.255000 128.320000 ;
      RECT 56.985000 128.250000 60.255000 128.320000 ;
      RECT 56.985000 128.320000 60.325000 128.390000 ;
      RECT 56.985000 128.320000 60.325000 128.390000 ;
      RECT 56.985000 128.390000 60.395000 128.460000 ;
      RECT 56.985000 128.390000 60.395000 128.460000 ;
      RECT 56.985000 128.460000 60.465000 128.530000 ;
      RECT 56.985000 128.460000 60.465000 128.530000 ;
      RECT 56.985000 128.530000 60.535000 128.600000 ;
      RECT 56.985000 128.530000 60.535000 128.600000 ;
      RECT 56.985000 128.600000 60.605000 128.670000 ;
      RECT 56.985000 128.600000 60.605000 128.670000 ;
      RECT 56.985000 128.670000 60.675000 128.740000 ;
      RECT 56.985000 128.670000 60.675000 128.740000 ;
      RECT 56.985000 128.740000 60.745000 128.810000 ;
      RECT 56.985000 128.740000 60.745000 128.810000 ;
      RECT 56.985000 128.770000 60.970000 135.760000 ;
      RECT 56.985000 128.810000 60.815000 128.825000 ;
      RECT 56.985000 128.810000 60.815000 128.825000 ;
      RECT 56.985000 128.825000 60.830000 135.740000 ;
      RECT 56.985000 135.740000 60.820000 135.750000 ;
      RECT 56.985000 135.740000 60.820000 135.750000 ;
      RECT 56.985000 135.750000 60.810000 135.760000 ;
      RECT 56.985000 135.750000 60.810000 135.760000 ;
      RECT 56.985000 148.435000 57.370000 148.505000 ;
      RECT 56.985000 148.435000 57.370000 148.505000 ;
      RECT 56.985000 148.505000 57.440000 148.575000 ;
      RECT 56.985000 148.505000 57.440000 148.575000 ;
      RECT 56.985000 148.575000 57.510000 148.645000 ;
      RECT 56.985000 148.575000 57.510000 148.645000 ;
      RECT 56.985000 148.645000 57.580000 148.715000 ;
      RECT 56.985000 148.645000 57.580000 148.715000 ;
      RECT 56.985000 148.715000 57.650000 148.785000 ;
      RECT 56.985000 148.715000 57.650000 148.785000 ;
      RECT 56.985000 148.785000 57.720000 148.855000 ;
      RECT 56.985000 148.785000 57.720000 148.855000 ;
      RECT 56.985000 148.855000 57.790000 148.925000 ;
      RECT 56.985000 148.855000 57.790000 148.925000 ;
      RECT 56.985000 148.925000 57.860000 148.995000 ;
      RECT 56.985000 148.925000 57.860000 148.995000 ;
      RECT 56.985000 148.995000 57.930000 149.065000 ;
      RECT 56.985000 148.995000 57.930000 149.065000 ;
      RECT 56.985000 149.065000 58.000000 149.135000 ;
      RECT 56.985000 149.065000 58.000000 149.135000 ;
      RECT 56.985000 149.135000 58.070000 149.205000 ;
      RECT 56.985000 149.135000 58.070000 149.205000 ;
      RECT 56.985000 149.205000 58.140000 149.275000 ;
      RECT 56.985000 149.205000 58.140000 149.275000 ;
      RECT 56.985000 149.275000 58.210000 149.345000 ;
      RECT 56.985000 149.275000 58.210000 149.345000 ;
      RECT 56.985000 149.345000 58.280000 149.415000 ;
      RECT 56.985000 149.345000 58.280000 149.415000 ;
      RECT 56.985000 149.415000 58.350000 149.485000 ;
      RECT 56.985000 149.415000 58.350000 149.485000 ;
      RECT 56.985000 149.485000 58.420000 149.500000 ;
      RECT 56.985000 149.485000 58.420000 149.500000 ;
      RECT 56.985000 149.500000 58.435000 149.570000 ;
      RECT 56.985000 149.500000 58.435000 149.570000 ;
      RECT 56.985000 149.500000 60.970000 151.840000 ;
      RECT 56.985000 149.570000 58.505000 149.640000 ;
      RECT 56.985000 149.570000 58.505000 149.640000 ;
      RECT 56.985000 149.640000 58.575000 149.710000 ;
      RECT 56.985000 149.640000 58.575000 149.710000 ;
      RECT 56.985000 149.710000 58.645000 149.780000 ;
      RECT 56.985000 149.710000 58.645000 149.780000 ;
      RECT 56.985000 149.780000 58.715000 149.850000 ;
      RECT 56.985000 149.780000 58.715000 149.850000 ;
      RECT 56.985000 149.850000 58.785000 149.920000 ;
      RECT 56.985000 149.850000 58.785000 149.920000 ;
      RECT 56.985000 149.920000 58.855000 149.990000 ;
      RECT 56.985000 149.920000 58.855000 149.990000 ;
      RECT 56.985000 149.990000 58.925000 150.060000 ;
      RECT 56.985000 149.990000 58.925000 150.060000 ;
      RECT 56.985000 150.060000 58.995000 150.130000 ;
      RECT 56.985000 150.060000 58.995000 150.130000 ;
      RECT 56.985000 150.130000 59.065000 150.200000 ;
      RECT 56.985000 150.130000 59.065000 150.200000 ;
      RECT 56.985000 150.200000 59.135000 150.270000 ;
      RECT 56.985000 150.200000 59.135000 150.270000 ;
      RECT 56.985000 150.270000 59.205000 150.340000 ;
      RECT 56.985000 150.270000 59.205000 150.340000 ;
      RECT 56.985000 150.340000 59.275000 150.410000 ;
      RECT 56.985000 150.340000 59.275000 150.410000 ;
      RECT 56.985000 150.410000 59.345000 150.480000 ;
      RECT 56.985000 150.410000 59.345000 150.480000 ;
      RECT 56.985000 150.480000 59.415000 150.550000 ;
      RECT 56.985000 150.480000 59.415000 150.550000 ;
      RECT 56.985000 150.550000 59.485000 150.620000 ;
      RECT 56.985000 150.550000 59.485000 150.620000 ;
      RECT 56.985000 150.620000 59.555000 150.690000 ;
      RECT 56.985000 150.620000 59.555000 150.690000 ;
      RECT 56.985000 150.690000 59.625000 150.760000 ;
      RECT 56.985000 150.690000 59.625000 150.760000 ;
      RECT 56.985000 150.760000 59.695000 150.830000 ;
      RECT 56.985000 150.760000 59.695000 150.830000 ;
      RECT 56.985000 150.830000 59.765000 150.900000 ;
      RECT 56.985000 150.830000 59.765000 150.900000 ;
      RECT 56.985000 150.900000 59.835000 150.970000 ;
      RECT 56.985000 150.900000 59.835000 150.970000 ;
      RECT 56.985000 150.970000 59.905000 151.040000 ;
      RECT 56.985000 150.970000 59.905000 151.040000 ;
      RECT 56.985000 151.040000 59.975000 151.110000 ;
      RECT 56.985000 151.040000 59.975000 151.110000 ;
      RECT 56.985000 151.110000 60.045000 151.180000 ;
      RECT 56.985000 151.110000 60.045000 151.180000 ;
      RECT 56.985000 151.180000 60.115000 151.250000 ;
      RECT 56.985000 151.180000 60.115000 151.250000 ;
      RECT 56.985000 151.250000 60.185000 151.320000 ;
      RECT 56.985000 151.250000 60.185000 151.320000 ;
      RECT 56.985000 151.320000 60.255000 151.390000 ;
      RECT 56.985000 151.320000 60.255000 151.390000 ;
      RECT 56.985000 151.390000 60.325000 151.460000 ;
      RECT 56.985000 151.390000 60.325000 151.460000 ;
      RECT 56.985000 151.460000 60.395000 151.530000 ;
      RECT 56.985000 151.460000 60.395000 151.530000 ;
      RECT 56.985000 151.530000 60.465000 151.600000 ;
      RECT 56.985000 151.530000 60.465000 151.600000 ;
      RECT 56.985000 151.600000 60.535000 151.670000 ;
      RECT 56.985000 151.600000 60.535000 151.670000 ;
      RECT 56.985000 151.670000 60.605000 151.740000 ;
      RECT 56.985000 151.670000 60.605000 151.740000 ;
      RECT 56.985000 151.740000 60.675000 151.810000 ;
      RECT 56.985000 151.740000 60.675000 151.810000 ;
      RECT 56.985000 151.810000 60.745000 151.880000 ;
      RECT 56.985000 151.810000 60.745000 151.880000 ;
      RECT 56.985000 151.840000 60.970000 158.760000 ;
      RECT 56.985000 151.880000 60.815000 151.895000 ;
      RECT 56.985000 151.880000 60.815000 151.895000 ;
      RECT 56.985000 151.895000 60.830000 158.755000 ;
      RECT 56.985000 158.755000 60.825000 158.760000 ;
      RECT 56.985000 158.755000 60.825000 158.760000 ;
      RECT 56.990000  56.435000 57.410000  56.505000 ;
      RECT 56.990000  56.435000 57.410000  56.505000 ;
      RECT 56.990000  56.505000 57.480000  56.575000 ;
      RECT 56.990000  56.505000 57.480000  56.575000 ;
      RECT 56.990000  56.575000 57.550000  56.645000 ;
      RECT 56.990000  56.575000 57.550000  56.645000 ;
      RECT 56.990000  56.645000 57.620000  56.715000 ;
      RECT 56.990000  56.645000 57.620000  56.715000 ;
      RECT 56.990000  56.715000 57.690000  56.785000 ;
      RECT 56.990000  56.715000 57.690000  56.785000 ;
      RECT 56.990000  56.785000 57.760000  56.855000 ;
      RECT 56.990000  56.785000 57.760000  56.855000 ;
      RECT 56.990000  56.855000 57.830000  56.925000 ;
      RECT 56.990000  56.855000 57.830000  56.925000 ;
      RECT 56.990000  56.925000 57.900000  56.995000 ;
      RECT 56.990000  56.925000 57.900000  56.995000 ;
      RECT 56.990000  56.995000 57.970000  57.065000 ;
      RECT 56.990000  56.995000 57.970000  57.065000 ;
      RECT 56.990000  57.065000 58.040000  57.135000 ;
      RECT 56.990000  57.065000 58.040000  57.135000 ;
      RECT 56.990000  57.135000 58.110000  57.205000 ;
      RECT 56.990000  57.135000 58.110000  57.205000 ;
      RECT 56.990000  57.205000 58.180000  57.275000 ;
      RECT 56.990000  57.205000 58.180000  57.275000 ;
      RECT 56.990000  57.275000 58.250000  57.345000 ;
      RECT 56.990000  57.275000 58.250000  57.345000 ;
      RECT 56.990000  57.345000 58.320000  57.415000 ;
      RECT 56.990000  57.345000 58.320000  57.415000 ;
      RECT 56.990000  57.415000 58.390000  57.485000 ;
      RECT 56.990000  57.415000 58.390000  57.485000 ;
      RECT 56.990000  57.485000 58.460000  57.500000 ;
      RECT 56.990000  57.485000 58.460000  57.500000 ;
      RECT 56.990000  57.500000 58.475000  57.570000 ;
      RECT 56.990000  57.500000 58.475000  57.570000 ;
      RECT 56.990000  57.500000 60.970000  59.800000 ;
      RECT 56.990000  57.570000 58.545000  57.640000 ;
      RECT 56.990000  57.570000 58.545000  57.640000 ;
      RECT 56.990000  57.640000 58.615000  57.710000 ;
      RECT 56.990000  57.640000 58.615000  57.710000 ;
      RECT 56.990000  57.710000 58.685000  57.780000 ;
      RECT 56.990000  57.710000 58.685000  57.780000 ;
      RECT 56.990000  57.780000 58.755000  57.850000 ;
      RECT 56.990000  57.780000 58.755000  57.850000 ;
      RECT 56.990000  57.850000 58.825000  57.920000 ;
      RECT 56.990000  57.850000 58.825000  57.920000 ;
      RECT 56.990000  57.920000 58.895000  57.990000 ;
      RECT 56.990000  57.920000 58.895000  57.990000 ;
      RECT 56.990000  57.990000 58.965000  58.060000 ;
      RECT 56.990000  57.990000 58.965000  58.060000 ;
      RECT 56.990000  58.060000 59.035000  58.130000 ;
      RECT 56.990000  58.060000 59.035000  58.130000 ;
      RECT 56.990000  58.130000 59.105000  58.200000 ;
      RECT 56.990000  58.130000 59.105000  58.200000 ;
      RECT 56.990000  58.200000 59.175000  58.270000 ;
      RECT 56.990000  58.200000 59.175000  58.270000 ;
      RECT 56.990000  58.270000 59.245000  58.340000 ;
      RECT 56.990000  58.270000 59.245000  58.340000 ;
      RECT 56.990000  58.340000 59.315000  58.410000 ;
      RECT 56.990000  58.340000 59.315000  58.410000 ;
      RECT 56.990000  58.410000 59.385000  58.480000 ;
      RECT 56.990000  58.410000 59.385000  58.480000 ;
      RECT 56.990000  58.480000 59.455000  58.550000 ;
      RECT 56.990000  58.480000 59.455000  58.550000 ;
      RECT 56.990000  58.550000 59.525000  58.620000 ;
      RECT 56.990000  58.550000 59.525000  58.620000 ;
      RECT 56.990000  58.620000 59.595000  58.690000 ;
      RECT 56.990000  58.620000 59.595000  58.690000 ;
      RECT 56.990000  58.690000 59.665000  58.760000 ;
      RECT 56.990000  58.690000 59.665000  58.760000 ;
      RECT 56.990000  58.760000 59.735000  58.830000 ;
      RECT 56.990000  58.760000 59.735000  58.830000 ;
      RECT 56.990000  58.830000 59.805000  58.900000 ;
      RECT 56.990000  58.830000 59.805000  58.900000 ;
      RECT 56.990000  58.900000 59.875000  58.970000 ;
      RECT 56.990000  58.900000 59.875000  58.970000 ;
      RECT 56.990000  58.970000 59.945000  59.040000 ;
      RECT 56.990000  58.970000 59.945000  59.040000 ;
      RECT 56.990000  59.040000 60.015000  59.110000 ;
      RECT 56.990000  59.040000 60.015000  59.110000 ;
      RECT 56.990000  59.110000 60.085000  59.180000 ;
      RECT 56.990000  59.110000 60.085000  59.180000 ;
      RECT 56.990000  59.180000 60.155000  59.250000 ;
      RECT 56.990000  59.180000 60.155000  59.250000 ;
      RECT 56.990000  59.250000 60.225000  59.320000 ;
      RECT 56.990000  59.250000 60.225000  59.320000 ;
      RECT 56.990000  59.320000 60.295000  59.390000 ;
      RECT 56.990000  59.320000 60.295000  59.390000 ;
      RECT 56.990000  59.390000 60.365000  59.460000 ;
      RECT 56.990000  59.390000 60.365000  59.460000 ;
      RECT 56.990000  59.460000 60.435000  59.530000 ;
      RECT 56.990000  59.460000 60.435000  59.530000 ;
      RECT 56.990000  59.530000 60.505000  59.600000 ;
      RECT 56.990000  59.530000 60.505000  59.600000 ;
      RECT 56.990000  59.600000 60.575000  59.670000 ;
      RECT 56.990000  59.600000 60.575000  59.670000 ;
      RECT 56.990000  59.670000 60.645000  59.740000 ;
      RECT 56.990000  59.670000 60.645000  59.740000 ;
      RECT 56.990000  59.740000 60.715000  59.810000 ;
      RECT 56.990000  59.740000 60.715000  59.810000 ;
      RECT 56.990000  59.800000 60.970000  66.760000 ;
      RECT 56.990000  59.810000 60.785000  59.855000 ;
      RECT 56.990000  59.810000 60.785000  59.855000 ;
      RECT 56.990000  59.855000 60.830000  66.735000 ;
      RECT 56.990000  66.735000 60.820000  66.745000 ;
      RECT 56.990000  66.735000 60.820000  66.745000 ;
      RECT 56.990000  66.745000 60.805000  66.760000 ;
      RECT 56.990000  66.745000 60.805000  66.760000 ;
      RECT 57.055000  35.975000 60.970000  39.725000 ;
      RECT 57.055000  39.725000 60.970000  42.520000 ;
      RECT 57.055000  39.920000 60.830000  39.990000 ;
      RECT 57.055000  39.920000 60.830000  39.990000 ;
      RECT 57.125000  39.850000 60.830000  39.920000 ;
      RECT 57.125000  39.850000 60.830000  39.920000 ;
      RECT 57.195000  35.835000 60.830000  39.780000 ;
      RECT 57.195000  39.780000 60.830000  39.850000 ;
      RECT 57.195000  39.780000 60.830000  39.850000 ;
      RECT 58.240000 172.500000 58.515000 172.570000 ;
      RECT 58.240000 172.500000 60.970000 174.760000 ;
      RECT 58.240000 172.570000 58.585000 172.640000 ;
      RECT 58.240000 172.640000 58.655000 172.710000 ;
      RECT 58.240000 172.710000 58.725000 172.780000 ;
      RECT 58.240000 172.780000 58.795000 172.850000 ;
      RECT 58.240000 172.850000 58.865000 172.920000 ;
      RECT 58.240000 172.920000 58.935000 172.990000 ;
      RECT 58.240000 172.990000 59.005000 173.060000 ;
      RECT 58.240000 173.060000 59.075000 173.130000 ;
      RECT 58.240000 173.130000 59.145000 173.200000 ;
      RECT 58.240000 173.200000 59.215000 173.270000 ;
      RECT 58.240000 173.270000 59.285000 173.340000 ;
      RECT 58.240000 173.340000 59.355000 173.410000 ;
      RECT 58.240000 173.410000 59.425000 173.480000 ;
      RECT 58.240000 173.480000 59.495000 173.550000 ;
      RECT 58.240000 173.550000 59.565000 173.620000 ;
      RECT 58.240000 173.620000 59.635000 173.690000 ;
      RECT 58.240000 173.690000 59.705000 173.760000 ;
      RECT 58.240000 173.760000 59.775000 173.830000 ;
      RECT 58.240000 173.830000 59.845000 173.900000 ;
      RECT 58.240000 173.900000 59.915000 173.970000 ;
      RECT 58.240000 173.970000 59.985000 174.040000 ;
      RECT 58.240000 174.040000 60.055000 174.110000 ;
      RECT 58.240000 174.110000 60.125000 174.180000 ;
      RECT 58.240000 174.180000 60.195000 174.250000 ;
      RECT 58.240000 174.250000 60.265000 174.320000 ;
      RECT 58.240000 174.320000 60.335000 174.390000 ;
      RECT 58.240000 174.390000 60.405000 174.460000 ;
      RECT 58.240000 174.460000 60.475000 174.530000 ;
      RECT 58.240000 174.530000 60.545000 174.600000 ;
      RECT 58.240000 174.600000 60.615000 174.670000 ;
      RECT 58.240000 174.670000 60.685000 174.740000 ;
      RECT 58.240000 174.740000 60.755000 174.810000 ;
      RECT 58.240000 174.760000 60.970000 181.760000 ;
      RECT 58.240000 174.810000 60.825000 174.815000 ;
      RECT 58.240000 174.815000 60.830000 181.760000 ;
      RECT 67.480000 190.280000 75.000000 195.355000 ;
      RECT 67.480000 190.295000 75.000000 200.000000 ;
      RECT 70.480000 193.295000 72.000000 197.000000 ;
      RECT 74.430000   0.000000 75.000000 190.155000 ;
      RECT 74.570000   0.000000 75.000000 190.295000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.195000  36.635000 ;
      RECT  0.000000  36.635000  0.810000  37.250000 ;
      RECT  0.000000  36.730000  0.150000  36.880000 ;
      RECT  0.000000  36.880000  0.300000  37.030000 ;
      RECT  0.000000  37.030000  0.450000  37.180000 ;
      RECT  0.000000  37.180000  0.600000  37.290000 ;
      RECT  0.000000  37.250000  0.810000  46.220000 ;
      RECT  0.000000  37.290000  0.710000  46.180000 ;
      RECT  0.000000  46.180000  0.560000  46.330000 ;
      RECT  0.000000  46.220000  0.195000  46.835000 ;
      RECT  0.000000  46.330000  0.410000  46.480000 ;
      RECT  0.000000  46.480000  0.260000  46.630000 ;
      RECT  0.000000  46.630000  0.110000  46.780000 ;
      RECT  0.000000  46.835000  0.195000 173.455000 ;
      RECT  0.000000 173.455000  2.760000 185.195000 ;
      RECT  0.000000 173.555000 14.250000 173.705000 ;
      RECT  0.000000 173.705000 14.100000 173.855000 ;
      RECT  0.000000 173.855000 13.950000 174.005000 ;
      RECT  0.000000 174.005000 13.800000 174.155000 ;
      RECT  0.000000 174.155000 13.650000 174.305000 ;
      RECT  0.000000 174.305000 13.500000 174.455000 ;
      RECT  0.000000 174.455000 13.350000 174.605000 ;
      RECT  0.000000 174.605000 13.200000 174.755000 ;
      RECT  0.000000 174.755000 13.050000 174.905000 ;
      RECT  0.000000 174.905000 12.900000 175.055000 ;
      RECT  0.000000 175.055000 12.750000 175.205000 ;
      RECT  0.000000 175.205000 12.600000 175.355000 ;
      RECT  0.000000 175.355000 12.450000 175.505000 ;
      RECT  0.000000 175.505000 12.300000 175.655000 ;
      RECT  0.000000 175.655000 12.150000 175.805000 ;
      RECT  0.000000 175.805000 12.000000 175.955000 ;
      RECT  0.000000 175.955000 11.850000 176.105000 ;
      RECT  0.000000 176.105000 11.700000 176.255000 ;
      RECT  0.000000 176.255000 11.550000 176.405000 ;
      RECT  0.000000 176.405000 11.400000 176.555000 ;
      RECT  0.000000 176.555000 11.250000 176.705000 ;
      RECT  0.000000 176.705000 11.100000 176.855000 ;
      RECT  0.000000 176.855000 10.950000 177.005000 ;
      RECT  0.000000 177.005000 10.800000 177.155000 ;
      RECT  0.000000 177.155000 10.650000 177.305000 ;
      RECT  0.000000 177.305000 10.500000 177.455000 ;
      RECT  0.000000 177.455000 10.350000 177.605000 ;
      RECT  0.000000 177.605000 10.200000 177.755000 ;
      RECT  0.000000 177.755000 10.050000 177.905000 ;
      RECT  0.000000 177.905000  9.900000 178.055000 ;
      RECT  0.000000 178.055000  9.750000 178.205000 ;
      RECT  0.000000 178.205000  9.600000 178.355000 ;
      RECT  0.000000 178.355000  9.450000 178.505000 ;
      RECT  0.000000 178.505000  9.300000 178.655000 ;
      RECT  0.000000 178.655000  9.150000 178.805000 ;
      RECT  0.000000 178.805000  9.000000 178.955000 ;
      RECT  0.000000 178.955000  8.850000 179.105000 ;
      RECT  0.000000 179.105000  8.700000 179.255000 ;
      RECT  0.000000 179.255000  8.550000 179.405000 ;
      RECT  0.000000 179.405000  8.400000 179.555000 ;
      RECT  0.000000 179.555000  8.250000 179.705000 ;
      RECT  0.000000 179.705000  8.100000 179.855000 ;
      RECT  0.000000 179.855000  7.950000 180.005000 ;
      RECT  0.000000 180.005000  7.800000 180.155000 ;
      RECT  0.000000 180.155000  7.650000 180.305000 ;
      RECT  0.000000 180.305000  7.500000 180.455000 ;
      RECT  0.000000 180.455000  7.350000 180.605000 ;
      RECT  0.000000 180.605000  7.200000 180.755000 ;
      RECT  0.000000 180.755000  7.050000 180.905000 ;
      RECT  0.000000 180.905000  6.900000 181.055000 ;
      RECT  0.000000 181.055000  6.750000 181.205000 ;
      RECT  0.000000 181.205000  6.600000 181.355000 ;
      RECT  0.000000 181.355000  6.450000 181.505000 ;
      RECT  0.000000 181.505000  6.300000 181.655000 ;
      RECT  0.000000 181.655000  6.150000 181.805000 ;
      RECT  0.000000 181.805000  6.000000 181.955000 ;
      RECT  0.000000 181.955000  5.850000 182.105000 ;
      RECT  0.000000 182.105000  5.700000 182.255000 ;
      RECT  0.000000 182.255000  5.550000 182.405000 ;
      RECT  0.000000 182.405000  5.400000 182.555000 ;
      RECT  0.000000 182.555000  5.250000 182.705000 ;
      RECT  0.000000 182.705000  5.100000 182.855000 ;
      RECT  0.000000 182.855000  4.950000 183.005000 ;
      RECT  0.000000 183.005000  4.800000 183.155000 ;
      RECT  0.000000 183.155000  4.650000 183.305000 ;
      RECT  0.000000 183.305000  4.500000 183.455000 ;
      RECT  0.000000 183.455000  4.350000 183.605000 ;
      RECT  0.000000 183.605000  4.200000 183.755000 ;
      RECT  0.000000 183.755000  4.050000 183.905000 ;
      RECT  0.000000 183.905000  3.900000 184.055000 ;
      RECT  0.000000 184.055000  3.750000 184.205000 ;
      RECT  0.000000 184.205000  3.600000 184.355000 ;
      RECT  0.000000 184.355000  3.450000 184.505000 ;
      RECT  0.000000 184.505000  3.300000 184.655000 ;
      RECT  0.000000 184.655000  3.150000 184.805000 ;
      RECT  0.000000 184.805000  3.000000 184.955000 ;
      RECT  0.000000 184.955000  2.850000 185.105000 ;
      RECT  0.000000 185.105000  2.760000 185.195000 ;
      RECT  0.000000 185.195000  2.760000 200.000000 ;
      RECT  0.000000 185.195000  2.760000 200.000000 ;
      RECT  3.000000 176.555000  7.005000 176.705000 ;
      RECT  3.000000 176.555000  7.005000 176.705000 ;
      RECT  3.000000 176.705000  6.855000 176.855000 ;
      RECT  3.000000 176.705000  6.855000 176.855000 ;
      RECT  3.000000 176.855000  6.705000 177.005000 ;
      RECT  3.000000 176.855000  6.705000 177.005000 ;
      RECT  3.000000 177.005000  6.555000 177.155000 ;
      RECT  3.000000 177.005000  6.555000 177.155000 ;
      RECT  3.000000 177.155000  6.405000 177.305000 ;
      RECT  3.000000 177.155000  6.405000 177.305000 ;
      RECT  3.000000 177.305000  6.255000 177.455000 ;
      RECT  3.000000 177.305000  6.255000 177.455000 ;
      RECT  3.000000 177.455000  6.105000 177.605000 ;
      RECT  3.000000 177.455000  6.105000 177.605000 ;
      RECT  3.000000 177.605000  5.955000 177.755000 ;
      RECT  3.000000 177.605000  5.955000 177.755000 ;
      RECT  3.000000 177.755000  5.805000 177.905000 ;
      RECT  3.000000 177.755000  5.805000 177.905000 ;
      RECT  3.000000 177.905000  5.655000 178.055000 ;
      RECT  3.000000 177.905000  5.655000 178.055000 ;
      RECT  3.000000 178.055000  5.505000 178.205000 ;
      RECT  3.000000 178.055000  5.505000 178.205000 ;
      RECT  3.000000 178.205000  5.355000 178.355000 ;
      RECT  3.000000 178.205000  5.355000 178.355000 ;
      RECT  3.000000 178.355000  5.205000 178.505000 ;
      RECT  3.000000 178.355000  5.205000 178.505000 ;
      RECT  3.000000 178.505000  5.055000 178.655000 ;
      RECT  3.000000 178.505000  5.055000 178.655000 ;
      RECT  3.000000 178.655000  4.905000 178.805000 ;
      RECT  3.000000 178.655000  4.905000 178.805000 ;
      RECT  3.000000 178.805000  4.755000 178.955000 ;
      RECT  3.000000 178.805000  4.755000 178.955000 ;
      RECT  3.000000 178.955000  4.605000 179.105000 ;
      RECT  3.000000 178.955000  4.605000 179.105000 ;
      RECT  3.000000 179.105000  4.455000 179.255000 ;
      RECT  3.000000 179.105000  4.455000 179.255000 ;
      RECT  3.000000 179.255000  4.305000 179.405000 ;
      RECT  3.000000 179.255000  4.305000 179.405000 ;
      RECT  3.000000 179.405000  4.155000 179.555000 ;
      RECT  3.000000 179.405000  4.155000 179.555000 ;
      RECT  3.000000 179.555000  4.005000 179.705000 ;
      RECT  3.000000 179.555000  4.005000 179.705000 ;
      RECT  3.000000 179.705000  3.855000 179.855000 ;
      RECT  3.000000 179.705000  3.855000 179.855000 ;
      RECT  3.000000 179.855000  3.705000 180.005000 ;
      RECT  3.000000 179.855000  3.705000 180.005000 ;
      RECT  3.000000 180.005000  3.555000 180.155000 ;
      RECT  3.000000 180.005000  3.555000 180.155000 ;
      RECT  3.000000 180.155000  3.405000 180.305000 ;
      RECT  3.000000 180.155000  3.405000 180.305000 ;
      RECT  3.000000 180.305000  3.255000 180.455000 ;
      RECT  3.000000 180.305000  3.255000 180.455000 ;
      RECT  3.000000 180.455000  3.105000 180.605000 ;
      RECT  3.000000 180.455000  3.105000 180.605000 ;
      RECT  3.000000 180.605000  3.005000 180.705000 ;
      RECT  3.000000 180.605000  3.005000 180.705000 ;
      RECT 13.800000 101.520000 15.100000 102.035000 ;
      RECT 13.800000 102.035000 15.100000 172.855000 ;
      RECT 13.800000 172.855000 14.500000 173.455000 ;
      RECT 13.900000 101.560000 15.425000 101.710000 ;
      RECT 13.900000 101.710000 15.275000 101.860000 ;
      RECT 13.900000 101.860000 15.125000 102.010000 ;
      RECT 13.900000 102.010000 15.100000 102.035000 ;
      RECT 13.900000 102.035000 15.100000 172.855000 ;
      RECT 13.900000 172.855000 14.950000 173.005000 ;
      RECT 13.900000 173.005000 14.800000 173.155000 ;
      RECT 13.900000 173.155000 14.650000 173.305000 ;
      RECT 13.900000 173.305000 14.500000 173.455000 ;
      RECT 13.900000 173.455000 14.400000 173.555000 ;
      RECT 14.020000 101.440000 15.575000 101.560000 ;
      RECT 14.170000 101.290000 15.695000 101.440000 ;
      RECT 14.320000 101.140000 15.845000 101.290000 ;
      RECT 14.470000 100.990000 15.995000 101.140000 ;
      RECT 14.620000 100.840000 16.145000 100.990000 ;
      RECT 14.770000 100.690000 16.295000 100.840000 ;
      RECT 14.920000 100.540000 16.445000 100.690000 ;
      RECT 15.070000 100.390000 16.595000 100.540000 ;
      RECT 15.220000 100.240000 16.745000 100.390000 ;
      RECT 15.370000 100.090000 16.895000 100.240000 ;
      RECT 15.520000  99.940000 17.045000 100.090000 ;
      RECT 15.670000  99.790000 17.195000  99.940000 ;
      RECT 15.820000  99.640000 17.345000  99.790000 ;
      RECT 15.970000  99.490000 17.495000  99.640000 ;
      RECT 16.120000  99.340000 17.645000  99.490000 ;
      RECT 16.270000  99.190000 17.795000  99.340000 ;
      RECT 16.420000  99.040000 17.945000  99.190000 ;
      RECT 16.570000  98.890000 18.095000  99.040000 ;
      RECT 16.720000  98.740000 18.245000  98.890000 ;
      RECT 16.870000  98.590000 18.395000  98.740000 ;
      RECT 17.020000  98.440000 18.545000  98.590000 ;
      RECT 17.170000  98.290000 18.695000  98.440000 ;
      RECT 17.320000  98.140000 18.845000  98.290000 ;
      RECT 17.470000  97.990000 18.995000  98.140000 ;
      RECT 17.620000  97.840000 19.145000  97.990000 ;
      RECT 17.770000  97.690000 19.295000  97.840000 ;
      RECT 17.920000  97.540000 19.445000  97.690000 ;
      RECT 18.070000  97.390000 19.595000  97.540000 ;
      RECT 18.220000  97.240000 19.745000  97.390000 ;
      RECT 18.370000  97.090000 19.895000  97.240000 ;
      RECT 18.520000  96.940000 20.045000  97.090000 ;
      RECT 18.670000  96.790000 20.195000  96.940000 ;
      RECT 18.820000  96.640000 20.345000  96.790000 ;
      RECT 18.970000  96.490000 20.495000  96.640000 ;
      RECT 19.120000  96.340000 20.645000  96.490000 ;
      RECT 19.270000  96.190000 20.795000  96.340000 ;
      RECT 19.420000  96.040000 20.945000  96.190000 ;
      RECT 19.570000  95.890000 21.095000  96.040000 ;
      RECT 19.720000  95.740000 21.245000  95.890000 ;
      RECT 19.870000  95.590000 21.395000  95.740000 ;
      RECT 20.020000  95.440000 21.545000  95.590000 ;
      RECT 20.170000  95.290000 21.695000  95.440000 ;
      RECT 20.320000  95.140000 21.845000  95.290000 ;
      RECT 20.470000  94.990000 21.995000  95.140000 ;
      RECT 20.620000  94.840000 22.145000  94.990000 ;
      RECT 20.770000  94.690000 22.295000  94.840000 ;
      RECT 20.920000  94.540000 22.445000  94.690000 ;
      RECT 21.070000  94.390000 22.595000  94.540000 ;
      RECT 21.220000  94.240000 22.745000  94.390000 ;
      RECT 21.370000  94.090000 22.895000  94.240000 ;
      RECT 21.520000  93.940000 23.045000  94.090000 ;
      RECT 21.670000  93.790000 23.195000  93.940000 ;
      RECT 21.695000  93.765000 23.345000  93.790000 ;
      RECT 21.845000  93.615000 23.345000  93.765000 ;
      RECT 21.900000 104.845000 25.530000 168.965000 ;
      RECT 21.900000 104.845000 25.530000 168.965000 ;
      RECT 21.900000 168.965000 25.530000 172.475000 ;
      RECT 21.970000 104.775000 25.530000 104.845000 ;
      RECT 21.995000  93.465000 23.345000  93.615000 ;
      RECT 22.050000 168.965000 25.530000 169.115000 ;
      RECT 22.120000 104.625000 25.530000 104.775000 ;
      RECT 22.145000  93.315000 23.345000  93.465000 ;
      RECT 22.200000 169.115000 25.530000 169.265000 ;
      RECT 22.270000 104.475000 25.530000 104.625000 ;
      RECT 22.295000  93.165000 23.345000  93.315000 ;
      RECT 22.350000 169.265000 25.530000 169.415000 ;
      RECT 22.420000 104.325000 25.530000 104.475000 ;
      RECT 22.445000  93.015000 23.345000  93.165000 ;
      RECT 22.500000 169.415000 25.530000 169.565000 ;
      RECT 22.570000 104.175000 25.530000 104.325000 ;
      RECT 22.595000  92.865000 23.345000  93.015000 ;
      RECT 22.650000 169.565000 25.530000 169.715000 ;
      RECT 22.720000 104.025000 25.530000 104.175000 ;
      RECT 22.745000  92.715000 23.345000  92.865000 ;
      RECT 22.800000 169.715000 25.530000 169.865000 ;
      RECT 22.870000 103.875000 25.530000 104.025000 ;
      RECT 22.895000  92.565000 23.345000  92.715000 ;
      RECT 22.945000  92.375000 23.345000  93.790000 ;
      RECT 22.950000 169.865000 25.530000 170.015000 ;
      RECT 23.020000 103.725000 25.530000 103.875000 ;
      RECT 23.045000  92.415000 23.345000  92.565000 ;
      RECT 23.100000 170.015000 25.530000 170.165000 ;
      RECT 23.170000 103.575000 25.530000 103.725000 ;
      RECT 23.195000  92.265000 23.345000  92.415000 ;
      RECT 23.250000 170.165000 25.530000 170.315000 ;
      RECT 23.320000 103.425000 25.530000 103.575000 ;
      RECT 23.400000 170.315000 25.530000 170.465000 ;
      RECT 23.470000 103.275000 25.530000 103.425000 ;
      RECT 23.550000 170.465000 25.530000 170.615000 ;
      RECT 23.620000 103.125000 25.530000 103.275000 ;
      RECT 23.700000 170.615000 25.530000 170.765000 ;
      RECT 23.770000 102.975000 25.530000 103.125000 ;
      RECT 23.850000 170.765000 25.530000 170.915000 ;
      RECT 23.920000 102.825000 25.530000 102.975000 ;
      RECT 24.000000 170.915000 25.530000 171.065000 ;
      RECT 24.070000 102.675000 25.530000 102.825000 ;
      RECT 24.150000 171.065000 25.530000 171.215000 ;
      RECT 24.220000 102.525000 25.530000 102.675000 ;
      RECT 24.300000 171.215000 25.530000 171.365000 ;
      RECT 24.370000 102.375000 25.530000 102.525000 ;
      RECT 24.450000 171.365000 25.530000 171.515000 ;
      RECT 24.520000 102.225000 25.530000 102.375000 ;
      RECT 24.520000 102.225000 25.530000 104.845000 ;
      RECT 24.525000 102.220000 25.530000 102.225000 ;
      RECT 24.600000 171.515000 25.530000 171.665000 ;
      RECT 24.675000 102.070000 25.535000 102.220000 ;
      RECT 24.695000   0.000000 25.495000  90.225000 ;
      RECT 24.695000  90.225000 25.095000  90.625000 ;
      RECT 24.750000 171.665000 25.530000 171.815000 ;
      RECT 24.795000   0.000000 25.495000  90.225000 ;
      RECT 24.795000  90.225000 25.345000  90.375000 ;
      RECT 24.795000  90.375000 25.195000  90.525000 ;
      RECT 24.795000  90.525000 25.045000  90.675000 ;
      RECT 24.795000  90.675000 24.895000  90.825000 ;
      RECT 24.825000 101.920000 25.685000 102.070000 ;
      RECT 24.900000 171.815000 25.530000 171.965000 ;
      RECT 24.975000 101.770000 25.835000 101.920000 ;
      RECT 25.050000 171.965000 25.530000 172.115000 ;
      RECT 25.125000 101.620000 25.985000 101.770000 ;
      RECT 25.200000 172.115000 25.530000 172.265000 ;
      RECT 25.275000 101.470000 26.135000 101.620000 ;
      RECT 25.350000 172.265000 25.530000 172.415000 ;
      RECT 25.410000 172.475000 25.530000 200.000000 ;
      RECT 25.425000 101.320000 26.285000 101.470000 ;
      RECT 25.500000 172.415000 25.530000 172.565000 ;
      RECT 25.575000 101.170000 26.435000 101.320000 ;
      RECT 25.725000 101.020000 26.585000 101.170000 ;
      RECT 25.875000 100.870000 26.735000 101.020000 ;
      RECT 26.025000 100.720000 26.885000 100.870000 ;
      RECT 26.175000 100.570000 27.035000 100.720000 ;
      RECT 26.325000 100.420000 27.185000 100.570000 ;
      RECT 26.475000 100.270000 27.335000 100.420000 ;
      RECT 26.625000 100.120000 27.485000 100.270000 ;
      RECT 26.775000  99.970000 27.635000 100.120000 ;
      RECT 26.925000  99.820000 27.785000  99.970000 ;
      RECT 27.075000  99.670000 27.935000  99.820000 ;
      RECT 27.225000  99.520000 28.085000  99.670000 ;
      RECT 27.375000  99.370000 28.235000  99.520000 ;
      RECT 27.525000  99.220000 28.385000  99.370000 ;
      RECT 27.675000  99.070000 28.535000  99.220000 ;
      RECT 27.825000  98.920000 28.685000  99.070000 ;
      RECT 27.975000  98.770000 28.835000  98.920000 ;
      RECT 28.125000  98.620000 28.985000  98.770000 ;
      RECT 28.275000  98.470000 29.135000  98.620000 ;
      RECT 28.425000  98.320000 29.285000  98.470000 ;
      RECT 28.575000  98.170000 29.435000  98.320000 ;
      RECT 28.725000  98.020000 29.585000  98.170000 ;
      RECT 28.875000  97.870000 29.735000  98.020000 ;
      RECT 29.025000  97.720000 29.885000  97.870000 ;
      RECT 29.175000  97.570000 30.035000  97.720000 ;
      RECT 29.325000  97.420000 30.185000  97.570000 ;
      RECT 29.475000  97.270000 30.335000  97.420000 ;
      RECT 29.625000  97.120000 30.485000  97.270000 ;
      RECT 29.775000  96.970000 30.635000  97.120000 ;
      RECT 29.925000  93.265000 31.545000  96.210000 ;
      RECT 29.925000  93.265000 31.545000  96.210000 ;
      RECT 29.925000  96.210000 30.935000  96.820000 ;
      RECT 29.925000  96.210000 31.395000  96.360000 ;
      RECT 29.925000  96.360000 31.245000  96.510000 ;
      RECT 29.925000  96.510000 31.095000  96.660000 ;
      RECT 29.925000  96.660000 30.945000  96.810000 ;
      RECT 29.925000  96.810000 30.935000  96.820000 ;
      RECT 29.925000  96.820000 30.785000  96.970000 ;
      RECT 29.950000  93.240000 31.520000  93.265000 ;
      RECT 30.100000  93.090000 31.370000  93.240000 ;
      RECT 30.250000  92.940000 31.220000  93.090000 ;
      RECT 30.400000  92.790000 31.070000  92.940000 ;
      RECT 30.400000  92.790000 31.545000  93.265000 ;
      RECT 32.330000  99.865000 37.490000 110.785000 ;
      RECT 32.330000 105.025000 37.490000 105.820000 ;
      RECT 32.330000 105.025000 37.490000 105.820000 ;
      RECT 32.330000 105.820000 37.490000 105.970000 ;
      RECT 32.330000 105.820000 37.490000 105.970000 ;
      RECT 32.330000 105.820000 42.455000 110.785000 ;
      RECT 32.330000 105.820000 42.455000 175.185000 ;
      RECT 32.330000 105.970000 37.640000 106.120000 ;
      RECT 32.330000 105.970000 37.640000 106.120000 ;
      RECT 32.330000 106.120000 37.790000 106.270000 ;
      RECT 32.330000 106.120000 37.790000 106.270000 ;
      RECT 32.330000 106.270000 37.940000 106.420000 ;
      RECT 32.330000 106.270000 37.940000 106.420000 ;
      RECT 32.330000 106.420000 38.090000 106.570000 ;
      RECT 32.330000 106.420000 38.090000 106.570000 ;
      RECT 32.330000 106.570000 38.240000 106.720000 ;
      RECT 32.330000 106.570000 38.240000 106.720000 ;
      RECT 32.330000 106.720000 38.390000 106.870000 ;
      RECT 32.330000 106.720000 38.390000 106.870000 ;
      RECT 32.330000 106.870000 38.540000 107.020000 ;
      RECT 32.330000 106.870000 38.540000 107.020000 ;
      RECT 32.330000 107.020000 38.690000 107.170000 ;
      RECT 32.330000 107.020000 38.690000 107.170000 ;
      RECT 32.330000 107.170000 38.840000 107.320000 ;
      RECT 32.330000 107.170000 38.840000 107.320000 ;
      RECT 32.330000 107.320000 38.990000 107.470000 ;
      RECT 32.330000 107.320000 38.990000 107.470000 ;
      RECT 32.330000 107.470000 39.140000 107.620000 ;
      RECT 32.330000 107.470000 39.140000 107.620000 ;
      RECT 32.330000 107.620000 39.290000 107.770000 ;
      RECT 32.330000 107.620000 39.290000 107.770000 ;
      RECT 32.330000 107.770000 39.440000 107.920000 ;
      RECT 32.330000 107.770000 39.440000 107.920000 ;
      RECT 32.330000 107.920000 39.590000 108.070000 ;
      RECT 32.330000 107.920000 39.590000 108.070000 ;
      RECT 32.330000 108.070000 39.740000 108.220000 ;
      RECT 32.330000 108.070000 39.740000 108.220000 ;
      RECT 32.330000 108.220000 39.890000 108.370000 ;
      RECT 32.330000 108.220000 39.890000 108.370000 ;
      RECT 32.330000 108.370000 40.040000 108.520000 ;
      RECT 32.330000 108.370000 40.040000 108.520000 ;
      RECT 32.330000 108.520000 40.190000 108.670000 ;
      RECT 32.330000 108.520000 40.190000 108.670000 ;
      RECT 32.330000 108.670000 40.340000 108.820000 ;
      RECT 32.330000 108.670000 40.340000 108.820000 ;
      RECT 32.330000 108.820000 40.490000 108.970000 ;
      RECT 32.330000 108.820000 40.490000 108.970000 ;
      RECT 32.330000 108.970000 40.640000 109.120000 ;
      RECT 32.330000 108.970000 40.640000 109.120000 ;
      RECT 32.330000 109.120000 40.790000 109.270000 ;
      RECT 32.330000 109.120000 40.790000 109.270000 ;
      RECT 32.330000 109.270000 40.940000 109.420000 ;
      RECT 32.330000 109.270000 40.940000 109.420000 ;
      RECT 32.330000 109.420000 41.090000 109.570000 ;
      RECT 32.330000 109.420000 41.090000 109.570000 ;
      RECT 32.330000 109.570000 41.240000 109.720000 ;
      RECT 32.330000 109.570000 41.240000 109.720000 ;
      RECT 32.330000 109.720000 41.390000 109.870000 ;
      RECT 32.330000 109.720000 41.390000 109.870000 ;
      RECT 32.330000 109.870000 41.540000 110.020000 ;
      RECT 32.330000 109.870000 41.540000 110.020000 ;
      RECT 32.330000 110.020000 41.690000 110.170000 ;
      RECT 32.330000 110.020000 41.690000 110.170000 ;
      RECT 32.330000 110.170000 41.840000 110.320000 ;
      RECT 32.330000 110.170000 41.840000 110.320000 ;
      RECT 32.330000 110.320000 41.990000 110.470000 ;
      RECT 32.330000 110.320000 41.990000 110.470000 ;
      RECT 32.330000 110.470000 42.140000 110.620000 ;
      RECT 32.330000 110.470000 42.140000 110.620000 ;
      RECT 32.330000 110.620000 42.290000 110.770000 ;
      RECT 32.330000 110.620000 42.290000 110.770000 ;
      RECT 32.330000 110.770000 42.440000 110.785000 ;
      RECT 32.330000 110.770000 42.440000 110.785000 ;
      RECT 32.330000 110.785000 42.455000 170.295000 ;
      RECT 32.330000 110.785000 42.455000 170.295000 ;
      RECT 32.330000 170.295000 37.565000 175.185000 ;
      RECT 32.390000 104.965000 37.490000 105.025000 ;
      RECT 32.390000 104.965000 37.490000 105.025000 ;
      RECT 32.480000 170.295000 42.305000 170.445000 ;
      RECT 32.480000 170.295000 42.305000 170.445000 ;
      RECT 32.540000 104.815000 37.490000 104.965000 ;
      RECT 32.540000 104.815000 37.490000 104.965000 ;
      RECT 32.630000 170.445000 42.155000 170.595000 ;
      RECT 32.630000 170.445000 42.155000 170.595000 ;
      RECT 32.690000 104.665000 37.490000 104.815000 ;
      RECT 32.690000 104.665000 37.490000 104.815000 ;
      RECT 32.780000 170.595000 42.005000 170.745000 ;
      RECT 32.780000 170.595000 42.005000 170.745000 ;
      RECT 32.840000 104.515000 37.490000 104.665000 ;
      RECT 32.840000 104.515000 37.490000 104.665000 ;
      RECT 32.930000 170.745000 41.855000 170.895000 ;
      RECT 32.930000 170.745000 41.855000 170.895000 ;
      RECT 32.990000 104.365000 37.490000 104.515000 ;
      RECT 32.990000 104.365000 37.490000 104.515000 ;
      RECT 33.080000 170.895000 41.705000 171.045000 ;
      RECT 33.080000 170.895000 41.705000 171.045000 ;
      RECT 33.140000 104.215000 37.490000 104.365000 ;
      RECT 33.140000 104.215000 37.490000 104.365000 ;
      RECT 33.230000 171.045000 41.555000 171.195000 ;
      RECT 33.230000 171.045000 41.555000 171.195000 ;
      RECT 33.290000 104.065000 37.490000 104.215000 ;
      RECT 33.290000 104.065000 37.490000 104.215000 ;
      RECT 33.380000 171.195000 41.405000 171.345000 ;
      RECT 33.380000 171.195000 41.405000 171.345000 ;
      RECT 33.440000 103.915000 37.490000 104.065000 ;
      RECT 33.440000 103.915000 37.490000 104.065000 ;
      RECT 33.530000 171.345000 41.255000 171.495000 ;
      RECT 33.530000 171.345000 41.255000 171.495000 ;
      RECT 33.590000 103.765000 37.490000 103.915000 ;
      RECT 33.590000 103.765000 37.490000 103.915000 ;
      RECT 33.680000 171.495000 41.105000 171.645000 ;
      RECT 33.680000 171.495000 41.105000 171.645000 ;
      RECT 33.740000 103.615000 37.490000 103.765000 ;
      RECT 33.740000 103.615000 37.490000 103.765000 ;
      RECT 33.830000 171.645000 40.955000 171.795000 ;
      RECT 33.830000 171.645000 40.955000 171.795000 ;
      RECT 33.890000 103.465000 37.490000 103.615000 ;
      RECT 33.890000 103.465000 37.490000 103.615000 ;
      RECT 33.980000 171.795000 40.805000 171.945000 ;
      RECT 33.980000 171.795000 40.805000 171.945000 ;
      RECT 34.040000 103.315000 37.490000 103.465000 ;
      RECT 34.040000 103.315000 37.490000 103.465000 ;
      RECT 34.130000 171.945000 40.655000 172.095000 ;
      RECT 34.130000 171.945000 40.655000 172.095000 ;
      RECT 34.190000 103.165000 37.490000 103.315000 ;
      RECT 34.190000 103.165000 37.490000 103.315000 ;
      RECT 34.280000 172.095000 40.505000 172.245000 ;
      RECT 34.280000 172.095000 40.505000 172.245000 ;
      RECT 34.340000 103.015000 37.490000 103.165000 ;
      RECT 34.340000 103.015000 37.490000 103.165000 ;
      RECT 34.430000 172.245000 40.355000 172.395000 ;
      RECT 34.430000 172.245000 40.355000 172.395000 ;
      RECT 34.490000 102.865000 37.490000 103.015000 ;
      RECT 34.490000 102.865000 37.490000 103.015000 ;
      RECT 34.580000 172.395000 40.205000 172.545000 ;
      RECT 34.580000 172.395000 40.205000 172.545000 ;
      RECT 34.640000 102.715000 37.490000 102.865000 ;
      RECT 34.640000 102.715000 37.490000 102.865000 ;
      RECT 34.730000 172.545000 40.055000 172.695000 ;
      RECT 34.730000 172.545000 40.055000 172.695000 ;
      RECT 34.790000 102.565000 37.490000 102.715000 ;
      RECT 34.790000 102.565000 37.490000 102.715000 ;
      RECT 34.880000 172.695000 39.905000 172.845000 ;
      RECT 34.880000 172.695000 39.905000 172.845000 ;
      RECT 34.940000 102.415000 37.490000 102.565000 ;
      RECT 34.940000 102.415000 37.490000 102.565000 ;
      RECT 35.030000 172.845000 39.755000 172.995000 ;
      RECT 35.030000 172.845000 39.755000 172.995000 ;
      RECT 35.090000 102.265000 37.490000 102.415000 ;
      RECT 35.090000 102.265000 37.490000 102.415000 ;
      RECT 35.180000 172.995000 39.605000 173.145000 ;
      RECT 35.180000 172.995000 39.605000 173.145000 ;
      RECT 35.240000 102.115000 37.490000 102.265000 ;
      RECT 35.240000 102.115000 37.490000 102.265000 ;
      RECT 35.330000 173.145000 39.455000 173.295000 ;
      RECT 35.330000 173.145000 39.455000 173.295000 ;
      RECT 35.390000 101.965000 37.490000 102.115000 ;
      RECT 35.390000 101.965000 37.490000 102.115000 ;
      RECT 35.480000 173.295000 39.305000 173.445000 ;
      RECT 35.480000 173.295000 39.305000 173.445000 ;
      RECT 35.540000 101.815000 37.490000 101.965000 ;
      RECT 35.540000 101.815000 37.490000 101.965000 ;
      RECT 35.630000 173.445000 39.155000 173.595000 ;
      RECT 35.630000 173.445000 39.155000 173.595000 ;
      RECT 35.690000 101.665000 37.490000 101.815000 ;
      RECT 35.690000 101.665000 37.490000 101.815000 ;
      RECT 35.780000 173.595000 39.005000 173.745000 ;
      RECT 35.780000 173.595000 39.005000 173.745000 ;
      RECT 35.840000 101.515000 37.490000 101.665000 ;
      RECT 35.840000 101.515000 37.490000 101.665000 ;
      RECT 35.930000 173.745000 38.855000 173.895000 ;
      RECT 35.930000 173.745000 38.855000 173.895000 ;
      RECT 35.990000 101.365000 37.490000 101.515000 ;
      RECT 35.990000 101.365000 37.490000 101.515000 ;
      RECT 36.080000 173.895000 38.705000 174.045000 ;
      RECT 36.080000 173.895000 38.705000 174.045000 ;
      RECT 36.140000 101.215000 37.490000 101.365000 ;
      RECT 36.140000 101.215000 37.490000 101.365000 ;
      RECT 36.230000 174.045000 38.555000 174.195000 ;
      RECT 36.230000 174.045000 38.555000 174.195000 ;
      RECT 36.290000 101.065000 37.490000 101.215000 ;
      RECT 36.290000 101.065000 37.490000 101.215000 ;
      RECT 36.380000 174.195000 38.405000 174.345000 ;
      RECT 36.380000 174.195000 38.405000 174.345000 ;
      RECT 36.440000 100.915000 37.490000 101.065000 ;
      RECT 36.440000 100.915000 37.490000 101.065000 ;
      RECT 36.530000 174.345000 38.255000 174.495000 ;
      RECT 36.530000 174.345000 38.255000 174.495000 ;
      RECT 36.590000 100.765000 37.490000 100.915000 ;
      RECT 36.590000 100.765000 37.490000 100.915000 ;
      RECT 36.680000 174.495000 38.105000 174.645000 ;
      RECT 36.680000 174.495000 38.105000 174.645000 ;
      RECT 36.740000 100.615000 37.490000 100.765000 ;
      RECT 36.740000 100.615000 37.490000 100.765000 ;
      RECT 36.830000 174.645000 37.955000 174.795000 ;
      RECT 36.830000 174.645000 37.955000 174.795000 ;
      RECT 36.890000 100.465000 37.490000 100.615000 ;
      RECT 36.890000 100.465000 37.490000 100.615000 ;
      RECT 36.980000 174.795000 37.805000 174.945000 ;
      RECT 36.980000 174.795000 37.805000 174.945000 ;
      RECT 37.040000 100.315000 37.490000 100.465000 ;
      RECT 37.040000 100.315000 37.490000 100.465000 ;
      RECT 37.130000 174.945000 37.655000 175.095000 ;
      RECT 37.130000 174.945000 37.655000 175.095000 ;
      RECT 37.190000 100.165000 37.490000 100.315000 ;
      RECT 37.190000 100.165000 37.490000 100.315000 ;
      RECT 37.220000 175.185000 37.565000 190.420000 ;
      RECT 37.220000 175.270000 37.305000 175.355000 ;
      RECT 37.220000 175.355000 37.565000 190.420000 ;
      RECT 37.220000 190.420000 49.375000 190.440000 ;
      RECT 37.220000 190.420000 49.375000 190.440000 ;
      RECT 37.220000 190.420000 49.375000 200.000000 ;
      RECT 37.220000 190.440000 75.000000 200.000000 ;
      RECT 37.220000 190.440000 75.000000 200.000000 ;
      RECT 37.280000 175.095000 37.505000 175.245000 ;
      RECT 37.280000 175.095000 37.505000 175.245000 ;
      RECT 37.295000   0.000000 37.490000 100.060000 ;
      RECT 37.295000 100.060000 37.490000 105.025000 ;
      RECT 37.340000 100.015000 37.490000 100.165000 ;
      RECT 37.340000 100.015000 37.490000 100.165000 ;
      RECT 37.390000 175.245000 37.395000 175.355000 ;
      RECT 37.390000 175.245000 37.395000 175.355000 ;
      RECT 37.480000 175.270000 37.565000 175.355000 ;
      RECT 43.240000 100.380000 44.860000 101.970000 ;
      RECT 43.240000 100.380000 44.860000 101.970000 ;
      RECT 43.240000 101.970000 44.860000 102.580000 ;
      RECT 43.265000 100.355000 44.835000 100.380000 ;
      RECT 43.390000 101.970000 44.860000 102.120000 ;
      RECT 43.415000 100.205000 44.685000 100.355000 ;
      RECT 43.540000 102.120000 44.860000 102.270000 ;
      RECT 43.565000 100.055000 44.535000 100.205000 ;
      RECT 43.690000 102.270000 44.860000 102.420000 ;
      RECT 43.715000  99.905000 44.385000 100.055000 ;
      RECT 43.715000  99.905000 44.860000 100.380000 ;
      RECT 43.840000 102.420000 44.860000 102.570000 ;
      RECT 43.850000 102.570000 44.860000 102.580000 ;
      RECT 43.850000 102.580000 50.265000 107.985000 ;
      RECT 44.000000 102.580000 44.860000 102.730000 ;
      RECT 44.150000 102.730000 45.010000 102.880000 ;
      RECT 44.300000 102.880000 45.160000 103.030000 ;
      RECT 44.450000 103.030000 45.310000 103.180000 ;
      RECT 44.600000 103.180000 45.460000 103.330000 ;
      RECT 44.750000 103.330000 45.610000 103.480000 ;
      RECT 44.900000 103.480000 45.760000 103.630000 ;
      RECT 45.050000 103.630000 45.910000 103.780000 ;
      RECT 45.200000 103.780000 46.060000 103.930000 ;
      RECT 45.350000 103.930000 46.210000 104.080000 ;
      RECT 45.500000 104.080000 46.360000 104.230000 ;
      RECT 45.650000 104.230000 46.510000 104.380000 ;
      RECT 45.800000 104.380000 46.660000 104.530000 ;
      RECT 45.950000 104.530000 46.810000 104.680000 ;
      RECT 46.100000 104.680000 46.960000 104.830000 ;
      RECT 46.250000 104.830000 47.110000 104.980000 ;
      RECT 46.400000 104.980000 47.260000 105.130000 ;
      RECT 46.550000 105.130000 47.410000 105.280000 ;
      RECT 46.700000 105.280000 47.560000 105.430000 ;
      RECT 46.850000 105.430000 47.710000 105.580000 ;
      RECT 47.000000 105.580000 47.860000 105.730000 ;
      RECT 47.150000 105.730000 48.010000 105.880000 ;
      RECT 47.300000 105.880000 48.160000 106.030000 ;
      RECT 47.450000 106.030000 48.310000 106.180000 ;
      RECT 47.600000 106.180000 48.460000 106.330000 ;
      RECT 47.750000 106.330000 48.610000 106.480000 ;
      RECT 47.900000 106.480000 48.760000 106.630000 ;
      RECT 48.050000 106.630000 48.910000 106.780000 ;
      RECT 48.200000 106.780000 49.060000 106.930000 ;
      RECT 48.350000 106.930000 49.210000 107.080000 ;
      RECT 48.500000 107.080000 49.360000 107.230000 ;
      RECT 48.650000 107.230000 49.510000 107.380000 ;
      RECT 48.800000 107.380000 49.660000 107.530000 ;
      RECT 48.950000 107.530000 49.810000 107.680000 ;
      RECT 49.100000 107.680000 49.960000 107.830000 ;
      RECT 49.250000 107.830000 50.110000 107.980000 ;
      RECT 49.255000 107.980000 50.260000 107.985000 ;
      RECT 49.255000 107.985000 50.265000 108.135000 ;
      RECT 49.255000 107.985000 52.885000 110.605000 ;
      RECT 49.255000 108.135000 50.415000 108.285000 ;
      RECT 49.255000 108.285000 50.565000 108.435000 ;
      RECT 49.255000 108.435000 50.715000 108.585000 ;
      RECT 49.255000 108.585000 50.865000 108.735000 ;
      RECT 49.255000 108.735000 51.015000 108.885000 ;
      RECT 49.255000 108.885000 51.165000 109.035000 ;
      RECT 49.255000 109.035000 51.315000 109.185000 ;
      RECT 49.255000 109.185000 51.465000 109.335000 ;
      RECT 49.255000 109.335000 51.615000 109.485000 ;
      RECT 49.255000 109.485000 51.765000 109.635000 ;
      RECT 49.255000 109.635000 51.915000 109.785000 ;
      RECT 49.255000 109.785000 52.065000 109.935000 ;
      RECT 49.255000 109.935000 52.215000 110.085000 ;
      RECT 49.255000 110.085000 52.365000 110.235000 ;
      RECT 49.255000 110.235000 52.515000 110.385000 ;
      RECT 49.255000 110.385000 52.665000 110.535000 ;
      RECT 49.255000 110.535000 52.815000 110.605000 ;
      RECT 49.255000 110.605000 52.885000 168.970000 ;
      RECT 49.255000 110.605000 52.885000 168.970000 ;
      RECT 49.255000 168.970000 49.375000 172.480000 ;
      RECT 49.255000 168.970000 52.735000 169.120000 ;
      RECT 49.255000 169.120000 52.585000 169.270000 ;
      RECT 49.255000 169.270000 52.435000 169.420000 ;
      RECT 49.255000 169.420000 52.285000 169.570000 ;
      RECT 49.255000 169.570000 52.135000 169.720000 ;
      RECT 49.255000 169.720000 51.985000 169.870000 ;
      RECT 49.255000 169.870000 51.835000 170.020000 ;
      RECT 49.255000 170.020000 51.685000 170.170000 ;
      RECT 49.255000 170.170000 51.535000 170.320000 ;
      RECT 49.255000 170.320000 51.385000 170.470000 ;
      RECT 49.255000 170.470000 51.235000 170.620000 ;
      RECT 49.255000 170.620000 51.085000 170.770000 ;
      RECT 49.255000 170.770000 50.935000 170.920000 ;
      RECT 49.255000 170.920000 50.785000 171.070000 ;
      RECT 49.255000 171.070000 50.635000 171.220000 ;
      RECT 49.255000 171.220000 50.485000 171.370000 ;
      RECT 49.255000 171.370000 50.335000 171.520000 ;
      RECT 49.255000 171.520000 50.185000 171.670000 ;
      RECT 49.255000 171.670000 50.035000 171.820000 ;
      RECT 49.255000 171.820000 49.885000 171.970000 ;
      RECT 49.255000 171.970000 49.735000 172.120000 ;
      RECT 49.255000 172.120000 49.585000 172.270000 ;
      RECT 49.255000 172.270000 49.435000 172.420000 ;
      RECT 49.255000 172.420000 49.285000 172.570000 ;
      RECT 49.255000 172.480000 49.375000 190.420000 ;
      RECT 49.290000   0.000000 49.990000  89.650000 ;
      RECT 49.290000   0.000000 50.090000  90.310000 ;
      RECT 49.290000  89.800000 49.440000  89.950000 ;
      RECT 49.290000  89.800000 49.440000  89.950000 ;
      RECT 49.290000  89.950000 49.590000  90.100000 ;
      RECT 49.290000  89.950000 49.590000  90.100000 ;
      RECT 49.290000  90.100000 49.740000  90.250000 ;
      RECT 49.290000  90.100000 49.740000  90.250000 ;
      RECT 49.290000  90.250000 49.890000  90.400000 ;
      RECT 49.290000  90.250000 49.890000  90.400000 ;
      RECT 49.290000  90.310000 55.765000  95.985000 ;
      RECT 49.290000  90.400000 50.040000  90.550000 ;
      RECT 49.290000  90.400000 50.040000  90.550000 ;
      RECT 49.290000  90.550000 50.190000  90.700000 ;
      RECT 49.290000  90.550000 50.190000  90.700000 ;
      RECT 49.290000  90.700000 50.340000  90.850000 ;
      RECT 49.290000  90.700000 50.340000  90.850000 ;
      RECT 49.290000  90.850000 50.490000  91.000000 ;
      RECT 49.290000  90.850000 50.490000  91.000000 ;
      RECT 49.290000  91.000000 50.640000  91.150000 ;
      RECT 49.290000  91.000000 50.640000  91.150000 ;
      RECT 49.290000  91.150000 50.790000  91.300000 ;
      RECT 49.290000  91.150000 50.790000  91.300000 ;
      RECT 49.290000  91.300000 50.940000  91.450000 ;
      RECT 49.290000  91.300000 50.940000  91.450000 ;
      RECT 49.290000  91.450000 51.090000  91.600000 ;
      RECT 49.290000  91.450000 51.090000  91.600000 ;
      RECT 49.290000  91.600000 51.240000  91.750000 ;
      RECT 49.290000  91.600000 51.240000  91.750000 ;
      RECT 49.290000  91.750000 51.390000  91.900000 ;
      RECT 49.290000  91.750000 51.390000  91.900000 ;
      RECT 49.290000  91.900000 51.540000  92.050000 ;
      RECT 49.290000  91.900000 51.540000  92.050000 ;
      RECT 49.290000  92.050000 51.690000  92.200000 ;
      RECT 49.290000  92.050000 51.690000  92.200000 ;
      RECT 49.290000  92.200000 51.840000  92.350000 ;
      RECT 49.290000  92.200000 51.840000  92.350000 ;
      RECT 49.290000  92.350000 51.990000  92.500000 ;
      RECT 49.290000  92.350000 51.990000  92.500000 ;
      RECT 49.290000  92.500000 52.140000  92.650000 ;
      RECT 49.290000  92.500000 52.140000  92.650000 ;
      RECT 49.290000  92.650000 52.290000  92.800000 ;
      RECT 49.290000  92.650000 52.290000  92.800000 ;
      RECT 49.290000  92.800000 52.440000  92.950000 ;
      RECT 49.290000  92.800000 52.440000  92.950000 ;
      RECT 49.290000  92.950000 52.590000  93.100000 ;
      RECT 49.290000  92.950000 52.590000  93.100000 ;
      RECT 49.290000  93.100000 52.740000  93.250000 ;
      RECT 49.290000  93.100000 52.740000  93.250000 ;
      RECT 49.290000  93.250000 52.890000  93.400000 ;
      RECT 49.290000  93.250000 52.890000  93.400000 ;
      RECT 49.290000  93.400000 53.040000  93.550000 ;
      RECT 49.290000  93.400000 53.040000  93.550000 ;
      RECT 49.290000  93.550000 53.190000  93.700000 ;
      RECT 49.290000  93.550000 53.190000  93.700000 ;
      RECT 49.290000  93.700000 53.340000  93.850000 ;
      RECT 49.290000  93.700000 53.340000  93.850000 ;
      RECT 49.290000  93.850000 53.490000  94.000000 ;
      RECT 49.290000  93.850000 53.490000  94.000000 ;
      RECT 49.290000  94.000000 53.640000  94.150000 ;
      RECT 49.290000  94.000000 53.640000  94.150000 ;
      RECT 49.290000  94.150000 53.790000  94.300000 ;
      RECT 49.290000  94.150000 53.790000  94.300000 ;
      RECT 49.290000  94.300000 53.940000  94.450000 ;
      RECT 49.290000  94.300000 53.940000  94.450000 ;
      RECT 49.290000  94.450000 54.090000  94.600000 ;
      RECT 49.290000  94.450000 54.090000  94.600000 ;
      RECT 49.290000  94.600000 54.240000  94.750000 ;
      RECT 49.290000  94.600000 54.240000  94.750000 ;
      RECT 49.290000  94.750000 54.390000  94.900000 ;
      RECT 49.290000  94.750000 54.390000  94.900000 ;
      RECT 49.290000  94.900000 54.540000  95.050000 ;
      RECT 49.290000  94.900000 54.540000  95.050000 ;
      RECT 49.290000  95.050000 54.690000  95.200000 ;
      RECT 49.290000  95.050000 54.690000  95.200000 ;
      RECT 49.290000  95.200000 54.840000  95.350000 ;
      RECT 49.290000  95.200000 54.840000  95.350000 ;
      RECT 49.290000  95.350000 54.990000  95.500000 ;
      RECT 49.290000  95.350000 54.990000  95.500000 ;
      RECT 49.290000  95.500000 55.140000  95.650000 ;
      RECT 49.290000  95.500000 55.140000  95.650000 ;
      RECT 49.290000  95.650000 55.290000  95.800000 ;
      RECT 49.290000  95.650000 55.290000  95.800000 ;
      RECT 49.290000  95.800000 55.440000  95.950000 ;
      RECT 49.290000  95.800000 55.440000  95.950000 ;
      RECT 49.290000  95.950000 55.590000  95.985000 ;
      RECT 49.290000  95.950000 55.590000  95.985000 ;
      RECT 49.290000  95.985000 57.915000  98.135000 ;
      RECT 49.440000  95.985000 55.625000  96.135000 ;
      RECT 49.440000  95.985000 55.625000  96.135000 ;
      RECT 49.590000  96.135000 55.775000  96.285000 ;
      RECT 49.590000  96.135000 55.775000  96.285000 ;
      RECT 49.740000  96.285000 55.925000  96.435000 ;
      RECT 49.740000  96.285000 55.925000  96.435000 ;
      RECT 49.890000  96.435000 56.075000  96.585000 ;
      RECT 49.890000  96.435000 56.075000  96.585000 ;
      RECT 50.040000  96.585000 56.225000  96.735000 ;
      RECT 50.040000  96.585000 56.225000  96.735000 ;
      RECT 50.190000  96.735000 56.375000  96.885000 ;
      RECT 50.190000  96.735000 56.375000  96.885000 ;
      RECT 50.340000  96.885000 56.525000  97.035000 ;
      RECT 50.340000  96.885000 56.525000  97.035000 ;
      RECT 50.490000  97.035000 56.675000  97.185000 ;
      RECT 50.490000  97.035000 56.675000  97.185000 ;
      RECT 50.640000  97.185000 56.825000  97.335000 ;
      RECT 50.640000  97.185000 56.825000  97.335000 ;
      RECT 50.790000  97.335000 56.975000  97.485000 ;
      RECT 50.790000  97.335000 56.975000  97.485000 ;
      RECT 50.940000  97.485000 57.125000  97.635000 ;
      RECT 50.940000  97.485000 57.125000  97.635000 ;
      RECT 51.090000  97.635000 57.275000  97.785000 ;
      RECT 51.090000  97.635000 57.275000  97.785000 ;
      RECT 51.240000  97.785000 57.425000  97.935000 ;
      RECT 51.240000  97.785000 57.425000  97.935000 ;
      RECT 51.390000  97.935000 57.575000  98.085000 ;
      RECT 51.390000  97.935000 57.575000  98.085000 ;
      RECT 51.440000  98.085000 57.725000  98.135000 ;
      RECT 51.440000  98.085000 57.725000  98.135000 ;
      RECT 51.440000  98.135000 57.775000  98.285000 ;
      RECT 51.440000  98.135000 57.775000  98.285000 ;
      RECT 51.440000  98.135000 59.330000  99.550000 ;
      RECT 51.440000  98.285000 57.925000  98.435000 ;
      RECT 51.440000  98.285000 57.925000  98.435000 ;
      RECT 51.440000  98.435000 58.075000  98.585000 ;
      RECT 51.440000  98.435000 58.075000  98.585000 ;
      RECT 51.440000  98.585000 58.225000  98.735000 ;
      RECT 51.440000  98.585000 58.225000  98.735000 ;
      RECT 51.440000  98.735000 58.375000  98.885000 ;
      RECT 51.440000  98.735000 58.375000  98.885000 ;
      RECT 51.440000  98.885000 58.525000  99.035000 ;
      RECT 51.440000  98.885000 58.525000  99.035000 ;
      RECT 51.440000  99.035000 58.675000  99.185000 ;
      RECT 51.440000  99.035000 58.675000  99.185000 ;
      RECT 51.440000  99.185000 58.825000  99.335000 ;
      RECT 51.440000  99.185000 58.825000  99.335000 ;
      RECT 51.440000  99.335000 58.975000  99.485000 ;
      RECT 51.440000  99.335000 58.975000  99.485000 ;
      RECT 51.440000  99.485000 59.125000  99.550000 ;
      RECT 51.440000  99.485000 59.125000  99.550000 ;
      RECT 51.440000  99.550000 61.200000 101.420000 ;
      RECT 51.590000  99.550000 59.190000  99.700000 ;
      RECT 51.590000  99.550000 59.190000  99.700000 ;
      RECT 51.740000  99.700000 59.340000  99.850000 ;
      RECT 51.740000  99.700000 59.340000  99.850000 ;
      RECT 51.890000  99.850000 59.490000 100.000000 ;
      RECT 51.890000  99.850000 59.490000 100.000000 ;
      RECT 52.040000 100.000000 59.640000 100.150000 ;
      RECT 52.040000 100.000000 59.640000 100.150000 ;
      RECT 52.190000 100.150000 59.790000 100.300000 ;
      RECT 52.190000 100.150000 59.790000 100.300000 ;
      RECT 52.340000 100.300000 59.940000 100.450000 ;
      RECT 52.340000 100.300000 59.940000 100.450000 ;
      RECT 52.490000 100.450000 60.090000 100.600000 ;
      RECT 52.490000 100.450000 60.090000 100.600000 ;
      RECT 52.640000 100.600000 60.240000 100.750000 ;
      RECT 52.640000 100.600000 60.240000 100.750000 ;
      RECT 52.790000 100.750000 60.390000 100.900000 ;
      RECT 52.790000 100.750000 60.390000 100.900000 ;
      RECT 52.940000 100.900000 60.540000 101.050000 ;
      RECT 52.940000 100.900000 60.540000 101.050000 ;
      RECT 53.090000 101.050000 60.690000 101.200000 ;
      RECT 53.090000 101.050000 60.690000 101.200000 ;
      RECT 53.240000 101.200000 60.840000 101.350000 ;
      RECT 53.240000 101.200000 60.840000 101.350000 ;
      RECT 53.310000 101.420000 61.200000 107.795000 ;
      RECT 53.350000 101.350000 60.990000 101.460000 ;
      RECT 53.350000 101.350000 60.990000 101.460000 ;
      RECT 53.500000 101.460000 61.100000 101.610000 ;
      RECT 53.500000 101.460000 61.100000 101.610000 ;
      RECT 53.650000 101.610000 61.100000 101.760000 ;
      RECT 53.650000 101.610000 61.100000 101.760000 ;
      RECT 53.800000 101.760000 61.100000 101.910000 ;
      RECT 53.800000 101.760000 61.100000 101.910000 ;
      RECT 53.950000 101.910000 61.100000 102.060000 ;
      RECT 53.950000 101.910000 61.100000 102.060000 ;
      RECT 54.100000 102.060000 61.100000 102.210000 ;
      RECT 54.100000 102.060000 61.100000 102.210000 ;
      RECT 54.250000 102.210000 61.100000 102.360000 ;
      RECT 54.250000 102.210000 61.100000 102.360000 ;
      RECT 54.400000 102.360000 61.100000 102.510000 ;
      RECT 54.400000 102.360000 61.100000 102.510000 ;
      RECT 54.550000 102.510000 61.100000 102.660000 ;
      RECT 54.550000 102.510000 61.100000 102.660000 ;
      RECT 54.700000 102.660000 61.100000 102.810000 ;
      RECT 54.700000 102.660000 61.100000 102.810000 ;
      RECT 54.850000 102.810000 61.100000 102.960000 ;
      RECT 54.850000 102.810000 61.100000 102.960000 ;
      RECT 55.000000 102.960000 61.100000 103.110000 ;
      RECT 55.000000 102.960000 61.100000 103.110000 ;
      RECT 55.150000 103.110000 61.100000 103.260000 ;
      RECT 55.150000 103.110000 61.100000 103.260000 ;
      RECT 55.300000 103.260000 61.100000 103.410000 ;
      RECT 55.300000 103.260000 61.100000 103.410000 ;
      RECT 55.450000 103.410000 61.100000 103.560000 ;
      RECT 55.450000 103.410000 61.100000 103.560000 ;
      RECT 55.600000 103.560000 61.100000 103.710000 ;
      RECT 55.600000 103.560000 61.100000 103.710000 ;
      RECT 55.750000 103.710000 61.100000 103.860000 ;
      RECT 55.750000 103.710000 61.100000 103.860000 ;
      RECT 55.900000 103.860000 61.100000 104.010000 ;
      RECT 55.900000 103.860000 61.100000 104.010000 ;
      RECT 56.050000 104.010000 61.100000 104.160000 ;
      RECT 56.050000 104.010000 61.100000 104.160000 ;
      RECT 56.200000 104.160000 61.100000 104.310000 ;
      RECT 56.200000 104.160000 61.100000 104.310000 ;
      RECT 56.350000 104.310000 61.100000 104.460000 ;
      RECT 56.350000 104.310000 61.100000 104.460000 ;
      RECT 56.500000 104.460000 61.100000 104.610000 ;
      RECT 56.500000 104.460000 61.100000 104.610000 ;
      RECT 56.650000 104.610000 61.100000 104.760000 ;
      RECT 56.650000 104.610000 61.100000 104.760000 ;
      RECT 56.800000 104.760000 61.100000 104.910000 ;
      RECT 56.800000 104.760000 61.100000 104.910000 ;
      RECT 56.950000 104.910000 61.100000 105.060000 ;
      RECT 56.950000 104.910000 61.100000 105.060000 ;
      RECT 57.100000 105.060000 61.100000 105.210000 ;
      RECT 57.100000 105.060000 61.100000 105.210000 ;
      RECT 57.250000 105.210000 61.100000 105.360000 ;
      RECT 57.250000 105.210000 61.100000 105.360000 ;
      RECT 57.400000 105.360000 61.100000 105.510000 ;
      RECT 57.400000 105.360000 61.100000 105.510000 ;
      RECT 57.550000 105.510000 61.100000 105.660000 ;
      RECT 57.550000 105.510000 61.100000 105.660000 ;
      RECT 57.700000 105.660000 61.100000 105.810000 ;
      RECT 57.700000 105.660000 61.100000 105.810000 ;
      RECT 57.850000 105.810000 61.100000 105.960000 ;
      RECT 57.850000 105.810000 61.100000 105.960000 ;
      RECT 58.000000 105.960000 61.100000 106.110000 ;
      RECT 58.000000 105.960000 61.100000 106.110000 ;
      RECT 58.150000 106.110000 61.100000 106.260000 ;
      RECT 58.150000 106.110000 61.100000 106.260000 ;
      RECT 58.300000 106.260000 61.100000 106.410000 ;
      RECT 58.300000 106.260000 61.100000 106.410000 ;
      RECT 58.450000 106.410000 61.100000 106.560000 ;
      RECT 58.450000 106.410000 61.100000 106.560000 ;
      RECT 58.600000 106.560000 61.100000 106.710000 ;
      RECT 58.600000 106.560000 61.100000 106.710000 ;
      RECT 58.750000 106.710000 61.100000 106.860000 ;
      RECT 58.750000 106.710000 61.100000 106.860000 ;
      RECT 58.900000 106.860000 61.100000 107.010000 ;
      RECT 58.900000 106.860000 61.100000 107.010000 ;
      RECT 59.050000 107.010000 61.100000 107.160000 ;
      RECT 59.050000 107.010000 61.100000 107.160000 ;
      RECT 59.200000 107.160000 61.100000 107.310000 ;
      RECT 59.200000 107.160000 61.100000 107.310000 ;
      RECT 59.350000 107.310000 61.100000 107.460000 ;
      RECT 59.350000 107.310000 61.100000 107.460000 ;
      RECT 59.500000 107.460000 61.100000 107.610000 ;
      RECT 59.500000 107.460000 61.100000 107.610000 ;
      RECT 59.650000 107.610000 61.100000 107.760000 ;
      RECT 59.650000 107.610000 61.100000 107.760000 ;
      RECT 59.685000 107.795000 61.200000 172.855000 ;
      RECT 59.685000 107.945000 59.835000 108.095000 ;
      RECT 59.685000 108.095000 59.985000 108.245000 ;
      RECT 59.685000 108.245000 60.135000 108.395000 ;
      RECT 59.685000 108.395000 60.285000 108.545000 ;
      RECT 59.685000 108.545000 60.435000 108.695000 ;
      RECT 59.685000 108.695000 60.585000 108.845000 ;
      RECT 59.685000 108.845000 60.735000 108.995000 ;
      RECT 59.685000 108.995000 60.885000 109.145000 ;
      RECT 59.685000 109.145000 61.035000 109.210000 ;
      RECT 59.685000 109.210000 61.100000 172.855000 ;
      RECT 59.685000 172.855000 61.200000 173.620000 ;
      RECT 59.800000 107.760000 61.100000 107.910000 ;
      RECT 59.800000 107.760000 61.100000 107.910000 ;
      RECT 59.835000 172.855000 61.100000 173.005000 ;
      RECT 59.950000 107.910000 61.100000 108.060000 ;
      RECT 59.950000 107.910000 61.100000 108.060000 ;
      RECT 59.985000 173.005000 61.100000 173.155000 ;
      RECT 60.100000 108.060000 61.100000 108.210000 ;
      RECT 60.100000 108.060000 61.100000 108.210000 ;
      RECT 60.135000 173.155000 61.100000 173.305000 ;
      RECT 60.250000 108.210000 61.100000 108.360000 ;
      RECT 60.250000 108.210000 61.100000 108.360000 ;
      RECT 60.285000 173.305000 61.100000 173.455000 ;
      RECT 60.400000 108.360000 61.100000 108.510000 ;
      RECT 60.400000 108.360000 61.100000 108.510000 ;
      RECT 60.435000 173.455000 61.100000 173.605000 ;
      RECT 60.450000 173.620000 75.000000 185.195000 ;
      RECT 60.550000 108.510000 61.100000 108.660000 ;
      RECT 60.550000 108.510000 61.100000 108.660000 ;
      RECT 60.550000 173.605000 61.100000 173.720000 ;
      RECT 60.700000 108.660000 61.100000 108.810000 ;
      RECT 60.700000 108.660000 61.100000 108.810000 ;
      RECT 60.700000 173.720000 75.000000 173.870000 ;
      RECT 60.700000 173.720000 75.000000 173.870000 ;
      RECT 60.850000 108.810000 61.100000 108.960000 ;
      RECT 60.850000 108.810000 61.100000 108.960000 ;
      RECT 60.850000 173.870000 75.000000 174.020000 ;
      RECT 60.850000 173.870000 75.000000 174.020000 ;
      RECT 61.000000 108.960000 61.100000 109.110000 ;
      RECT 61.000000 108.960000 61.100000 109.110000 ;
      RECT 61.000000 174.020000 75.000000 174.170000 ;
      RECT 61.000000 174.020000 75.000000 174.170000 ;
      RECT 61.150000 174.170000 75.000000 174.320000 ;
      RECT 61.150000 174.170000 75.000000 174.320000 ;
      RECT 61.300000 174.320000 75.000000 174.470000 ;
      RECT 61.300000 174.320000 75.000000 174.470000 ;
      RECT 61.450000 174.470000 75.000000 174.620000 ;
      RECT 61.450000 174.470000 75.000000 174.620000 ;
      RECT 61.600000 174.620000 75.000000 174.770000 ;
      RECT 61.600000 174.620000 75.000000 174.770000 ;
      RECT 61.750000 174.770000 75.000000 174.920000 ;
      RECT 61.750000 174.770000 75.000000 174.920000 ;
      RECT 61.900000 174.920000 75.000000 175.070000 ;
      RECT 61.900000 174.920000 75.000000 175.070000 ;
      RECT 62.050000 175.070000 75.000000 175.220000 ;
      RECT 62.050000 175.070000 75.000000 175.220000 ;
      RECT 62.200000 175.220000 75.000000 175.370000 ;
      RECT 62.200000 175.220000 75.000000 175.370000 ;
      RECT 62.350000 175.370000 75.000000 175.520000 ;
      RECT 62.350000 175.370000 75.000000 175.520000 ;
      RECT 62.500000 175.520000 75.000000 175.670000 ;
      RECT 62.500000 175.520000 75.000000 175.670000 ;
      RECT 62.650000 175.670000 75.000000 175.820000 ;
      RECT 62.650000 175.670000 75.000000 175.820000 ;
      RECT 62.800000 175.820000 75.000000 175.970000 ;
      RECT 62.800000 175.820000 75.000000 175.970000 ;
      RECT 62.950000 175.970000 75.000000 176.120000 ;
      RECT 62.950000 175.970000 75.000000 176.120000 ;
      RECT 63.100000 176.120000 75.000000 176.270000 ;
      RECT 63.100000 176.120000 75.000000 176.270000 ;
      RECT 63.250000 176.270000 75.000000 176.420000 ;
      RECT 63.250000 176.270000 75.000000 176.420000 ;
      RECT 63.400000 176.420000 75.000000 176.570000 ;
      RECT 63.400000 176.420000 75.000000 176.570000 ;
      RECT 63.550000 176.570000 75.000000 176.720000 ;
      RECT 63.550000 176.570000 75.000000 176.720000 ;
      RECT 63.700000 176.720000 75.000000 176.870000 ;
      RECT 63.700000 176.720000 75.000000 176.870000 ;
      RECT 63.850000 176.870000 75.000000 177.020000 ;
      RECT 63.850000 176.870000 75.000000 177.020000 ;
      RECT 64.000000 177.020000 75.000000 177.170000 ;
      RECT 64.000000 177.020000 75.000000 177.170000 ;
      RECT 64.150000 177.170000 75.000000 177.320000 ;
      RECT 64.150000 177.170000 75.000000 177.320000 ;
      RECT 64.300000 177.320000 75.000000 177.470000 ;
      RECT 64.300000 177.320000 75.000000 177.470000 ;
      RECT 64.450000 177.470000 75.000000 177.620000 ;
      RECT 64.450000 177.470000 75.000000 177.620000 ;
      RECT 64.600000 177.620000 75.000000 177.770000 ;
      RECT 64.600000 177.620000 75.000000 177.770000 ;
      RECT 64.750000 177.770000 75.000000 177.920000 ;
      RECT 64.750000 177.770000 75.000000 177.920000 ;
      RECT 64.900000 177.920000 75.000000 178.070000 ;
      RECT 64.900000 177.920000 75.000000 178.070000 ;
      RECT 65.050000 178.070000 75.000000 178.220000 ;
      RECT 65.050000 178.070000 75.000000 178.220000 ;
      RECT 65.200000 178.220000 75.000000 178.370000 ;
      RECT 65.200000 178.220000 75.000000 178.370000 ;
      RECT 65.350000 178.370000 75.000000 178.520000 ;
      RECT 65.350000 178.370000 75.000000 178.520000 ;
      RECT 65.500000 178.520000 75.000000 178.670000 ;
      RECT 65.500000 178.520000 75.000000 178.670000 ;
      RECT 65.650000 178.670000 75.000000 178.820000 ;
      RECT 65.650000 178.670000 75.000000 178.820000 ;
      RECT 65.800000 178.820000 75.000000 178.970000 ;
      RECT 65.800000 178.820000 75.000000 178.970000 ;
      RECT 65.950000 178.970000 75.000000 179.120000 ;
      RECT 65.950000 178.970000 75.000000 179.120000 ;
      RECT 66.100000 179.120000 75.000000 179.270000 ;
      RECT 66.100000 179.120000 75.000000 179.270000 ;
      RECT 66.250000 179.270000 75.000000 179.420000 ;
      RECT 66.250000 179.270000 75.000000 179.420000 ;
      RECT 66.400000 179.420000 75.000000 179.570000 ;
      RECT 66.400000 179.420000 75.000000 179.570000 ;
      RECT 66.550000 179.570000 75.000000 179.720000 ;
      RECT 66.550000 179.570000 75.000000 179.720000 ;
      RECT 66.700000 179.720000 75.000000 179.870000 ;
      RECT 66.700000 179.720000 75.000000 179.870000 ;
      RECT 66.850000 179.870000 75.000000 180.020000 ;
      RECT 66.850000 179.870000 75.000000 180.020000 ;
      RECT 67.000000 180.020000 75.000000 180.170000 ;
      RECT 67.000000 180.020000 75.000000 180.170000 ;
      RECT 67.150000 180.170000 75.000000 180.320000 ;
      RECT 67.150000 180.170000 75.000000 180.320000 ;
      RECT 67.300000 180.320000 75.000000 180.470000 ;
      RECT 67.300000 180.320000 75.000000 180.470000 ;
      RECT 67.450000 180.470000 75.000000 180.620000 ;
      RECT 67.450000 180.470000 75.000000 180.620000 ;
      RECT 67.600000 180.620000 75.000000 180.770000 ;
      RECT 67.600000 180.620000 75.000000 180.770000 ;
      RECT 67.750000 180.770000 75.000000 180.920000 ;
      RECT 67.750000 180.770000 75.000000 180.920000 ;
      RECT 67.900000 180.920000 75.000000 181.070000 ;
      RECT 67.900000 180.920000 75.000000 181.070000 ;
      RECT 68.050000 181.070000 75.000000 181.220000 ;
      RECT 68.050000 181.070000 75.000000 181.220000 ;
      RECT 68.200000 181.220000 75.000000 181.370000 ;
      RECT 68.200000 181.220000 75.000000 181.370000 ;
      RECT 68.350000 181.370000 75.000000 181.520000 ;
      RECT 68.350000 181.370000 75.000000 181.520000 ;
      RECT 68.500000 181.520000 75.000000 181.670000 ;
      RECT 68.500000 181.520000 75.000000 181.670000 ;
      RECT 68.650000 181.670000 75.000000 181.820000 ;
      RECT 68.650000 181.670000 75.000000 181.820000 ;
      RECT 68.800000 181.820000 75.000000 181.970000 ;
      RECT 68.800000 181.820000 75.000000 181.970000 ;
      RECT 68.950000 181.970000 75.000000 182.120000 ;
      RECT 68.950000 181.970000 75.000000 182.120000 ;
      RECT 69.100000 182.120000 75.000000 182.270000 ;
      RECT 69.100000 182.120000 75.000000 182.270000 ;
      RECT 69.250000 182.270000 75.000000 182.420000 ;
      RECT 69.250000 182.270000 75.000000 182.420000 ;
      RECT 69.400000 182.420000 75.000000 182.570000 ;
      RECT 69.400000 182.420000 75.000000 182.570000 ;
      RECT 69.550000 182.570000 75.000000 182.720000 ;
      RECT 69.550000 182.570000 75.000000 182.720000 ;
      RECT 69.700000 182.720000 75.000000 182.870000 ;
      RECT 69.700000 182.720000 75.000000 182.870000 ;
      RECT 69.850000 182.870000 75.000000 183.020000 ;
      RECT 69.850000 182.870000 75.000000 183.020000 ;
      RECT 70.000000 183.020000 75.000000 183.170000 ;
      RECT 70.000000 183.020000 75.000000 183.170000 ;
      RECT 70.150000 183.170000 75.000000 183.320000 ;
      RECT 70.150000 183.170000 75.000000 183.320000 ;
      RECT 70.300000 183.320000 75.000000 183.470000 ;
      RECT 70.300000 183.320000 75.000000 183.470000 ;
      RECT 70.450000 183.470000 75.000000 183.620000 ;
      RECT 70.450000 183.470000 75.000000 183.620000 ;
      RECT 70.600000 183.620000 75.000000 183.770000 ;
      RECT 70.600000 183.620000 75.000000 183.770000 ;
      RECT 70.750000 183.770000 75.000000 183.920000 ;
      RECT 70.750000 183.770000 75.000000 183.920000 ;
      RECT 70.900000 183.920000 75.000000 184.070000 ;
      RECT 70.900000 183.920000 75.000000 184.070000 ;
      RECT 71.050000 184.070000 75.000000 184.220000 ;
      RECT 71.050000 184.070000 75.000000 184.220000 ;
      RECT 71.200000 184.220000 75.000000 184.370000 ;
      RECT 71.200000 184.220000 75.000000 184.370000 ;
      RECT 71.350000 184.370000 75.000000 184.520000 ;
      RECT 71.350000 184.370000 75.000000 184.520000 ;
      RECT 71.500000 184.520000 75.000000 184.670000 ;
      RECT 71.500000 184.520000 75.000000 184.670000 ;
      RECT 71.650000 184.670000 75.000000 184.820000 ;
      RECT 71.650000 184.670000 75.000000 184.820000 ;
      RECT 71.800000 184.820000 75.000000 184.970000 ;
      RECT 71.800000 184.820000 75.000000 184.970000 ;
      RECT 71.950000 184.970000 75.000000 185.120000 ;
      RECT 71.950000 184.970000 75.000000 185.120000 ;
      RECT 72.025000 185.195000 75.000000 190.440000 ;
      RECT 72.025000 185.345000 72.175000 185.495000 ;
      RECT 72.025000 185.495000 72.325000 185.645000 ;
      RECT 72.025000 185.645000 72.475000 185.795000 ;
      RECT 72.025000 185.795000 72.625000 185.945000 ;
      RECT 72.025000 185.945000 72.775000 186.095000 ;
      RECT 72.025000 186.095000 72.925000 186.245000 ;
      RECT 72.025000 186.245000 73.075000 186.395000 ;
      RECT 72.025000 186.395000 73.225000 186.545000 ;
      RECT 72.025000 186.545000 73.375000 186.695000 ;
      RECT 72.025000 186.695000 73.525000 186.845000 ;
      RECT 72.025000 186.845000 73.675000 186.995000 ;
      RECT 72.025000 186.995000 73.825000 187.145000 ;
      RECT 72.025000 187.145000 73.975000 187.295000 ;
      RECT 72.025000 187.295000 74.125000 187.445000 ;
      RECT 72.025000 187.445000 74.275000 187.595000 ;
      RECT 72.025000 187.595000 74.425000 187.745000 ;
      RECT 72.025000 187.745000 74.575000 187.895000 ;
      RECT 72.025000 187.895000 74.725000 188.045000 ;
      RECT 72.025000 188.045000 74.875000 188.170000 ;
      RECT 72.025000 188.170000 75.000000 190.440000 ;
      RECT 72.100000 185.120000 75.000000 185.270000 ;
      RECT 72.100000 185.120000 75.000000 185.270000 ;
      RECT 72.250000 185.270000 75.000000 185.420000 ;
      RECT 72.250000 185.270000 75.000000 185.420000 ;
      RECT 72.400000 185.420000 75.000000 185.570000 ;
      RECT 72.400000 185.420000 75.000000 185.570000 ;
      RECT 72.550000 185.570000 75.000000 185.720000 ;
      RECT 72.550000 185.570000 75.000000 185.720000 ;
      RECT 72.700000 185.720000 75.000000 185.870000 ;
      RECT 72.700000 185.720000 75.000000 185.870000 ;
      RECT 72.850000 185.870000 75.000000 186.020000 ;
      RECT 72.850000 185.870000 75.000000 186.020000 ;
      RECT 73.000000 186.020000 75.000000 186.170000 ;
      RECT 73.000000 186.020000 75.000000 186.170000 ;
      RECT 73.150000 186.170000 75.000000 186.320000 ;
      RECT 73.150000 186.170000 75.000000 186.320000 ;
      RECT 73.300000 186.320000 75.000000 186.470000 ;
      RECT 73.300000 186.320000 75.000000 186.470000 ;
      RECT 73.450000 186.470000 75.000000 186.620000 ;
      RECT 73.450000 186.470000 75.000000 186.620000 ;
      RECT 73.600000 186.620000 75.000000 186.770000 ;
      RECT 73.600000 186.620000 75.000000 186.770000 ;
      RECT 73.750000 186.770000 75.000000 186.920000 ;
      RECT 73.750000 186.770000 75.000000 186.920000 ;
      RECT 73.900000 186.920000 75.000000 187.070000 ;
      RECT 73.900000 186.920000 75.000000 187.070000 ;
      RECT 74.050000 187.070000 75.000000 187.220000 ;
      RECT 74.050000 187.070000 75.000000 187.220000 ;
      RECT 74.200000 187.220000 75.000000 187.370000 ;
      RECT 74.200000 187.220000 75.000000 187.370000 ;
      RECT 74.350000 187.370000 75.000000 187.520000 ;
      RECT 74.350000 187.370000 75.000000 187.520000 ;
      RECT 74.500000 187.520000 75.000000 187.670000 ;
      RECT 74.500000 187.520000 75.000000 187.670000 ;
      RECT 74.590000   0.000000 75.000000 173.620000 ;
      RECT 74.650000 187.670000 75.000000 187.820000 ;
      RECT 74.650000 187.670000 75.000000 187.820000 ;
      RECT 74.690000   0.000000 75.000000 173.720000 ;
      RECT 74.800000 187.820000 75.000000 187.970000 ;
      RECT 74.800000 187.820000 75.000000 187.970000 ;
      RECT 74.950000 187.970000 75.000000 188.120000 ;
      RECT 74.950000 187.970000 75.000000 188.120000 ;
    LAYER met4 ;
      RECT  4.800000 104.380000  5.160000 104.530000 ;
      RECT  4.800000 104.530000  5.525000 104.680000 ;
      RECT  4.800000 104.680000  5.885000 104.830000 ;
      RECT  4.800000 104.830000  6.245000 104.980000 ;
      RECT  4.800000 104.980000  6.610000 105.130000 ;
      RECT  4.800000 105.130000  6.970000 105.280000 ;
      RECT  4.800000 105.280000  7.330000 105.350000 ;
      RECT  4.800000 105.350000  7.500000 165.450000 ;
      RECT  4.800000 165.450000  7.500000 165.600000 ;
      RECT  4.800000 165.600000  7.650000 165.750000 ;
      RECT  4.800000 165.750000  7.800000 165.900000 ;
      RECT  4.800000 165.900000  7.950000 166.050000 ;
      RECT  4.800000 166.050000  8.100000 166.200000 ;
      RECT  4.800000 166.200000  8.250000 166.350000 ;
      RECT  4.800000 166.350000  8.400000 166.500000 ;
      RECT  4.800000 166.500000  8.550000 166.570000 ;
      RECT  4.840000 104.265000  7.460000 165.545000 ;
      RECT  4.880000 104.150000  8.620000 104.230000 ;
      RECT  4.950000 166.570000  8.620000 166.720000 ;
      RECT  5.030000 104.000000  8.700000 104.150000 ;
      RECT  5.100000 166.720000  8.770000 166.870000 ;
      RECT  5.160000 104.230000  8.470000 104.380000 ;
      RECT  5.180000 103.850000  8.850000 104.000000 ;
      RECT  5.250000 166.870000  8.920000 167.020000 ;
      RECT  5.330000 103.700000  9.000000 103.850000 ;
      RECT  5.400000 167.020000  9.070000 167.170000 ;
      RECT  5.470000 165.675000  7.595000 167.175000 ;
      RECT  5.480000 103.550000  9.150000 103.700000 ;
      RECT  5.525000 104.380000  8.320000 104.530000 ;
      RECT  5.550000 167.170000  9.220000 167.320000 ;
      RECT  5.630000 103.400000  9.300000 103.550000 ;
      RECT  5.655000 103.425000  6.280000 104.075000 ;
      RECT  5.700000 167.320000  9.370000 167.470000 ;
      RECT  5.780000 103.250000  9.450000 103.400000 ;
      RECT  5.850000 167.470000  9.520000 167.620000 ;
      RECT  5.885000 104.530000  8.170000 104.680000 ;
      RECT  5.930000 103.100000  9.600000 103.250000 ;
      RECT  6.000000 167.620000  9.670000 167.770000 ;
      RECT  6.080000 102.950000  9.750000 103.100000 ;
      RECT  6.150000 167.770000  9.820000 167.920000 ;
      RECT  6.230000 102.800000  9.900000 102.950000 ;
      RECT  6.235000 167.300000  6.860000 167.950000 ;
      RECT  6.245000 104.680000  8.020000 104.830000 ;
      RECT  6.300000 167.920000  9.970000 168.070000 ;
      RECT  6.380000 102.650000 10.050000 102.800000 ;
      RECT  6.450000 168.070000 10.120000 168.220000 ;
      RECT  6.510000 102.630000  8.635000 104.130000 ;
      RECT  6.530000 102.500000 10.200000 102.650000 ;
      RECT  6.600000 168.220000 10.270000 168.370000 ;
      RECT  6.610000 104.830000  7.870000 104.980000 ;
      RECT  6.680000 102.350000 10.350000 102.500000 ;
      RECT  6.750000 168.370000 10.420000 168.520000 ;
      RECT  6.830000 102.200000 10.500000 102.350000 ;
      RECT  6.900000 168.520000 10.570000 168.670000 ;
      RECT  6.970000 104.980000  7.720000 105.130000 ;
      RECT  6.980000 102.050000 10.650000 102.200000 ;
      RECT  7.050000 168.670000 10.720000 168.820000 ;
      RECT  7.070000 167.275000  9.195000 168.775000 ;
      RECT  7.130000 101.900000 10.800000 102.050000 ;
      RECT  7.200000 168.820000 10.870000 168.970000 ;
      RECT  7.275000 101.855000  7.900000 102.505000 ;
      RECT  7.280000 101.750000 10.950000 101.900000 ;
      RECT  7.310000 104.205000  7.935000 104.855000 ;
      RECT  7.330000 105.130000  7.570000 105.280000 ;
      RECT  7.350000 168.970000 11.020000 169.120000 ;
      RECT  7.430000 101.600000 11.100000 101.750000 ;
      RECT  7.500000 169.120000 11.170000 169.270000 ;
      RECT  7.580000 101.450000 11.250000 101.600000 ;
      RECT  7.650000 169.270000 11.320000 169.420000 ;
      RECT  7.675000 166.490000  8.300000 167.140000 ;
      RECT  7.730000 101.300000 11.400000 101.450000 ;
      RECT  7.800000 169.420000 11.470000 169.570000 ;
      RECT  7.875000 168.940000  8.500000 169.590000 ;
      RECT  7.880000 101.150000 11.550000 101.300000 ;
      RECT  7.950000 169.570000 11.620000 169.720000 ;
      RECT  8.030000 101.000000 11.700000 101.150000 ;
      RECT  8.100000 169.720000 11.770000 169.870000 ;
      RECT  8.110000 101.030000 10.235000 102.530000 ;
      RECT  8.180000 100.850000 11.850000 101.000000 ;
      RECT  8.250000 169.870000 11.920000 170.020000 ;
      RECT  8.330000 100.700000 12.000000 100.850000 ;
      RECT  8.400000 170.020000 12.070000 170.170000 ;
      RECT  8.480000 100.550000 12.150000 100.700000 ;
      RECT  8.550000 170.170000 12.220000 170.320000 ;
      RECT  8.630000 100.400000 12.300000 100.550000 ;
      RECT  8.630000 170.320000 12.370000 170.400000 ;
      RECT  8.690000 168.895000 10.815000 170.395000 ;
      RECT  8.715000 102.665000  9.340000 103.315000 ;
      RECT  8.780000 100.250000 62.550000 100.400000 ;
      RECT  8.780000 170.400000 12.390000 170.550000 ;
      RECT  8.915000 100.215000  9.540000 100.865000 ;
      RECT  8.930000 100.100000 62.610000 100.250000 ;
      RECT  8.930000 170.550000 12.325000 170.700000 ;
      RECT  9.080000  99.950000 62.675000 100.100000 ;
      RECT  9.080000 170.700000 12.265000 170.850000 ;
      RECT  9.230000  99.800000 62.735000  99.950000 ;
      RECT  9.230000 170.850000 12.200000 171.000000 ;
      RECT  9.300000 168.115000  9.925000 168.765000 ;
      RECT  9.320000 170.425000  9.730000 171.075000 ;
      RECT  9.380000  99.650000 62.800000  99.800000 ;
      RECT  9.380000 171.000000 12.140000 171.150000 ;
      RECT  9.530000  99.500000 62.860000  99.650000 ;
      RECT  9.530000 171.150000 12.075000 171.300000 ;
      RECT  9.680000  99.350000 62.925000  99.500000 ;
      RECT  9.680000 171.300000 12.015000 171.450000 ;
      RECT  9.730000  99.410000 11.855000 100.910000 ;
      RECT  9.830000  99.200000 62.985000  99.350000 ;
      RECT  9.830000 171.450000 11.950000 171.600000 ;
      RECT  9.965000 170.770000 11.105000 171.580000 ;
      RECT  9.980000  99.050000 63.050000  99.200000 ;
      RECT  9.980000 171.600000 11.890000 171.750000 ;
      RECT 10.130000  98.900000 63.110000  99.050000 ;
      RECT 10.130000 171.750000 11.830000 171.900000 ;
      RECT 10.280000  98.750000 63.170000  98.900000 ;
      RECT 10.280000 171.900000 11.765000 172.050000 ;
      RECT 10.340000 101.040000 10.965000 101.690000 ;
      RECT 10.430000  98.600000 63.235000  98.750000 ;
      RECT 10.430000 172.050000 11.705000 172.200000 ;
      RECT 10.580000  98.450000 63.295000  98.600000 ;
      RECT 10.580000 172.200000 11.640000 172.350000 ;
      RECT 10.610000 171.715000 11.020000 172.365000 ;
      RECT 10.620000  98.510000 11.245000  99.160000 ;
      RECT 10.730000  98.300000 63.360000  98.450000 ;
      RECT 10.730000 172.350000 11.580000 172.500000 ;
      RECT 10.880000  98.150000 63.420000  98.300000 ;
      RECT 10.880000 172.500000 11.515000 172.650000 ;
      RECT 10.890000 169.555000 11.515000 170.205000 ;
      RECT 11.030000  98.000000 63.485000  98.150000 ;
      RECT 11.030000 172.650000 11.455000 172.800000 ;
      RECT 11.180000  97.850000 63.545000  98.000000 ;
      RECT 11.180000 172.800000 11.390000 172.950000 ;
      RECT 11.330000  97.700000 63.610000  97.850000 ;
      RECT 11.330000 170.400000 13.335000 173.100000 ;
      RECT 11.390000 172.950000 63.670000 173.100000 ;
      RECT 11.455000 172.800000 63.820000 172.950000 ;
      RECT 11.515000 172.650000 63.970000 172.800000 ;
      RECT 11.580000 172.500000 64.120000 172.650000 ;
      RECT 11.640000 172.350000 64.270000 172.500000 ;
      RECT 11.705000 172.200000 64.420000 172.350000 ;
      RECT 11.765000 172.050000 64.570000 172.200000 ;
      RECT 11.830000 171.900000 64.720000 172.050000 ;
      RECT 11.890000 171.750000 64.870000 171.900000 ;
      RECT 11.950000 171.600000 65.020000 171.750000 ;
      RECT 12.015000 171.450000 65.170000 171.600000 ;
      RECT 12.075000 171.300000 65.320000 171.450000 ;
      RECT 12.140000 171.150000 65.470000 171.300000 ;
      RECT 12.200000 171.000000 65.620000 171.150000 ;
      RECT 12.265000 170.850000 65.770000 171.000000 ;
      RECT 12.325000 170.700000 65.920000 170.850000 ;
      RECT 12.390000 170.550000 66.070000 170.700000 ;
      RECT 12.450000 170.400000 66.220000 170.550000 ;
      RECT 58.800000  97.740000 59.420000  98.535000 ;
      RECT 59.465000  97.725000 63.575000  99.225000 ;
      RECT 60.180000  99.285000 60.630000  99.935000 ;
      RECT 60.700000  99.420000 62.760000 100.350000 ;
      RECT 61.655000 170.400000 63.665000 173.100000 ;
      RECT 62.610000 100.250000 66.220000 100.400000 ;
      RECT 62.630000 170.320000 66.370000 170.400000 ;
      RECT 62.675000 100.100000 66.070000 100.250000 ;
      RECT 62.700000 100.400000 66.370000 100.550000 ;
      RECT 62.735000  99.950000 65.920000 100.100000 ;
      RECT 62.780000 170.170000 66.450000 170.320000 ;
      RECT 62.800000  99.800000 65.770000  99.950000 ;
      RECT 62.850000 100.550000 66.520000 100.700000 ;
      RECT 62.860000  99.650000 65.620000  99.800000 ;
      RECT 62.925000  99.500000 65.470000  99.650000 ;
      RECT 62.930000 170.020000 66.600000 170.170000 ;
      RECT 62.985000  99.350000 65.320000  99.500000 ;
      RECT 63.000000 100.700000 66.670000 100.850000 ;
      RECT 63.050000  99.200000 65.170000  99.350000 ;
      RECT 63.080000 169.870000 66.750000 170.020000 ;
      RECT 63.110000  99.050000 65.020000  99.200000 ;
      RECT 63.135000  99.410000 65.260000 100.910000 ;
      RECT 63.150000 100.850000 66.820000 101.000000 ;
      RECT 63.170000  98.900000 64.870000  99.050000 ;
      RECT 63.230000 169.720000 66.900000 169.870000 ;
      RECT 63.235000  98.750000 64.720000  98.900000 ;
      RECT 63.295000  98.600000 64.570000  98.750000 ;
      RECT 63.300000 101.000000 66.970000 101.150000 ;
      RECT 63.360000  98.450000 64.420000  98.600000 ;
      RECT 63.380000 169.570000 67.050000 169.720000 ;
      RECT 63.420000  98.300000 64.270000  98.450000 ;
      RECT 63.450000 101.150000 67.120000 101.300000 ;
      RECT 63.475000 169.555000 64.100000 170.205000 ;
      RECT 63.485000  98.150000 64.120000  98.300000 ;
      RECT 63.530000 169.420000 67.200000 169.570000 ;
      RECT 63.545000  98.000000 63.970000  98.150000 ;
      RECT 63.600000 101.300000 67.270000 101.450000 ;
      RECT 63.610000  97.850000 63.820000  98.000000 ;
      RECT 63.680000 169.270000 67.350000 169.420000 ;
      RECT 63.745000  98.510000 64.370000  99.160000 ;
      RECT 63.750000 101.450000 67.420000 101.600000 ;
      RECT 63.830000 169.120000 67.500000 169.270000 ;
      RECT 63.885000 170.770000 65.025000 171.580000 ;
      RECT 63.900000 101.600000 67.570000 101.750000 ;
      RECT 63.970000 171.715000 64.380000 172.365000 ;
      RECT 63.980000 168.970000 67.650000 169.120000 ;
      RECT 64.025000 101.040000 64.650000 101.690000 ;
      RECT 64.050000 101.750000 67.720000 101.900000 ;
      RECT 64.130000 168.820000 67.800000 168.970000 ;
      RECT 64.175000 168.895000 66.300000 170.395000 ;
      RECT 64.200000 101.900000 67.870000 102.050000 ;
      RECT 64.280000 168.670000 67.950000 168.820000 ;
      RECT 64.350000 102.050000 68.020000 102.200000 ;
      RECT 64.430000 168.520000 68.100000 168.670000 ;
      RECT 64.500000 102.200000 68.170000 102.350000 ;
      RECT 64.580000 168.370000 68.250000 168.520000 ;
      RECT 64.650000 102.350000 68.320000 102.500000 ;
      RECT 64.730000 168.220000 68.400000 168.370000 ;
      RECT 64.755000 101.030000 66.880000 102.530000 ;
      RECT 64.800000 102.500000 68.470000 102.650000 ;
      RECT 64.880000 168.070000 68.550000 168.220000 ;
      RECT 64.950000 102.650000 68.620000 102.800000 ;
      RECT 65.030000 167.920000 68.700000 168.070000 ;
      RECT 65.065000 168.115000 65.690000 168.765000 ;
      RECT 65.100000 102.800000 68.770000 102.950000 ;
      RECT 65.180000 167.770000 68.850000 167.920000 ;
      RECT 65.250000 102.950000 68.920000 103.100000 ;
      RECT 65.260000 170.425000 65.670000 171.075000 ;
      RECT 65.330000 167.620000 69.000000 167.770000 ;
      RECT 65.400000 103.100000 69.070000 103.250000 ;
      RECT 65.450000 100.215000 66.075000 100.865000 ;
      RECT 65.480000 167.470000 69.150000 167.620000 ;
      RECT 65.550000 103.250000 69.220000 103.400000 ;
      RECT 65.630000 167.320000 69.300000 167.470000 ;
      RECT 65.650000 102.665000 66.275000 103.315000 ;
      RECT 65.700000 103.400000 69.370000 103.550000 ;
      RECT 65.780000 167.170000 69.450000 167.320000 ;
      RECT 65.795000 167.275000 67.920000 168.775000 ;
      RECT 65.850000 103.550000 69.520000 103.700000 ;
      RECT 65.930000 167.020000 69.600000 167.170000 ;
      RECT 66.000000 103.700000 69.670000 103.850000 ;
      RECT 66.080000 166.870000 69.750000 167.020000 ;
      RECT 66.150000 103.850000 69.820000 104.000000 ;
      RECT 66.230000 166.720000 69.900000 166.870000 ;
      RECT 66.300000 104.000000 69.970000 104.150000 ;
      RECT 66.355000 102.630000 68.480000 104.130000 ;
      RECT 66.380000 104.150000 70.120000 104.230000 ;
      RECT 66.380000 166.570000 70.050000 166.720000 ;
      RECT 66.450000 166.500000 70.030000 166.570000 ;
      RECT 66.490000 168.940000 67.115000 169.590000 ;
      RECT 66.530000 104.230000 70.200000 104.380000 ;
      RECT 66.600000 166.350000 69.670000 166.500000 ;
      RECT 66.680000 104.380000 70.200000 104.530000 ;
      RECT 66.690000 166.490000 67.315000 167.140000 ;
      RECT 66.750000 166.200000 69.310000 166.350000 ;
      RECT 66.830000 104.530000 70.200000 104.680000 ;
      RECT 66.900000 166.050000 68.945000 166.200000 ;
      RECT 66.980000 104.680000 70.200000 104.830000 ;
      RECT 67.050000 165.900000 68.585000 166.050000 ;
      RECT 67.055000 104.205000 67.680000 104.855000 ;
      RECT 67.090000 101.855000 67.715000 102.505000 ;
      RECT 67.130000 104.830000 70.200000 104.980000 ;
      RECT 67.200000 165.750000 68.225000 165.900000 ;
      RECT 67.280000 104.980000 70.200000 105.130000 ;
      RECT 67.350000 165.600000 67.860000 165.750000 ;
      RECT 67.395000 165.675000 69.520000 167.175000 ;
      RECT 67.430000 105.130000 70.200000 105.280000 ;
      RECT 67.500000 105.280000 70.200000 105.350000 ;
      RECT 67.500000 105.350000 70.200000 165.450000 ;
      RECT 67.530000 104.265000 70.150000 165.545000 ;
      RECT 67.860000 165.450000 70.200000 165.600000 ;
      RECT 68.130000 167.300000 68.755000 167.950000 ;
      RECT 68.225000 165.600000 70.200000 165.750000 ;
      RECT 68.550000 103.230000 69.170000 104.115000 ;
      RECT 68.585000 165.750000 70.200000 165.900000 ;
      RECT 68.945000 165.900000 70.200000 166.050000 ;
      RECT 69.200000 103.590000 69.535000 104.240000 ;
      RECT 69.310000 166.050000 70.200000 166.200000 ;
      RECT 69.670000 166.200000 70.200000 166.350000 ;
      RECT 70.030000 166.350000 70.200000 166.500000 ;
  END
END sky130_fd_io__top_power_hvc_wpad


MACRO sky130_fd_io__overlay_vssa_lvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.500000 34.740000 24.400000 38.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500000 49.650000 24.400000 50.820000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 34.740000 74.655000 38.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 49.650000 74.655000 50.820000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 24.375000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 24.375000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.590000 34.820000  0.790000 35.020000 ;
        RECT  0.590000 35.260000  0.790000 35.460000 ;
        RECT  0.590000 35.700000  0.790000 35.900000 ;
        RECT  0.590000 36.140000  0.790000 36.340000 ;
        RECT  0.590000 36.580000  0.790000 36.780000 ;
        RECT  0.590000 37.020000  0.790000 37.220000 ;
        RECT  0.590000 37.460000  0.790000 37.660000 ;
        RECT  0.590000 37.900000  0.790000 38.100000 ;
        RECT  0.590000 49.715000  0.790000 49.915000 ;
        RECT  0.590000 50.135000  0.790000 50.335000 ;
        RECT  0.590000 50.555000  0.790000 50.755000 ;
        RECT  1.000000 34.820000  1.200000 35.020000 ;
        RECT  1.000000 35.260000  1.200000 35.460000 ;
        RECT  1.000000 35.700000  1.200000 35.900000 ;
        RECT  1.000000 36.140000  1.200000 36.340000 ;
        RECT  1.000000 36.580000  1.200000 36.780000 ;
        RECT  1.000000 37.020000  1.200000 37.220000 ;
        RECT  1.000000 37.460000  1.200000 37.660000 ;
        RECT  1.000000 37.900000  1.200000 38.100000 ;
        RECT  1.000000 49.715000  1.200000 49.915000 ;
        RECT  1.000000 50.135000  1.200000 50.335000 ;
        RECT  1.000000 50.555000  1.200000 50.755000 ;
        RECT  1.410000 34.820000  1.610000 35.020000 ;
        RECT  1.410000 35.260000  1.610000 35.460000 ;
        RECT  1.410000 35.700000  1.610000 35.900000 ;
        RECT  1.410000 36.140000  1.610000 36.340000 ;
        RECT  1.410000 36.580000  1.610000 36.780000 ;
        RECT  1.410000 37.020000  1.610000 37.220000 ;
        RECT  1.410000 37.460000  1.610000 37.660000 ;
        RECT  1.410000 37.900000  1.610000 38.100000 ;
        RECT  1.410000 49.715000  1.610000 49.915000 ;
        RECT  1.410000 50.135000  1.610000 50.335000 ;
        RECT  1.410000 50.555000  1.610000 50.755000 ;
        RECT  1.820000 34.820000  2.020000 35.020000 ;
        RECT  1.820000 35.260000  2.020000 35.460000 ;
        RECT  1.820000 35.700000  2.020000 35.900000 ;
        RECT  1.820000 36.140000  2.020000 36.340000 ;
        RECT  1.820000 36.580000  2.020000 36.780000 ;
        RECT  1.820000 37.020000  2.020000 37.220000 ;
        RECT  1.820000 37.460000  2.020000 37.660000 ;
        RECT  1.820000 37.900000  2.020000 38.100000 ;
        RECT  1.820000 49.715000  2.020000 49.915000 ;
        RECT  1.820000 50.135000  2.020000 50.335000 ;
        RECT  1.820000 50.555000  2.020000 50.755000 ;
        RECT  2.230000 34.820000  2.430000 35.020000 ;
        RECT  2.230000 35.260000  2.430000 35.460000 ;
        RECT  2.230000 35.700000  2.430000 35.900000 ;
        RECT  2.230000 36.140000  2.430000 36.340000 ;
        RECT  2.230000 36.580000  2.430000 36.780000 ;
        RECT  2.230000 37.020000  2.430000 37.220000 ;
        RECT  2.230000 37.460000  2.430000 37.660000 ;
        RECT  2.230000 37.900000  2.430000 38.100000 ;
        RECT  2.230000 49.715000  2.430000 49.915000 ;
        RECT  2.230000 50.135000  2.430000 50.335000 ;
        RECT  2.230000 50.555000  2.430000 50.755000 ;
        RECT  2.640000 34.820000  2.840000 35.020000 ;
        RECT  2.640000 35.260000  2.840000 35.460000 ;
        RECT  2.640000 35.700000  2.840000 35.900000 ;
        RECT  2.640000 36.140000  2.840000 36.340000 ;
        RECT  2.640000 36.580000  2.840000 36.780000 ;
        RECT  2.640000 37.020000  2.840000 37.220000 ;
        RECT  2.640000 37.460000  2.840000 37.660000 ;
        RECT  2.640000 37.900000  2.840000 38.100000 ;
        RECT  2.640000 49.715000  2.840000 49.915000 ;
        RECT  2.640000 50.135000  2.840000 50.335000 ;
        RECT  2.640000 50.555000  2.840000 50.755000 ;
        RECT  3.050000 34.820000  3.250000 35.020000 ;
        RECT  3.050000 35.260000  3.250000 35.460000 ;
        RECT  3.050000 35.700000  3.250000 35.900000 ;
        RECT  3.050000 36.140000  3.250000 36.340000 ;
        RECT  3.050000 36.580000  3.250000 36.780000 ;
        RECT  3.050000 37.020000  3.250000 37.220000 ;
        RECT  3.050000 37.460000  3.250000 37.660000 ;
        RECT  3.050000 37.900000  3.250000 38.100000 ;
        RECT  3.050000 49.715000  3.250000 49.915000 ;
        RECT  3.050000 50.135000  3.250000 50.335000 ;
        RECT  3.050000 50.555000  3.250000 50.755000 ;
        RECT  3.455000 34.820000  3.655000 35.020000 ;
        RECT  3.455000 35.260000  3.655000 35.460000 ;
        RECT  3.455000 35.700000  3.655000 35.900000 ;
        RECT  3.455000 36.140000  3.655000 36.340000 ;
        RECT  3.455000 36.580000  3.655000 36.780000 ;
        RECT  3.455000 37.020000  3.655000 37.220000 ;
        RECT  3.455000 37.460000  3.655000 37.660000 ;
        RECT  3.455000 37.900000  3.655000 38.100000 ;
        RECT  3.455000 49.715000  3.655000 49.915000 ;
        RECT  3.455000 50.135000  3.655000 50.335000 ;
        RECT  3.455000 50.555000  3.655000 50.755000 ;
        RECT  3.860000 34.820000  4.060000 35.020000 ;
        RECT  3.860000 35.260000  4.060000 35.460000 ;
        RECT  3.860000 35.700000  4.060000 35.900000 ;
        RECT  3.860000 36.140000  4.060000 36.340000 ;
        RECT  3.860000 36.580000  4.060000 36.780000 ;
        RECT  3.860000 37.020000  4.060000 37.220000 ;
        RECT  3.860000 37.460000  4.060000 37.660000 ;
        RECT  3.860000 37.900000  4.060000 38.100000 ;
        RECT  3.860000 49.715000  4.060000 49.915000 ;
        RECT  3.860000 50.135000  4.060000 50.335000 ;
        RECT  3.860000 50.555000  4.060000 50.755000 ;
        RECT  4.265000 34.820000  4.465000 35.020000 ;
        RECT  4.265000 35.260000  4.465000 35.460000 ;
        RECT  4.265000 35.700000  4.465000 35.900000 ;
        RECT  4.265000 36.140000  4.465000 36.340000 ;
        RECT  4.265000 36.580000  4.465000 36.780000 ;
        RECT  4.265000 37.020000  4.465000 37.220000 ;
        RECT  4.265000 37.460000  4.465000 37.660000 ;
        RECT  4.265000 37.900000  4.465000 38.100000 ;
        RECT  4.265000 49.715000  4.465000 49.915000 ;
        RECT  4.265000 50.135000  4.465000 50.335000 ;
        RECT  4.265000 50.555000  4.465000 50.755000 ;
        RECT  4.670000 34.820000  4.870000 35.020000 ;
        RECT  4.670000 35.260000  4.870000 35.460000 ;
        RECT  4.670000 35.700000  4.870000 35.900000 ;
        RECT  4.670000 36.140000  4.870000 36.340000 ;
        RECT  4.670000 36.580000  4.870000 36.780000 ;
        RECT  4.670000 37.020000  4.870000 37.220000 ;
        RECT  4.670000 37.460000  4.870000 37.660000 ;
        RECT  4.670000 37.900000  4.870000 38.100000 ;
        RECT  4.670000 49.715000  4.870000 49.915000 ;
        RECT  4.670000 50.135000  4.870000 50.335000 ;
        RECT  4.670000 50.555000  4.870000 50.755000 ;
        RECT  5.075000 34.820000  5.275000 35.020000 ;
        RECT  5.075000 35.260000  5.275000 35.460000 ;
        RECT  5.075000 35.700000  5.275000 35.900000 ;
        RECT  5.075000 36.140000  5.275000 36.340000 ;
        RECT  5.075000 36.580000  5.275000 36.780000 ;
        RECT  5.075000 37.020000  5.275000 37.220000 ;
        RECT  5.075000 37.460000  5.275000 37.660000 ;
        RECT  5.075000 37.900000  5.275000 38.100000 ;
        RECT  5.075000 49.715000  5.275000 49.915000 ;
        RECT  5.075000 50.135000  5.275000 50.335000 ;
        RECT  5.075000 50.555000  5.275000 50.755000 ;
        RECT  5.480000 34.820000  5.680000 35.020000 ;
        RECT  5.480000 35.260000  5.680000 35.460000 ;
        RECT  5.480000 35.700000  5.680000 35.900000 ;
        RECT  5.480000 36.140000  5.680000 36.340000 ;
        RECT  5.480000 36.580000  5.680000 36.780000 ;
        RECT  5.480000 37.020000  5.680000 37.220000 ;
        RECT  5.480000 37.460000  5.680000 37.660000 ;
        RECT  5.480000 37.900000  5.680000 38.100000 ;
        RECT  5.480000 49.715000  5.680000 49.915000 ;
        RECT  5.480000 50.135000  5.680000 50.335000 ;
        RECT  5.480000 50.555000  5.680000 50.755000 ;
        RECT  5.885000 34.820000  6.085000 35.020000 ;
        RECT  5.885000 35.260000  6.085000 35.460000 ;
        RECT  5.885000 35.700000  6.085000 35.900000 ;
        RECT  5.885000 36.140000  6.085000 36.340000 ;
        RECT  5.885000 36.580000  6.085000 36.780000 ;
        RECT  5.885000 37.020000  6.085000 37.220000 ;
        RECT  5.885000 37.460000  6.085000 37.660000 ;
        RECT  5.885000 37.900000  6.085000 38.100000 ;
        RECT  5.885000 49.715000  6.085000 49.915000 ;
        RECT  5.885000 50.135000  6.085000 50.335000 ;
        RECT  5.885000 50.555000  6.085000 50.755000 ;
        RECT  6.290000 34.820000  6.490000 35.020000 ;
        RECT  6.290000 35.260000  6.490000 35.460000 ;
        RECT  6.290000 35.700000  6.490000 35.900000 ;
        RECT  6.290000 36.140000  6.490000 36.340000 ;
        RECT  6.290000 36.580000  6.490000 36.780000 ;
        RECT  6.290000 37.020000  6.490000 37.220000 ;
        RECT  6.290000 37.460000  6.490000 37.660000 ;
        RECT  6.290000 37.900000  6.490000 38.100000 ;
        RECT  6.290000 49.715000  6.490000 49.915000 ;
        RECT  6.290000 50.135000  6.490000 50.335000 ;
        RECT  6.290000 50.555000  6.490000 50.755000 ;
        RECT  6.695000 34.820000  6.895000 35.020000 ;
        RECT  6.695000 35.260000  6.895000 35.460000 ;
        RECT  6.695000 35.700000  6.895000 35.900000 ;
        RECT  6.695000 36.140000  6.895000 36.340000 ;
        RECT  6.695000 36.580000  6.895000 36.780000 ;
        RECT  6.695000 37.020000  6.895000 37.220000 ;
        RECT  6.695000 37.460000  6.895000 37.660000 ;
        RECT  6.695000 37.900000  6.895000 38.100000 ;
        RECT  6.695000 49.715000  6.895000 49.915000 ;
        RECT  6.695000 50.135000  6.895000 50.335000 ;
        RECT  6.695000 50.555000  6.895000 50.755000 ;
        RECT  7.100000 34.820000  7.300000 35.020000 ;
        RECT  7.100000 35.260000  7.300000 35.460000 ;
        RECT  7.100000 35.700000  7.300000 35.900000 ;
        RECT  7.100000 36.140000  7.300000 36.340000 ;
        RECT  7.100000 36.580000  7.300000 36.780000 ;
        RECT  7.100000 37.020000  7.300000 37.220000 ;
        RECT  7.100000 37.460000  7.300000 37.660000 ;
        RECT  7.100000 37.900000  7.300000 38.100000 ;
        RECT  7.100000 49.715000  7.300000 49.915000 ;
        RECT  7.100000 50.135000  7.300000 50.335000 ;
        RECT  7.100000 50.555000  7.300000 50.755000 ;
        RECT  7.505000 34.820000  7.705000 35.020000 ;
        RECT  7.505000 35.260000  7.705000 35.460000 ;
        RECT  7.505000 35.700000  7.705000 35.900000 ;
        RECT  7.505000 36.140000  7.705000 36.340000 ;
        RECT  7.505000 36.580000  7.705000 36.780000 ;
        RECT  7.505000 37.020000  7.705000 37.220000 ;
        RECT  7.505000 37.460000  7.705000 37.660000 ;
        RECT  7.505000 37.900000  7.705000 38.100000 ;
        RECT  7.505000 49.715000  7.705000 49.915000 ;
        RECT  7.505000 50.135000  7.705000 50.335000 ;
        RECT  7.505000 50.555000  7.705000 50.755000 ;
        RECT  7.910000 34.820000  8.110000 35.020000 ;
        RECT  7.910000 35.260000  8.110000 35.460000 ;
        RECT  7.910000 35.700000  8.110000 35.900000 ;
        RECT  7.910000 36.140000  8.110000 36.340000 ;
        RECT  7.910000 36.580000  8.110000 36.780000 ;
        RECT  7.910000 37.020000  8.110000 37.220000 ;
        RECT  7.910000 37.460000  8.110000 37.660000 ;
        RECT  7.910000 37.900000  8.110000 38.100000 ;
        RECT  7.910000 49.715000  8.110000 49.915000 ;
        RECT  7.910000 50.135000  8.110000 50.335000 ;
        RECT  7.910000 50.555000  8.110000 50.755000 ;
        RECT  8.315000 34.820000  8.515000 35.020000 ;
        RECT  8.315000 35.260000  8.515000 35.460000 ;
        RECT  8.315000 35.700000  8.515000 35.900000 ;
        RECT  8.315000 36.140000  8.515000 36.340000 ;
        RECT  8.315000 36.580000  8.515000 36.780000 ;
        RECT  8.315000 37.020000  8.515000 37.220000 ;
        RECT  8.315000 37.460000  8.515000 37.660000 ;
        RECT  8.315000 37.900000  8.515000 38.100000 ;
        RECT  8.315000 49.715000  8.515000 49.915000 ;
        RECT  8.315000 50.135000  8.515000 50.335000 ;
        RECT  8.315000 50.555000  8.515000 50.755000 ;
        RECT  8.720000 34.820000  8.920000 35.020000 ;
        RECT  8.720000 35.260000  8.920000 35.460000 ;
        RECT  8.720000 35.700000  8.920000 35.900000 ;
        RECT  8.720000 36.140000  8.920000 36.340000 ;
        RECT  8.720000 36.580000  8.920000 36.780000 ;
        RECT  8.720000 37.020000  8.920000 37.220000 ;
        RECT  8.720000 37.460000  8.920000 37.660000 ;
        RECT  8.720000 37.900000  8.920000 38.100000 ;
        RECT  8.720000 49.715000  8.920000 49.915000 ;
        RECT  8.720000 50.135000  8.920000 50.335000 ;
        RECT  8.720000 50.555000  8.920000 50.755000 ;
        RECT  9.125000 34.820000  9.325000 35.020000 ;
        RECT  9.125000 35.260000  9.325000 35.460000 ;
        RECT  9.125000 35.700000  9.325000 35.900000 ;
        RECT  9.125000 36.140000  9.325000 36.340000 ;
        RECT  9.125000 36.580000  9.325000 36.780000 ;
        RECT  9.125000 37.020000  9.325000 37.220000 ;
        RECT  9.125000 37.460000  9.325000 37.660000 ;
        RECT  9.125000 37.900000  9.325000 38.100000 ;
        RECT  9.125000 49.715000  9.325000 49.915000 ;
        RECT  9.125000 50.135000  9.325000 50.335000 ;
        RECT  9.125000 50.555000  9.325000 50.755000 ;
        RECT  9.530000 34.820000  9.730000 35.020000 ;
        RECT  9.530000 35.260000  9.730000 35.460000 ;
        RECT  9.530000 35.700000  9.730000 35.900000 ;
        RECT  9.530000 36.140000  9.730000 36.340000 ;
        RECT  9.530000 36.580000  9.730000 36.780000 ;
        RECT  9.530000 37.020000  9.730000 37.220000 ;
        RECT  9.530000 37.460000  9.730000 37.660000 ;
        RECT  9.530000 37.900000  9.730000 38.100000 ;
        RECT  9.530000 49.715000  9.730000 49.915000 ;
        RECT  9.530000 50.135000  9.730000 50.335000 ;
        RECT  9.530000 50.555000  9.730000 50.755000 ;
        RECT  9.935000 34.820000 10.135000 35.020000 ;
        RECT  9.935000 35.260000 10.135000 35.460000 ;
        RECT  9.935000 35.700000 10.135000 35.900000 ;
        RECT  9.935000 36.140000 10.135000 36.340000 ;
        RECT  9.935000 36.580000 10.135000 36.780000 ;
        RECT  9.935000 37.020000 10.135000 37.220000 ;
        RECT  9.935000 37.460000 10.135000 37.660000 ;
        RECT  9.935000 37.900000 10.135000 38.100000 ;
        RECT  9.935000 49.715000 10.135000 49.915000 ;
        RECT  9.935000 50.135000 10.135000 50.335000 ;
        RECT  9.935000 50.555000 10.135000 50.755000 ;
        RECT 10.340000 34.820000 10.540000 35.020000 ;
        RECT 10.340000 35.260000 10.540000 35.460000 ;
        RECT 10.340000 35.700000 10.540000 35.900000 ;
        RECT 10.340000 36.140000 10.540000 36.340000 ;
        RECT 10.340000 36.580000 10.540000 36.780000 ;
        RECT 10.340000 37.020000 10.540000 37.220000 ;
        RECT 10.340000 37.460000 10.540000 37.660000 ;
        RECT 10.340000 37.900000 10.540000 38.100000 ;
        RECT 10.340000 49.715000 10.540000 49.915000 ;
        RECT 10.340000 50.135000 10.540000 50.335000 ;
        RECT 10.340000 50.555000 10.540000 50.755000 ;
        RECT 10.745000 34.820000 10.945000 35.020000 ;
        RECT 10.745000 35.260000 10.945000 35.460000 ;
        RECT 10.745000 35.700000 10.945000 35.900000 ;
        RECT 10.745000 36.140000 10.945000 36.340000 ;
        RECT 10.745000 36.580000 10.945000 36.780000 ;
        RECT 10.745000 37.020000 10.945000 37.220000 ;
        RECT 10.745000 37.460000 10.945000 37.660000 ;
        RECT 10.745000 37.900000 10.945000 38.100000 ;
        RECT 10.745000 49.715000 10.945000 49.915000 ;
        RECT 10.745000 50.135000 10.945000 50.335000 ;
        RECT 10.745000 50.555000 10.945000 50.755000 ;
        RECT 11.150000 34.820000 11.350000 35.020000 ;
        RECT 11.150000 35.260000 11.350000 35.460000 ;
        RECT 11.150000 35.700000 11.350000 35.900000 ;
        RECT 11.150000 36.140000 11.350000 36.340000 ;
        RECT 11.150000 36.580000 11.350000 36.780000 ;
        RECT 11.150000 37.020000 11.350000 37.220000 ;
        RECT 11.150000 37.460000 11.350000 37.660000 ;
        RECT 11.150000 37.900000 11.350000 38.100000 ;
        RECT 11.150000 49.715000 11.350000 49.915000 ;
        RECT 11.150000 50.135000 11.350000 50.335000 ;
        RECT 11.150000 50.555000 11.350000 50.755000 ;
        RECT 11.555000 34.820000 11.755000 35.020000 ;
        RECT 11.555000 35.260000 11.755000 35.460000 ;
        RECT 11.555000 35.700000 11.755000 35.900000 ;
        RECT 11.555000 36.140000 11.755000 36.340000 ;
        RECT 11.555000 36.580000 11.755000 36.780000 ;
        RECT 11.555000 37.020000 11.755000 37.220000 ;
        RECT 11.555000 37.460000 11.755000 37.660000 ;
        RECT 11.555000 37.900000 11.755000 38.100000 ;
        RECT 11.555000 49.715000 11.755000 49.915000 ;
        RECT 11.555000 50.135000 11.755000 50.335000 ;
        RECT 11.555000 50.555000 11.755000 50.755000 ;
        RECT 11.960000 34.820000 12.160000 35.020000 ;
        RECT 11.960000 35.260000 12.160000 35.460000 ;
        RECT 11.960000 35.700000 12.160000 35.900000 ;
        RECT 11.960000 36.140000 12.160000 36.340000 ;
        RECT 11.960000 36.580000 12.160000 36.780000 ;
        RECT 11.960000 37.020000 12.160000 37.220000 ;
        RECT 11.960000 37.460000 12.160000 37.660000 ;
        RECT 11.960000 37.900000 12.160000 38.100000 ;
        RECT 11.960000 49.715000 12.160000 49.915000 ;
        RECT 11.960000 50.135000 12.160000 50.335000 ;
        RECT 11.960000 50.555000 12.160000 50.755000 ;
        RECT 12.365000 34.820000 12.565000 35.020000 ;
        RECT 12.365000 35.260000 12.565000 35.460000 ;
        RECT 12.365000 35.700000 12.565000 35.900000 ;
        RECT 12.365000 36.140000 12.565000 36.340000 ;
        RECT 12.365000 36.580000 12.565000 36.780000 ;
        RECT 12.365000 37.020000 12.565000 37.220000 ;
        RECT 12.365000 37.460000 12.565000 37.660000 ;
        RECT 12.365000 37.900000 12.565000 38.100000 ;
        RECT 12.365000 49.715000 12.565000 49.915000 ;
        RECT 12.365000 50.135000 12.565000 50.335000 ;
        RECT 12.365000 50.555000 12.565000 50.755000 ;
        RECT 12.770000 34.820000 12.970000 35.020000 ;
        RECT 12.770000 35.260000 12.970000 35.460000 ;
        RECT 12.770000 35.700000 12.970000 35.900000 ;
        RECT 12.770000 36.140000 12.970000 36.340000 ;
        RECT 12.770000 36.580000 12.970000 36.780000 ;
        RECT 12.770000 37.020000 12.970000 37.220000 ;
        RECT 12.770000 37.460000 12.970000 37.660000 ;
        RECT 12.770000 37.900000 12.970000 38.100000 ;
        RECT 12.770000 49.715000 12.970000 49.915000 ;
        RECT 12.770000 50.135000 12.970000 50.335000 ;
        RECT 12.770000 50.555000 12.970000 50.755000 ;
        RECT 13.175000 34.820000 13.375000 35.020000 ;
        RECT 13.175000 35.260000 13.375000 35.460000 ;
        RECT 13.175000 35.700000 13.375000 35.900000 ;
        RECT 13.175000 36.140000 13.375000 36.340000 ;
        RECT 13.175000 36.580000 13.375000 36.780000 ;
        RECT 13.175000 37.020000 13.375000 37.220000 ;
        RECT 13.175000 37.460000 13.375000 37.660000 ;
        RECT 13.175000 37.900000 13.375000 38.100000 ;
        RECT 13.175000 49.715000 13.375000 49.915000 ;
        RECT 13.175000 50.135000 13.375000 50.335000 ;
        RECT 13.175000 50.555000 13.375000 50.755000 ;
        RECT 13.580000 34.820000 13.780000 35.020000 ;
        RECT 13.580000 35.260000 13.780000 35.460000 ;
        RECT 13.580000 35.700000 13.780000 35.900000 ;
        RECT 13.580000 36.140000 13.780000 36.340000 ;
        RECT 13.580000 36.580000 13.780000 36.780000 ;
        RECT 13.580000 37.020000 13.780000 37.220000 ;
        RECT 13.580000 37.460000 13.780000 37.660000 ;
        RECT 13.580000 37.900000 13.780000 38.100000 ;
        RECT 13.580000 49.715000 13.780000 49.915000 ;
        RECT 13.580000 50.135000 13.780000 50.335000 ;
        RECT 13.580000 50.555000 13.780000 50.755000 ;
        RECT 13.985000 34.820000 14.185000 35.020000 ;
        RECT 13.985000 35.260000 14.185000 35.460000 ;
        RECT 13.985000 35.700000 14.185000 35.900000 ;
        RECT 13.985000 36.140000 14.185000 36.340000 ;
        RECT 13.985000 36.580000 14.185000 36.780000 ;
        RECT 13.985000 37.020000 14.185000 37.220000 ;
        RECT 13.985000 37.460000 14.185000 37.660000 ;
        RECT 13.985000 37.900000 14.185000 38.100000 ;
        RECT 13.985000 49.715000 14.185000 49.915000 ;
        RECT 13.985000 50.135000 14.185000 50.335000 ;
        RECT 13.985000 50.555000 14.185000 50.755000 ;
        RECT 14.390000 34.820000 14.590000 35.020000 ;
        RECT 14.390000 35.260000 14.590000 35.460000 ;
        RECT 14.390000 35.700000 14.590000 35.900000 ;
        RECT 14.390000 36.140000 14.590000 36.340000 ;
        RECT 14.390000 36.580000 14.590000 36.780000 ;
        RECT 14.390000 37.020000 14.590000 37.220000 ;
        RECT 14.390000 37.460000 14.590000 37.660000 ;
        RECT 14.390000 37.900000 14.590000 38.100000 ;
        RECT 14.390000 49.715000 14.590000 49.915000 ;
        RECT 14.390000 50.135000 14.590000 50.335000 ;
        RECT 14.390000 50.555000 14.590000 50.755000 ;
        RECT 14.795000 34.820000 14.995000 35.020000 ;
        RECT 14.795000 35.260000 14.995000 35.460000 ;
        RECT 14.795000 35.700000 14.995000 35.900000 ;
        RECT 14.795000 36.140000 14.995000 36.340000 ;
        RECT 14.795000 36.580000 14.995000 36.780000 ;
        RECT 14.795000 37.020000 14.995000 37.220000 ;
        RECT 14.795000 37.460000 14.995000 37.660000 ;
        RECT 14.795000 37.900000 14.995000 38.100000 ;
        RECT 14.795000 49.715000 14.995000 49.915000 ;
        RECT 14.795000 50.135000 14.995000 50.335000 ;
        RECT 14.795000 50.555000 14.995000 50.755000 ;
        RECT 15.200000 34.820000 15.400000 35.020000 ;
        RECT 15.200000 35.260000 15.400000 35.460000 ;
        RECT 15.200000 35.700000 15.400000 35.900000 ;
        RECT 15.200000 36.140000 15.400000 36.340000 ;
        RECT 15.200000 36.580000 15.400000 36.780000 ;
        RECT 15.200000 37.020000 15.400000 37.220000 ;
        RECT 15.200000 37.460000 15.400000 37.660000 ;
        RECT 15.200000 37.900000 15.400000 38.100000 ;
        RECT 15.200000 49.715000 15.400000 49.915000 ;
        RECT 15.200000 50.135000 15.400000 50.335000 ;
        RECT 15.200000 50.555000 15.400000 50.755000 ;
        RECT 15.605000 34.820000 15.805000 35.020000 ;
        RECT 15.605000 35.260000 15.805000 35.460000 ;
        RECT 15.605000 35.700000 15.805000 35.900000 ;
        RECT 15.605000 36.140000 15.805000 36.340000 ;
        RECT 15.605000 36.580000 15.805000 36.780000 ;
        RECT 15.605000 37.020000 15.805000 37.220000 ;
        RECT 15.605000 37.460000 15.805000 37.660000 ;
        RECT 15.605000 37.900000 15.805000 38.100000 ;
        RECT 15.605000 49.715000 15.805000 49.915000 ;
        RECT 15.605000 50.135000 15.805000 50.335000 ;
        RECT 15.605000 50.555000 15.805000 50.755000 ;
        RECT 16.010000 34.820000 16.210000 35.020000 ;
        RECT 16.010000 35.260000 16.210000 35.460000 ;
        RECT 16.010000 35.700000 16.210000 35.900000 ;
        RECT 16.010000 36.140000 16.210000 36.340000 ;
        RECT 16.010000 36.580000 16.210000 36.780000 ;
        RECT 16.010000 37.020000 16.210000 37.220000 ;
        RECT 16.010000 37.460000 16.210000 37.660000 ;
        RECT 16.010000 37.900000 16.210000 38.100000 ;
        RECT 16.010000 49.715000 16.210000 49.915000 ;
        RECT 16.010000 50.135000 16.210000 50.335000 ;
        RECT 16.010000 50.555000 16.210000 50.755000 ;
        RECT 16.415000 34.820000 16.615000 35.020000 ;
        RECT 16.415000 35.260000 16.615000 35.460000 ;
        RECT 16.415000 35.700000 16.615000 35.900000 ;
        RECT 16.415000 36.140000 16.615000 36.340000 ;
        RECT 16.415000 36.580000 16.615000 36.780000 ;
        RECT 16.415000 37.020000 16.615000 37.220000 ;
        RECT 16.415000 37.460000 16.615000 37.660000 ;
        RECT 16.415000 37.900000 16.615000 38.100000 ;
        RECT 16.415000 49.715000 16.615000 49.915000 ;
        RECT 16.415000 50.135000 16.615000 50.335000 ;
        RECT 16.415000 50.555000 16.615000 50.755000 ;
        RECT 16.820000 34.820000 17.020000 35.020000 ;
        RECT 16.820000 35.260000 17.020000 35.460000 ;
        RECT 16.820000 35.700000 17.020000 35.900000 ;
        RECT 16.820000 36.140000 17.020000 36.340000 ;
        RECT 16.820000 36.580000 17.020000 36.780000 ;
        RECT 16.820000 37.020000 17.020000 37.220000 ;
        RECT 16.820000 37.460000 17.020000 37.660000 ;
        RECT 16.820000 37.900000 17.020000 38.100000 ;
        RECT 16.820000 49.715000 17.020000 49.915000 ;
        RECT 16.820000 50.135000 17.020000 50.335000 ;
        RECT 16.820000 50.555000 17.020000 50.755000 ;
        RECT 17.225000 34.820000 17.425000 35.020000 ;
        RECT 17.225000 35.260000 17.425000 35.460000 ;
        RECT 17.225000 35.700000 17.425000 35.900000 ;
        RECT 17.225000 36.140000 17.425000 36.340000 ;
        RECT 17.225000 36.580000 17.425000 36.780000 ;
        RECT 17.225000 37.020000 17.425000 37.220000 ;
        RECT 17.225000 37.460000 17.425000 37.660000 ;
        RECT 17.225000 37.900000 17.425000 38.100000 ;
        RECT 17.225000 49.715000 17.425000 49.915000 ;
        RECT 17.225000 50.135000 17.425000 50.335000 ;
        RECT 17.225000 50.555000 17.425000 50.755000 ;
        RECT 17.630000 34.820000 17.830000 35.020000 ;
        RECT 17.630000 35.260000 17.830000 35.460000 ;
        RECT 17.630000 35.700000 17.830000 35.900000 ;
        RECT 17.630000 36.140000 17.830000 36.340000 ;
        RECT 17.630000 36.580000 17.830000 36.780000 ;
        RECT 17.630000 37.020000 17.830000 37.220000 ;
        RECT 17.630000 37.460000 17.830000 37.660000 ;
        RECT 17.630000 37.900000 17.830000 38.100000 ;
        RECT 17.630000 49.715000 17.830000 49.915000 ;
        RECT 17.630000 50.135000 17.830000 50.335000 ;
        RECT 17.630000 50.555000 17.830000 50.755000 ;
        RECT 18.035000 34.820000 18.235000 35.020000 ;
        RECT 18.035000 35.260000 18.235000 35.460000 ;
        RECT 18.035000 35.700000 18.235000 35.900000 ;
        RECT 18.035000 36.140000 18.235000 36.340000 ;
        RECT 18.035000 36.580000 18.235000 36.780000 ;
        RECT 18.035000 37.020000 18.235000 37.220000 ;
        RECT 18.035000 37.460000 18.235000 37.660000 ;
        RECT 18.035000 37.900000 18.235000 38.100000 ;
        RECT 18.035000 49.715000 18.235000 49.915000 ;
        RECT 18.035000 50.135000 18.235000 50.335000 ;
        RECT 18.035000 50.555000 18.235000 50.755000 ;
        RECT 18.440000 34.820000 18.640000 35.020000 ;
        RECT 18.440000 35.260000 18.640000 35.460000 ;
        RECT 18.440000 35.700000 18.640000 35.900000 ;
        RECT 18.440000 36.140000 18.640000 36.340000 ;
        RECT 18.440000 36.580000 18.640000 36.780000 ;
        RECT 18.440000 37.020000 18.640000 37.220000 ;
        RECT 18.440000 37.460000 18.640000 37.660000 ;
        RECT 18.440000 37.900000 18.640000 38.100000 ;
        RECT 18.440000 49.715000 18.640000 49.915000 ;
        RECT 18.440000 50.135000 18.640000 50.335000 ;
        RECT 18.440000 50.555000 18.640000 50.755000 ;
        RECT 18.845000 34.820000 19.045000 35.020000 ;
        RECT 18.845000 35.260000 19.045000 35.460000 ;
        RECT 18.845000 35.700000 19.045000 35.900000 ;
        RECT 18.845000 36.140000 19.045000 36.340000 ;
        RECT 18.845000 36.580000 19.045000 36.780000 ;
        RECT 18.845000 37.020000 19.045000 37.220000 ;
        RECT 18.845000 37.460000 19.045000 37.660000 ;
        RECT 18.845000 37.900000 19.045000 38.100000 ;
        RECT 18.845000 49.715000 19.045000 49.915000 ;
        RECT 18.845000 50.135000 19.045000 50.335000 ;
        RECT 18.845000 50.555000 19.045000 50.755000 ;
        RECT 19.250000 34.820000 19.450000 35.020000 ;
        RECT 19.250000 35.260000 19.450000 35.460000 ;
        RECT 19.250000 35.700000 19.450000 35.900000 ;
        RECT 19.250000 36.140000 19.450000 36.340000 ;
        RECT 19.250000 36.580000 19.450000 36.780000 ;
        RECT 19.250000 37.020000 19.450000 37.220000 ;
        RECT 19.250000 37.460000 19.450000 37.660000 ;
        RECT 19.250000 37.900000 19.450000 38.100000 ;
        RECT 19.250000 49.715000 19.450000 49.915000 ;
        RECT 19.250000 50.135000 19.450000 50.335000 ;
        RECT 19.250000 50.555000 19.450000 50.755000 ;
        RECT 19.655000 34.820000 19.855000 35.020000 ;
        RECT 19.655000 35.260000 19.855000 35.460000 ;
        RECT 19.655000 35.700000 19.855000 35.900000 ;
        RECT 19.655000 36.140000 19.855000 36.340000 ;
        RECT 19.655000 36.580000 19.855000 36.780000 ;
        RECT 19.655000 37.020000 19.855000 37.220000 ;
        RECT 19.655000 37.460000 19.855000 37.660000 ;
        RECT 19.655000 37.900000 19.855000 38.100000 ;
        RECT 19.655000 49.715000 19.855000 49.915000 ;
        RECT 19.655000 50.135000 19.855000 50.335000 ;
        RECT 19.655000 50.555000 19.855000 50.755000 ;
        RECT 20.060000 34.820000 20.260000 35.020000 ;
        RECT 20.060000 35.260000 20.260000 35.460000 ;
        RECT 20.060000 35.700000 20.260000 35.900000 ;
        RECT 20.060000 36.140000 20.260000 36.340000 ;
        RECT 20.060000 36.580000 20.260000 36.780000 ;
        RECT 20.060000 37.020000 20.260000 37.220000 ;
        RECT 20.060000 37.460000 20.260000 37.660000 ;
        RECT 20.060000 37.900000 20.260000 38.100000 ;
        RECT 20.060000 49.715000 20.260000 49.915000 ;
        RECT 20.060000 50.135000 20.260000 50.335000 ;
        RECT 20.060000 50.555000 20.260000 50.755000 ;
        RECT 20.465000 34.820000 20.665000 35.020000 ;
        RECT 20.465000 35.260000 20.665000 35.460000 ;
        RECT 20.465000 35.700000 20.665000 35.900000 ;
        RECT 20.465000 36.140000 20.665000 36.340000 ;
        RECT 20.465000 36.580000 20.665000 36.780000 ;
        RECT 20.465000 37.020000 20.665000 37.220000 ;
        RECT 20.465000 37.460000 20.665000 37.660000 ;
        RECT 20.465000 37.900000 20.665000 38.100000 ;
        RECT 20.465000 49.715000 20.665000 49.915000 ;
        RECT 20.465000 50.135000 20.665000 50.335000 ;
        RECT 20.465000 50.555000 20.665000 50.755000 ;
        RECT 20.870000 34.820000 21.070000 35.020000 ;
        RECT 20.870000 35.260000 21.070000 35.460000 ;
        RECT 20.870000 35.700000 21.070000 35.900000 ;
        RECT 20.870000 36.140000 21.070000 36.340000 ;
        RECT 20.870000 36.580000 21.070000 36.780000 ;
        RECT 20.870000 37.020000 21.070000 37.220000 ;
        RECT 20.870000 37.460000 21.070000 37.660000 ;
        RECT 20.870000 37.900000 21.070000 38.100000 ;
        RECT 20.870000 49.715000 21.070000 49.915000 ;
        RECT 20.870000 50.135000 21.070000 50.335000 ;
        RECT 20.870000 50.555000 21.070000 50.755000 ;
        RECT 21.275000 34.820000 21.475000 35.020000 ;
        RECT 21.275000 35.260000 21.475000 35.460000 ;
        RECT 21.275000 35.700000 21.475000 35.900000 ;
        RECT 21.275000 36.140000 21.475000 36.340000 ;
        RECT 21.275000 36.580000 21.475000 36.780000 ;
        RECT 21.275000 37.020000 21.475000 37.220000 ;
        RECT 21.275000 37.460000 21.475000 37.660000 ;
        RECT 21.275000 37.900000 21.475000 38.100000 ;
        RECT 21.275000 49.715000 21.475000 49.915000 ;
        RECT 21.275000 50.135000 21.475000 50.335000 ;
        RECT 21.275000 50.555000 21.475000 50.755000 ;
        RECT 21.680000 34.820000 21.880000 35.020000 ;
        RECT 21.680000 35.260000 21.880000 35.460000 ;
        RECT 21.680000 35.700000 21.880000 35.900000 ;
        RECT 21.680000 36.140000 21.880000 36.340000 ;
        RECT 21.680000 36.580000 21.880000 36.780000 ;
        RECT 21.680000 37.020000 21.880000 37.220000 ;
        RECT 21.680000 37.460000 21.880000 37.660000 ;
        RECT 21.680000 37.900000 21.880000 38.100000 ;
        RECT 21.680000 49.715000 21.880000 49.915000 ;
        RECT 21.680000 50.135000 21.880000 50.335000 ;
        RECT 21.680000 50.555000 21.880000 50.755000 ;
        RECT 22.085000 34.820000 22.285000 35.020000 ;
        RECT 22.085000 35.260000 22.285000 35.460000 ;
        RECT 22.085000 35.700000 22.285000 35.900000 ;
        RECT 22.085000 36.140000 22.285000 36.340000 ;
        RECT 22.085000 36.580000 22.285000 36.780000 ;
        RECT 22.085000 37.020000 22.285000 37.220000 ;
        RECT 22.085000 37.460000 22.285000 37.660000 ;
        RECT 22.085000 37.900000 22.285000 38.100000 ;
        RECT 22.085000 49.715000 22.285000 49.915000 ;
        RECT 22.085000 50.135000 22.285000 50.335000 ;
        RECT 22.085000 50.555000 22.285000 50.755000 ;
        RECT 22.490000 34.820000 22.690000 35.020000 ;
        RECT 22.490000 35.260000 22.690000 35.460000 ;
        RECT 22.490000 35.700000 22.690000 35.900000 ;
        RECT 22.490000 36.140000 22.690000 36.340000 ;
        RECT 22.490000 36.580000 22.690000 36.780000 ;
        RECT 22.490000 37.020000 22.690000 37.220000 ;
        RECT 22.490000 37.460000 22.690000 37.660000 ;
        RECT 22.490000 37.900000 22.690000 38.100000 ;
        RECT 22.490000 49.715000 22.690000 49.915000 ;
        RECT 22.490000 50.135000 22.690000 50.335000 ;
        RECT 22.490000 50.555000 22.690000 50.755000 ;
        RECT 22.895000 34.820000 23.095000 35.020000 ;
        RECT 22.895000 35.260000 23.095000 35.460000 ;
        RECT 22.895000 35.700000 23.095000 35.900000 ;
        RECT 22.895000 36.140000 23.095000 36.340000 ;
        RECT 22.895000 36.580000 23.095000 36.780000 ;
        RECT 22.895000 37.020000 23.095000 37.220000 ;
        RECT 22.895000 37.460000 23.095000 37.660000 ;
        RECT 22.895000 37.900000 23.095000 38.100000 ;
        RECT 22.895000 49.715000 23.095000 49.915000 ;
        RECT 22.895000 50.135000 23.095000 50.335000 ;
        RECT 22.895000 50.555000 23.095000 50.755000 ;
        RECT 23.300000 34.820000 23.500000 35.020000 ;
        RECT 23.300000 35.260000 23.500000 35.460000 ;
        RECT 23.300000 35.700000 23.500000 35.900000 ;
        RECT 23.300000 36.140000 23.500000 36.340000 ;
        RECT 23.300000 36.580000 23.500000 36.780000 ;
        RECT 23.300000 37.020000 23.500000 37.220000 ;
        RECT 23.300000 37.460000 23.500000 37.660000 ;
        RECT 23.300000 37.900000 23.500000 38.100000 ;
        RECT 23.300000 49.715000 23.500000 49.915000 ;
        RECT 23.300000 50.135000 23.500000 50.335000 ;
        RECT 23.300000 50.555000 23.500000 50.755000 ;
        RECT 23.705000 34.820000 23.905000 35.020000 ;
        RECT 23.705000 35.260000 23.905000 35.460000 ;
        RECT 23.705000 35.700000 23.905000 35.900000 ;
        RECT 23.705000 36.140000 23.905000 36.340000 ;
        RECT 23.705000 36.580000 23.905000 36.780000 ;
        RECT 23.705000 37.020000 23.905000 37.220000 ;
        RECT 23.705000 37.460000 23.905000 37.660000 ;
        RECT 23.705000 37.900000 23.905000 38.100000 ;
        RECT 23.705000 49.715000 23.905000 49.915000 ;
        RECT 23.705000 50.135000 23.905000 50.335000 ;
        RECT 23.705000 50.555000 23.905000 50.755000 ;
        RECT 24.110000 34.820000 24.310000 35.020000 ;
        RECT 24.110000 35.260000 24.310000 35.460000 ;
        RECT 24.110000 35.700000 24.310000 35.900000 ;
        RECT 24.110000 36.140000 24.310000 36.340000 ;
        RECT 24.110000 36.580000 24.310000 36.780000 ;
        RECT 24.110000 37.020000 24.310000 37.220000 ;
        RECT 24.110000 37.460000 24.310000 37.660000 ;
        RECT 24.110000 37.900000 24.310000 38.100000 ;
        RECT 24.110000 49.715000 24.310000 49.915000 ;
        RECT 24.110000 50.135000 24.310000 50.335000 ;
        RECT 24.110000 50.555000 24.310000 50.755000 ;
        RECT 50.845000 34.820000 51.045000 35.020000 ;
        RECT 50.845000 35.260000 51.045000 35.460000 ;
        RECT 50.845000 35.700000 51.045000 35.900000 ;
        RECT 50.845000 36.140000 51.045000 36.340000 ;
        RECT 50.845000 36.580000 51.045000 36.780000 ;
        RECT 50.845000 37.020000 51.045000 37.220000 ;
        RECT 50.845000 37.460000 51.045000 37.660000 ;
        RECT 50.845000 37.900000 51.045000 38.100000 ;
        RECT 50.845000 49.715000 51.045000 49.915000 ;
        RECT 50.845000 50.135000 51.045000 50.335000 ;
        RECT 50.845000 50.555000 51.045000 50.755000 ;
        RECT 51.255000 34.820000 51.455000 35.020000 ;
        RECT 51.255000 35.260000 51.455000 35.460000 ;
        RECT 51.255000 35.700000 51.455000 35.900000 ;
        RECT 51.255000 36.140000 51.455000 36.340000 ;
        RECT 51.255000 36.580000 51.455000 36.780000 ;
        RECT 51.255000 37.020000 51.455000 37.220000 ;
        RECT 51.255000 37.460000 51.455000 37.660000 ;
        RECT 51.255000 37.900000 51.455000 38.100000 ;
        RECT 51.255000 49.715000 51.455000 49.915000 ;
        RECT 51.255000 50.135000 51.455000 50.335000 ;
        RECT 51.255000 50.555000 51.455000 50.755000 ;
        RECT 51.665000 34.820000 51.865000 35.020000 ;
        RECT 51.665000 35.260000 51.865000 35.460000 ;
        RECT 51.665000 35.700000 51.865000 35.900000 ;
        RECT 51.665000 36.140000 51.865000 36.340000 ;
        RECT 51.665000 36.580000 51.865000 36.780000 ;
        RECT 51.665000 37.020000 51.865000 37.220000 ;
        RECT 51.665000 37.460000 51.865000 37.660000 ;
        RECT 51.665000 37.900000 51.865000 38.100000 ;
        RECT 51.665000 49.715000 51.865000 49.915000 ;
        RECT 51.665000 50.135000 51.865000 50.335000 ;
        RECT 51.665000 50.555000 51.865000 50.755000 ;
        RECT 52.075000 34.820000 52.275000 35.020000 ;
        RECT 52.075000 35.260000 52.275000 35.460000 ;
        RECT 52.075000 35.700000 52.275000 35.900000 ;
        RECT 52.075000 36.140000 52.275000 36.340000 ;
        RECT 52.075000 36.580000 52.275000 36.780000 ;
        RECT 52.075000 37.020000 52.275000 37.220000 ;
        RECT 52.075000 37.460000 52.275000 37.660000 ;
        RECT 52.075000 37.900000 52.275000 38.100000 ;
        RECT 52.075000 49.715000 52.275000 49.915000 ;
        RECT 52.075000 50.135000 52.275000 50.335000 ;
        RECT 52.075000 50.555000 52.275000 50.755000 ;
        RECT 52.485000 34.820000 52.685000 35.020000 ;
        RECT 52.485000 35.260000 52.685000 35.460000 ;
        RECT 52.485000 35.700000 52.685000 35.900000 ;
        RECT 52.485000 36.140000 52.685000 36.340000 ;
        RECT 52.485000 36.580000 52.685000 36.780000 ;
        RECT 52.485000 37.020000 52.685000 37.220000 ;
        RECT 52.485000 37.460000 52.685000 37.660000 ;
        RECT 52.485000 37.900000 52.685000 38.100000 ;
        RECT 52.485000 49.715000 52.685000 49.915000 ;
        RECT 52.485000 50.135000 52.685000 50.335000 ;
        RECT 52.485000 50.555000 52.685000 50.755000 ;
        RECT 52.895000 34.820000 53.095000 35.020000 ;
        RECT 52.895000 35.260000 53.095000 35.460000 ;
        RECT 52.895000 35.700000 53.095000 35.900000 ;
        RECT 52.895000 36.140000 53.095000 36.340000 ;
        RECT 52.895000 36.580000 53.095000 36.780000 ;
        RECT 52.895000 37.020000 53.095000 37.220000 ;
        RECT 52.895000 37.460000 53.095000 37.660000 ;
        RECT 52.895000 37.900000 53.095000 38.100000 ;
        RECT 52.895000 49.715000 53.095000 49.915000 ;
        RECT 52.895000 50.135000 53.095000 50.335000 ;
        RECT 52.895000 50.555000 53.095000 50.755000 ;
        RECT 53.305000 34.820000 53.505000 35.020000 ;
        RECT 53.305000 35.260000 53.505000 35.460000 ;
        RECT 53.305000 35.700000 53.505000 35.900000 ;
        RECT 53.305000 36.140000 53.505000 36.340000 ;
        RECT 53.305000 36.580000 53.505000 36.780000 ;
        RECT 53.305000 37.020000 53.505000 37.220000 ;
        RECT 53.305000 37.460000 53.505000 37.660000 ;
        RECT 53.305000 37.900000 53.505000 38.100000 ;
        RECT 53.305000 49.715000 53.505000 49.915000 ;
        RECT 53.305000 50.135000 53.505000 50.335000 ;
        RECT 53.305000 50.555000 53.505000 50.755000 ;
        RECT 53.710000 34.820000 53.910000 35.020000 ;
        RECT 53.710000 35.260000 53.910000 35.460000 ;
        RECT 53.710000 35.700000 53.910000 35.900000 ;
        RECT 53.710000 36.140000 53.910000 36.340000 ;
        RECT 53.710000 36.580000 53.910000 36.780000 ;
        RECT 53.710000 37.020000 53.910000 37.220000 ;
        RECT 53.710000 37.460000 53.910000 37.660000 ;
        RECT 53.710000 37.900000 53.910000 38.100000 ;
        RECT 53.710000 49.715000 53.910000 49.915000 ;
        RECT 53.710000 50.135000 53.910000 50.335000 ;
        RECT 53.710000 50.555000 53.910000 50.755000 ;
        RECT 54.115000 34.820000 54.315000 35.020000 ;
        RECT 54.115000 35.260000 54.315000 35.460000 ;
        RECT 54.115000 35.700000 54.315000 35.900000 ;
        RECT 54.115000 36.140000 54.315000 36.340000 ;
        RECT 54.115000 36.580000 54.315000 36.780000 ;
        RECT 54.115000 37.020000 54.315000 37.220000 ;
        RECT 54.115000 37.460000 54.315000 37.660000 ;
        RECT 54.115000 37.900000 54.315000 38.100000 ;
        RECT 54.115000 49.715000 54.315000 49.915000 ;
        RECT 54.115000 50.135000 54.315000 50.335000 ;
        RECT 54.115000 50.555000 54.315000 50.755000 ;
        RECT 54.520000 34.820000 54.720000 35.020000 ;
        RECT 54.520000 35.260000 54.720000 35.460000 ;
        RECT 54.520000 35.700000 54.720000 35.900000 ;
        RECT 54.520000 36.140000 54.720000 36.340000 ;
        RECT 54.520000 36.580000 54.720000 36.780000 ;
        RECT 54.520000 37.020000 54.720000 37.220000 ;
        RECT 54.520000 37.460000 54.720000 37.660000 ;
        RECT 54.520000 37.900000 54.720000 38.100000 ;
        RECT 54.520000 49.715000 54.720000 49.915000 ;
        RECT 54.520000 50.135000 54.720000 50.335000 ;
        RECT 54.520000 50.555000 54.720000 50.755000 ;
        RECT 54.925000 34.820000 55.125000 35.020000 ;
        RECT 54.925000 35.260000 55.125000 35.460000 ;
        RECT 54.925000 35.700000 55.125000 35.900000 ;
        RECT 54.925000 36.140000 55.125000 36.340000 ;
        RECT 54.925000 36.580000 55.125000 36.780000 ;
        RECT 54.925000 37.020000 55.125000 37.220000 ;
        RECT 54.925000 37.460000 55.125000 37.660000 ;
        RECT 54.925000 37.900000 55.125000 38.100000 ;
        RECT 54.925000 49.715000 55.125000 49.915000 ;
        RECT 54.925000 50.135000 55.125000 50.335000 ;
        RECT 54.925000 50.555000 55.125000 50.755000 ;
        RECT 55.330000 34.820000 55.530000 35.020000 ;
        RECT 55.330000 35.260000 55.530000 35.460000 ;
        RECT 55.330000 35.700000 55.530000 35.900000 ;
        RECT 55.330000 36.140000 55.530000 36.340000 ;
        RECT 55.330000 36.580000 55.530000 36.780000 ;
        RECT 55.330000 37.020000 55.530000 37.220000 ;
        RECT 55.330000 37.460000 55.530000 37.660000 ;
        RECT 55.330000 37.900000 55.530000 38.100000 ;
        RECT 55.330000 49.715000 55.530000 49.915000 ;
        RECT 55.330000 50.135000 55.530000 50.335000 ;
        RECT 55.330000 50.555000 55.530000 50.755000 ;
        RECT 55.735000 34.820000 55.935000 35.020000 ;
        RECT 55.735000 35.260000 55.935000 35.460000 ;
        RECT 55.735000 35.700000 55.935000 35.900000 ;
        RECT 55.735000 36.140000 55.935000 36.340000 ;
        RECT 55.735000 36.580000 55.935000 36.780000 ;
        RECT 55.735000 37.020000 55.935000 37.220000 ;
        RECT 55.735000 37.460000 55.935000 37.660000 ;
        RECT 55.735000 37.900000 55.935000 38.100000 ;
        RECT 55.735000 49.715000 55.935000 49.915000 ;
        RECT 55.735000 50.135000 55.935000 50.335000 ;
        RECT 55.735000 50.555000 55.935000 50.755000 ;
        RECT 56.140000 34.820000 56.340000 35.020000 ;
        RECT 56.140000 35.260000 56.340000 35.460000 ;
        RECT 56.140000 35.700000 56.340000 35.900000 ;
        RECT 56.140000 36.140000 56.340000 36.340000 ;
        RECT 56.140000 36.580000 56.340000 36.780000 ;
        RECT 56.140000 37.020000 56.340000 37.220000 ;
        RECT 56.140000 37.460000 56.340000 37.660000 ;
        RECT 56.140000 37.900000 56.340000 38.100000 ;
        RECT 56.140000 49.715000 56.340000 49.915000 ;
        RECT 56.140000 50.135000 56.340000 50.335000 ;
        RECT 56.140000 50.555000 56.340000 50.755000 ;
        RECT 56.545000 34.820000 56.745000 35.020000 ;
        RECT 56.545000 35.260000 56.745000 35.460000 ;
        RECT 56.545000 35.700000 56.745000 35.900000 ;
        RECT 56.545000 36.140000 56.745000 36.340000 ;
        RECT 56.545000 36.580000 56.745000 36.780000 ;
        RECT 56.545000 37.020000 56.745000 37.220000 ;
        RECT 56.545000 37.460000 56.745000 37.660000 ;
        RECT 56.545000 37.900000 56.745000 38.100000 ;
        RECT 56.545000 49.715000 56.745000 49.915000 ;
        RECT 56.545000 50.135000 56.745000 50.335000 ;
        RECT 56.545000 50.555000 56.745000 50.755000 ;
        RECT 56.950000 34.820000 57.150000 35.020000 ;
        RECT 56.950000 35.260000 57.150000 35.460000 ;
        RECT 56.950000 35.700000 57.150000 35.900000 ;
        RECT 56.950000 36.140000 57.150000 36.340000 ;
        RECT 56.950000 36.580000 57.150000 36.780000 ;
        RECT 56.950000 37.020000 57.150000 37.220000 ;
        RECT 56.950000 37.460000 57.150000 37.660000 ;
        RECT 56.950000 37.900000 57.150000 38.100000 ;
        RECT 56.950000 49.715000 57.150000 49.915000 ;
        RECT 56.950000 50.135000 57.150000 50.335000 ;
        RECT 56.950000 50.555000 57.150000 50.755000 ;
        RECT 57.355000 34.820000 57.555000 35.020000 ;
        RECT 57.355000 35.260000 57.555000 35.460000 ;
        RECT 57.355000 35.700000 57.555000 35.900000 ;
        RECT 57.355000 36.140000 57.555000 36.340000 ;
        RECT 57.355000 36.580000 57.555000 36.780000 ;
        RECT 57.355000 37.020000 57.555000 37.220000 ;
        RECT 57.355000 37.460000 57.555000 37.660000 ;
        RECT 57.355000 37.900000 57.555000 38.100000 ;
        RECT 57.355000 49.715000 57.555000 49.915000 ;
        RECT 57.355000 50.135000 57.555000 50.335000 ;
        RECT 57.355000 50.555000 57.555000 50.755000 ;
        RECT 57.760000 34.820000 57.960000 35.020000 ;
        RECT 57.760000 35.260000 57.960000 35.460000 ;
        RECT 57.760000 35.700000 57.960000 35.900000 ;
        RECT 57.760000 36.140000 57.960000 36.340000 ;
        RECT 57.760000 36.580000 57.960000 36.780000 ;
        RECT 57.760000 37.020000 57.960000 37.220000 ;
        RECT 57.760000 37.460000 57.960000 37.660000 ;
        RECT 57.760000 37.900000 57.960000 38.100000 ;
        RECT 57.760000 49.715000 57.960000 49.915000 ;
        RECT 57.760000 50.135000 57.960000 50.335000 ;
        RECT 57.760000 50.555000 57.960000 50.755000 ;
        RECT 58.165000 34.820000 58.365000 35.020000 ;
        RECT 58.165000 35.260000 58.365000 35.460000 ;
        RECT 58.165000 35.700000 58.365000 35.900000 ;
        RECT 58.165000 36.140000 58.365000 36.340000 ;
        RECT 58.165000 36.580000 58.365000 36.780000 ;
        RECT 58.165000 37.020000 58.365000 37.220000 ;
        RECT 58.165000 37.460000 58.365000 37.660000 ;
        RECT 58.165000 37.900000 58.365000 38.100000 ;
        RECT 58.165000 49.715000 58.365000 49.915000 ;
        RECT 58.165000 50.135000 58.365000 50.335000 ;
        RECT 58.165000 50.555000 58.365000 50.755000 ;
        RECT 58.570000 34.820000 58.770000 35.020000 ;
        RECT 58.570000 35.260000 58.770000 35.460000 ;
        RECT 58.570000 35.700000 58.770000 35.900000 ;
        RECT 58.570000 36.140000 58.770000 36.340000 ;
        RECT 58.570000 36.580000 58.770000 36.780000 ;
        RECT 58.570000 37.020000 58.770000 37.220000 ;
        RECT 58.570000 37.460000 58.770000 37.660000 ;
        RECT 58.570000 37.900000 58.770000 38.100000 ;
        RECT 58.570000 49.715000 58.770000 49.915000 ;
        RECT 58.570000 50.135000 58.770000 50.335000 ;
        RECT 58.570000 50.555000 58.770000 50.755000 ;
        RECT 58.975000 34.820000 59.175000 35.020000 ;
        RECT 58.975000 35.260000 59.175000 35.460000 ;
        RECT 58.975000 35.700000 59.175000 35.900000 ;
        RECT 58.975000 36.140000 59.175000 36.340000 ;
        RECT 58.975000 36.580000 59.175000 36.780000 ;
        RECT 58.975000 37.020000 59.175000 37.220000 ;
        RECT 58.975000 37.460000 59.175000 37.660000 ;
        RECT 58.975000 37.900000 59.175000 38.100000 ;
        RECT 58.975000 49.715000 59.175000 49.915000 ;
        RECT 58.975000 50.135000 59.175000 50.335000 ;
        RECT 58.975000 50.555000 59.175000 50.755000 ;
        RECT 59.380000 34.820000 59.580000 35.020000 ;
        RECT 59.380000 35.260000 59.580000 35.460000 ;
        RECT 59.380000 35.700000 59.580000 35.900000 ;
        RECT 59.380000 36.140000 59.580000 36.340000 ;
        RECT 59.380000 36.580000 59.580000 36.780000 ;
        RECT 59.380000 37.020000 59.580000 37.220000 ;
        RECT 59.380000 37.460000 59.580000 37.660000 ;
        RECT 59.380000 37.900000 59.580000 38.100000 ;
        RECT 59.380000 49.715000 59.580000 49.915000 ;
        RECT 59.380000 50.135000 59.580000 50.335000 ;
        RECT 59.380000 50.555000 59.580000 50.755000 ;
        RECT 59.785000 34.820000 59.985000 35.020000 ;
        RECT 59.785000 35.260000 59.985000 35.460000 ;
        RECT 59.785000 35.700000 59.985000 35.900000 ;
        RECT 59.785000 36.140000 59.985000 36.340000 ;
        RECT 59.785000 36.580000 59.985000 36.780000 ;
        RECT 59.785000 37.020000 59.985000 37.220000 ;
        RECT 59.785000 37.460000 59.985000 37.660000 ;
        RECT 59.785000 37.900000 59.985000 38.100000 ;
        RECT 59.785000 49.715000 59.985000 49.915000 ;
        RECT 59.785000 50.135000 59.985000 50.335000 ;
        RECT 59.785000 50.555000 59.985000 50.755000 ;
        RECT 60.190000 34.820000 60.390000 35.020000 ;
        RECT 60.190000 35.260000 60.390000 35.460000 ;
        RECT 60.190000 35.700000 60.390000 35.900000 ;
        RECT 60.190000 36.140000 60.390000 36.340000 ;
        RECT 60.190000 36.580000 60.390000 36.780000 ;
        RECT 60.190000 37.020000 60.390000 37.220000 ;
        RECT 60.190000 37.460000 60.390000 37.660000 ;
        RECT 60.190000 37.900000 60.390000 38.100000 ;
        RECT 60.190000 49.715000 60.390000 49.915000 ;
        RECT 60.190000 50.135000 60.390000 50.335000 ;
        RECT 60.190000 50.555000 60.390000 50.755000 ;
        RECT 60.595000 34.820000 60.795000 35.020000 ;
        RECT 60.595000 35.260000 60.795000 35.460000 ;
        RECT 60.595000 35.700000 60.795000 35.900000 ;
        RECT 60.595000 36.140000 60.795000 36.340000 ;
        RECT 60.595000 36.580000 60.795000 36.780000 ;
        RECT 60.595000 37.020000 60.795000 37.220000 ;
        RECT 60.595000 37.460000 60.795000 37.660000 ;
        RECT 60.595000 37.900000 60.795000 38.100000 ;
        RECT 60.595000 49.715000 60.795000 49.915000 ;
        RECT 60.595000 50.135000 60.795000 50.335000 ;
        RECT 60.595000 50.555000 60.795000 50.755000 ;
        RECT 61.000000 34.820000 61.200000 35.020000 ;
        RECT 61.000000 35.260000 61.200000 35.460000 ;
        RECT 61.000000 35.700000 61.200000 35.900000 ;
        RECT 61.000000 36.140000 61.200000 36.340000 ;
        RECT 61.000000 36.580000 61.200000 36.780000 ;
        RECT 61.000000 37.020000 61.200000 37.220000 ;
        RECT 61.000000 37.460000 61.200000 37.660000 ;
        RECT 61.000000 37.900000 61.200000 38.100000 ;
        RECT 61.000000 49.715000 61.200000 49.915000 ;
        RECT 61.000000 50.135000 61.200000 50.335000 ;
        RECT 61.000000 50.555000 61.200000 50.755000 ;
        RECT 61.405000 34.820000 61.605000 35.020000 ;
        RECT 61.405000 35.260000 61.605000 35.460000 ;
        RECT 61.405000 35.700000 61.605000 35.900000 ;
        RECT 61.405000 36.140000 61.605000 36.340000 ;
        RECT 61.405000 36.580000 61.605000 36.780000 ;
        RECT 61.405000 37.020000 61.605000 37.220000 ;
        RECT 61.405000 37.460000 61.605000 37.660000 ;
        RECT 61.405000 37.900000 61.605000 38.100000 ;
        RECT 61.405000 49.715000 61.605000 49.915000 ;
        RECT 61.405000 50.135000 61.605000 50.335000 ;
        RECT 61.405000 50.555000 61.605000 50.755000 ;
        RECT 61.810000 34.820000 62.010000 35.020000 ;
        RECT 61.810000 35.260000 62.010000 35.460000 ;
        RECT 61.810000 35.700000 62.010000 35.900000 ;
        RECT 61.810000 36.140000 62.010000 36.340000 ;
        RECT 61.810000 36.580000 62.010000 36.780000 ;
        RECT 61.810000 37.020000 62.010000 37.220000 ;
        RECT 61.810000 37.460000 62.010000 37.660000 ;
        RECT 61.810000 37.900000 62.010000 38.100000 ;
        RECT 61.810000 49.715000 62.010000 49.915000 ;
        RECT 61.810000 50.135000 62.010000 50.335000 ;
        RECT 61.810000 50.555000 62.010000 50.755000 ;
        RECT 62.215000 34.820000 62.415000 35.020000 ;
        RECT 62.215000 35.260000 62.415000 35.460000 ;
        RECT 62.215000 35.700000 62.415000 35.900000 ;
        RECT 62.215000 36.140000 62.415000 36.340000 ;
        RECT 62.215000 36.580000 62.415000 36.780000 ;
        RECT 62.215000 37.020000 62.415000 37.220000 ;
        RECT 62.215000 37.460000 62.415000 37.660000 ;
        RECT 62.215000 37.900000 62.415000 38.100000 ;
        RECT 62.215000 49.715000 62.415000 49.915000 ;
        RECT 62.215000 50.135000 62.415000 50.335000 ;
        RECT 62.215000 50.555000 62.415000 50.755000 ;
        RECT 62.620000 34.820000 62.820000 35.020000 ;
        RECT 62.620000 35.260000 62.820000 35.460000 ;
        RECT 62.620000 35.700000 62.820000 35.900000 ;
        RECT 62.620000 36.140000 62.820000 36.340000 ;
        RECT 62.620000 36.580000 62.820000 36.780000 ;
        RECT 62.620000 37.020000 62.820000 37.220000 ;
        RECT 62.620000 37.460000 62.820000 37.660000 ;
        RECT 62.620000 37.900000 62.820000 38.100000 ;
        RECT 62.620000 49.715000 62.820000 49.915000 ;
        RECT 62.620000 50.135000 62.820000 50.335000 ;
        RECT 62.620000 50.555000 62.820000 50.755000 ;
        RECT 63.025000 34.820000 63.225000 35.020000 ;
        RECT 63.025000 35.260000 63.225000 35.460000 ;
        RECT 63.025000 35.700000 63.225000 35.900000 ;
        RECT 63.025000 36.140000 63.225000 36.340000 ;
        RECT 63.025000 36.580000 63.225000 36.780000 ;
        RECT 63.025000 37.020000 63.225000 37.220000 ;
        RECT 63.025000 37.460000 63.225000 37.660000 ;
        RECT 63.025000 37.900000 63.225000 38.100000 ;
        RECT 63.025000 49.715000 63.225000 49.915000 ;
        RECT 63.025000 50.135000 63.225000 50.335000 ;
        RECT 63.025000 50.555000 63.225000 50.755000 ;
        RECT 63.430000 34.820000 63.630000 35.020000 ;
        RECT 63.430000 35.260000 63.630000 35.460000 ;
        RECT 63.430000 35.700000 63.630000 35.900000 ;
        RECT 63.430000 36.140000 63.630000 36.340000 ;
        RECT 63.430000 36.580000 63.630000 36.780000 ;
        RECT 63.430000 37.020000 63.630000 37.220000 ;
        RECT 63.430000 37.460000 63.630000 37.660000 ;
        RECT 63.430000 37.900000 63.630000 38.100000 ;
        RECT 63.430000 49.715000 63.630000 49.915000 ;
        RECT 63.430000 50.135000 63.630000 50.335000 ;
        RECT 63.430000 50.555000 63.630000 50.755000 ;
        RECT 63.835000 34.820000 64.035000 35.020000 ;
        RECT 63.835000 35.260000 64.035000 35.460000 ;
        RECT 63.835000 35.700000 64.035000 35.900000 ;
        RECT 63.835000 36.140000 64.035000 36.340000 ;
        RECT 63.835000 36.580000 64.035000 36.780000 ;
        RECT 63.835000 37.020000 64.035000 37.220000 ;
        RECT 63.835000 37.460000 64.035000 37.660000 ;
        RECT 63.835000 37.900000 64.035000 38.100000 ;
        RECT 63.835000 49.715000 64.035000 49.915000 ;
        RECT 63.835000 50.135000 64.035000 50.335000 ;
        RECT 63.835000 50.555000 64.035000 50.755000 ;
        RECT 64.240000 34.820000 64.440000 35.020000 ;
        RECT 64.240000 35.260000 64.440000 35.460000 ;
        RECT 64.240000 35.700000 64.440000 35.900000 ;
        RECT 64.240000 36.140000 64.440000 36.340000 ;
        RECT 64.240000 36.580000 64.440000 36.780000 ;
        RECT 64.240000 37.020000 64.440000 37.220000 ;
        RECT 64.240000 37.460000 64.440000 37.660000 ;
        RECT 64.240000 37.900000 64.440000 38.100000 ;
        RECT 64.240000 49.715000 64.440000 49.915000 ;
        RECT 64.240000 50.135000 64.440000 50.335000 ;
        RECT 64.240000 50.555000 64.440000 50.755000 ;
        RECT 64.645000 34.820000 64.845000 35.020000 ;
        RECT 64.645000 35.260000 64.845000 35.460000 ;
        RECT 64.645000 35.700000 64.845000 35.900000 ;
        RECT 64.645000 36.140000 64.845000 36.340000 ;
        RECT 64.645000 36.580000 64.845000 36.780000 ;
        RECT 64.645000 37.020000 64.845000 37.220000 ;
        RECT 64.645000 37.460000 64.845000 37.660000 ;
        RECT 64.645000 37.900000 64.845000 38.100000 ;
        RECT 64.645000 49.715000 64.845000 49.915000 ;
        RECT 64.645000 50.135000 64.845000 50.335000 ;
        RECT 64.645000 50.555000 64.845000 50.755000 ;
        RECT 65.050000 34.820000 65.250000 35.020000 ;
        RECT 65.050000 35.260000 65.250000 35.460000 ;
        RECT 65.050000 35.700000 65.250000 35.900000 ;
        RECT 65.050000 36.140000 65.250000 36.340000 ;
        RECT 65.050000 36.580000 65.250000 36.780000 ;
        RECT 65.050000 37.020000 65.250000 37.220000 ;
        RECT 65.050000 37.460000 65.250000 37.660000 ;
        RECT 65.050000 37.900000 65.250000 38.100000 ;
        RECT 65.050000 49.715000 65.250000 49.915000 ;
        RECT 65.050000 50.135000 65.250000 50.335000 ;
        RECT 65.050000 50.555000 65.250000 50.755000 ;
        RECT 65.455000 34.820000 65.655000 35.020000 ;
        RECT 65.455000 35.260000 65.655000 35.460000 ;
        RECT 65.455000 35.700000 65.655000 35.900000 ;
        RECT 65.455000 36.140000 65.655000 36.340000 ;
        RECT 65.455000 36.580000 65.655000 36.780000 ;
        RECT 65.455000 37.020000 65.655000 37.220000 ;
        RECT 65.455000 37.460000 65.655000 37.660000 ;
        RECT 65.455000 37.900000 65.655000 38.100000 ;
        RECT 65.455000 49.715000 65.655000 49.915000 ;
        RECT 65.455000 50.135000 65.655000 50.335000 ;
        RECT 65.455000 50.555000 65.655000 50.755000 ;
        RECT 65.860000 34.820000 66.060000 35.020000 ;
        RECT 65.860000 35.260000 66.060000 35.460000 ;
        RECT 65.860000 35.700000 66.060000 35.900000 ;
        RECT 65.860000 36.140000 66.060000 36.340000 ;
        RECT 65.860000 36.580000 66.060000 36.780000 ;
        RECT 65.860000 37.020000 66.060000 37.220000 ;
        RECT 65.860000 37.460000 66.060000 37.660000 ;
        RECT 65.860000 37.900000 66.060000 38.100000 ;
        RECT 65.860000 49.715000 66.060000 49.915000 ;
        RECT 65.860000 50.135000 66.060000 50.335000 ;
        RECT 65.860000 50.555000 66.060000 50.755000 ;
        RECT 66.265000 34.820000 66.465000 35.020000 ;
        RECT 66.265000 35.260000 66.465000 35.460000 ;
        RECT 66.265000 35.700000 66.465000 35.900000 ;
        RECT 66.265000 36.140000 66.465000 36.340000 ;
        RECT 66.265000 36.580000 66.465000 36.780000 ;
        RECT 66.265000 37.020000 66.465000 37.220000 ;
        RECT 66.265000 37.460000 66.465000 37.660000 ;
        RECT 66.265000 37.900000 66.465000 38.100000 ;
        RECT 66.265000 49.715000 66.465000 49.915000 ;
        RECT 66.265000 50.135000 66.465000 50.335000 ;
        RECT 66.265000 50.555000 66.465000 50.755000 ;
        RECT 66.670000 34.820000 66.870000 35.020000 ;
        RECT 66.670000 35.260000 66.870000 35.460000 ;
        RECT 66.670000 35.700000 66.870000 35.900000 ;
        RECT 66.670000 36.140000 66.870000 36.340000 ;
        RECT 66.670000 36.580000 66.870000 36.780000 ;
        RECT 66.670000 37.020000 66.870000 37.220000 ;
        RECT 66.670000 37.460000 66.870000 37.660000 ;
        RECT 66.670000 37.900000 66.870000 38.100000 ;
        RECT 66.670000 49.715000 66.870000 49.915000 ;
        RECT 66.670000 50.135000 66.870000 50.335000 ;
        RECT 66.670000 50.555000 66.870000 50.755000 ;
        RECT 67.075000 34.820000 67.275000 35.020000 ;
        RECT 67.075000 35.260000 67.275000 35.460000 ;
        RECT 67.075000 35.700000 67.275000 35.900000 ;
        RECT 67.075000 36.140000 67.275000 36.340000 ;
        RECT 67.075000 36.580000 67.275000 36.780000 ;
        RECT 67.075000 37.020000 67.275000 37.220000 ;
        RECT 67.075000 37.460000 67.275000 37.660000 ;
        RECT 67.075000 37.900000 67.275000 38.100000 ;
        RECT 67.075000 49.715000 67.275000 49.915000 ;
        RECT 67.075000 50.135000 67.275000 50.335000 ;
        RECT 67.075000 50.555000 67.275000 50.755000 ;
        RECT 67.480000 34.820000 67.680000 35.020000 ;
        RECT 67.480000 35.260000 67.680000 35.460000 ;
        RECT 67.480000 35.700000 67.680000 35.900000 ;
        RECT 67.480000 36.140000 67.680000 36.340000 ;
        RECT 67.480000 36.580000 67.680000 36.780000 ;
        RECT 67.480000 37.020000 67.680000 37.220000 ;
        RECT 67.480000 37.460000 67.680000 37.660000 ;
        RECT 67.480000 37.900000 67.680000 38.100000 ;
        RECT 67.480000 49.715000 67.680000 49.915000 ;
        RECT 67.480000 50.135000 67.680000 50.335000 ;
        RECT 67.480000 50.555000 67.680000 50.755000 ;
        RECT 67.885000 34.820000 68.085000 35.020000 ;
        RECT 67.885000 35.260000 68.085000 35.460000 ;
        RECT 67.885000 35.700000 68.085000 35.900000 ;
        RECT 67.885000 36.140000 68.085000 36.340000 ;
        RECT 67.885000 36.580000 68.085000 36.780000 ;
        RECT 67.885000 37.020000 68.085000 37.220000 ;
        RECT 67.885000 37.460000 68.085000 37.660000 ;
        RECT 67.885000 37.900000 68.085000 38.100000 ;
        RECT 67.885000 49.715000 68.085000 49.915000 ;
        RECT 67.885000 50.135000 68.085000 50.335000 ;
        RECT 67.885000 50.555000 68.085000 50.755000 ;
        RECT 68.290000 34.820000 68.490000 35.020000 ;
        RECT 68.290000 35.260000 68.490000 35.460000 ;
        RECT 68.290000 35.700000 68.490000 35.900000 ;
        RECT 68.290000 36.140000 68.490000 36.340000 ;
        RECT 68.290000 36.580000 68.490000 36.780000 ;
        RECT 68.290000 37.020000 68.490000 37.220000 ;
        RECT 68.290000 37.460000 68.490000 37.660000 ;
        RECT 68.290000 37.900000 68.490000 38.100000 ;
        RECT 68.290000 49.715000 68.490000 49.915000 ;
        RECT 68.290000 50.135000 68.490000 50.335000 ;
        RECT 68.290000 50.555000 68.490000 50.755000 ;
        RECT 68.695000 34.820000 68.895000 35.020000 ;
        RECT 68.695000 35.260000 68.895000 35.460000 ;
        RECT 68.695000 35.700000 68.895000 35.900000 ;
        RECT 68.695000 36.140000 68.895000 36.340000 ;
        RECT 68.695000 36.580000 68.895000 36.780000 ;
        RECT 68.695000 37.020000 68.895000 37.220000 ;
        RECT 68.695000 37.460000 68.895000 37.660000 ;
        RECT 68.695000 37.900000 68.895000 38.100000 ;
        RECT 68.695000 49.715000 68.895000 49.915000 ;
        RECT 68.695000 50.135000 68.895000 50.335000 ;
        RECT 68.695000 50.555000 68.895000 50.755000 ;
        RECT 69.100000 34.820000 69.300000 35.020000 ;
        RECT 69.100000 35.260000 69.300000 35.460000 ;
        RECT 69.100000 35.700000 69.300000 35.900000 ;
        RECT 69.100000 36.140000 69.300000 36.340000 ;
        RECT 69.100000 36.580000 69.300000 36.780000 ;
        RECT 69.100000 37.020000 69.300000 37.220000 ;
        RECT 69.100000 37.460000 69.300000 37.660000 ;
        RECT 69.100000 37.900000 69.300000 38.100000 ;
        RECT 69.100000 49.715000 69.300000 49.915000 ;
        RECT 69.100000 50.135000 69.300000 50.335000 ;
        RECT 69.100000 50.555000 69.300000 50.755000 ;
        RECT 69.505000 34.820000 69.705000 35.020000 ;
        RECT 69.505000 35.260000 69.705000 35.460000 ;
        RECT 69.505000 35.700000 69.705000 35.900000 ;
        RECT 69.505000 36.140000 69.705000 36.340000 ;
        RECT 69.505000 36.580000 69.705000 36.780000 ;
        RECT 69.505000 37.020000 69.705000 37.220000 ;
        RECT 69.505000 37.460000 69.705000 37.660000 ;
        RECT 69.505000 37.900000 69.705000 38.100000 ;
        RECT 69.505000 49.715000 69.705000 49.915000 ;
        RECT 69.505000 50.135000 69.705000 50.335000 ;
        RECT 69.505000 50.555000 69.705000 50.755000 ;
        RECT 69.910000 34.820000 70.110000 35.020000 ;
        RECT 69.910000 35.260000 70.110000 35.460000 ;
        RECT 69.910000 35.700000 70.110000 35.900000 ;
        RECT 69.910000 36.140000 70.110000 36.340000 ;
        RECT 69.910000 36.580000 70.110000 36.780000 ;
        RECT 69.910000 37.020000 70.110000 37.220000 ;
        RECT 69.910000 37.460000 70.110000 37.660000 ;
        RECT 69.910000 37.900000 70.110000 38.100000 ;
        RECT 69.910000 49.715000 70.110000 49.915000 ;
        RECT 69.910000 50.135000 70.110000 50.335000 ;
        RECT 69.910000 50.555000 70.110000 50.755000 ;
        RECT 70.315000 34.820000 70.515000 35.020000 ;
        RECT 70.315000 35.260000 70.515000 35.460000 ;
        RECT 70.315000 35.700000 70.515000 35.900000 ;
        RECT 70.315000 36.140000 70.515000 36.340000 ;
        RECT 70.315000 36.580000 70.515000 36.780000 ;
        RECT 70.315000 37.020000 70.515000 37.220000 ;
        RECT 70.315000 37.460000 70.515000 37.660000 ;
        RECT 70.315000 37.900000 70.515000 38.100000 ;
        RECT 70.315000 49.715000 70.515000 49.915000 ;
        RECT 70.315000 50.135000 70.515000 50.335000 ;
        RECT 70.315000 50.555000 70.515000 50.755000 ;
        RECT 70.720000 34.820000 70.920000 35.020000 ;
        RECT 70.720000 35.260000 70.920000 35.460000 ;
        RECT 70.720000 35.700000 70.920000 35.900000 ;
        RECT 70.720000 36.140000 70.920000 36.340000 ;
        RECT 70.720000 36.580000 70.920000 36.780000 ;
        RECT 70.720000 37.020000 70.920000 37.220000 ;
        RECT 70.720000 37.460000 70.920000 37.660000 ;
        RECT 70.720000 37.900000 70.920000 38.100000 ;
        RECT 70.720000 49.715000 70.920000 49.915000 ;
        RECT 70.720000 50.135000 70.920000 50.335000 ;
        RECT 70.720000 50.555000 70.920000 50.755000 ;
        RECT 71.125000 34.820000 71.325000 35.020000 ;
        RECT 71.125000 35.260000 71.325000 35.460000 ;
        RECT 71.125000 35.700000 71.325000 35.900000 ;
        RECT 71.125000 36.140000 71.325000 36.340000 ;
        RECT 71.125000 36.580000 71.325000 36.780000 ;
        RECT 71.125000 37.020000 71.325000 37.220000 ;
        RECT 71.125000 37.460000 71.325000 37.660000 ;
        RECT 71.125000 37.900000 71.325000 38.100000 ;
        RECT 71.125000 49.715000 71.325000 49.915000 ;
        RECT 71.125000 50.135000 71.325000 50.335000 ;
        RECT 71.125000 50.555000 71.325000 50.755000 ;
        RECT 71.530000 34.820000 71.730000 35.020000 ;
        RECT 71.530000 35.260000 71.730000 35.460000 ;
        RECT 71.530000 35.700000 71.730000 35.900000 ;
        RECT 71.530000 36.140000 71.730000 36.340000 ;
        RECT 71.530000 36.580000 71.730000 36.780000 ;
        RECT 71.530000 37.020000 71.730000 37.220000 ;
        RECT 71.530000 37.460000 71.730000 37.660000 ;
        RECT 71.530000 37.900000 71.730000 38.100000 ;
        RECT 71.530000 49.715000 71.730000 49.915000 ;
        RECT 71.530000 50.135000 71.730000 50.335000 ;
        RECT 71.530000 50.555000 71.730000 50.755000 ;
        RECT 71.935000 34.820000 72.135000 35.020000 ;
        RECT 71.935000 35.260000 72.135000 35.460000 ;
        RECT 71.935000 35.700000 72.135000 35.900000 ;
        RECT 71.935000 36.140000 72.135000 36.340000 ;
        RECT 71.935000 36.580000 72.135000 36.780000 ;
        RECT 71.935000 37.020000 72.135000 37.220000 ;
        RECT 71.935000 37.460000 72.135000 37.660000 ;
        RECT 71.935000 37.900000 72.135000 38.100000 ;
        RECT 71.935000 49.715000 72.135000 49.915000 ;
        RECT 71.935000 50.135000 72.135000 50.335000 ;
        RECT 71.935000 50.555000 72.135000 50.755000 ;
        RECT 72.340000 34.820000 72.540000 35.020000 ;
        RECT 72.340000 35.260000 72.540000 35.460000 ;
        RECT 72.340000 35.700000 72.540000 35.900000 ;
        RECT 72.340000 36.140000 72.540000 36.340000 ;
        RECT 72.340000 36.580000 72.540000 36.780000 ;
        RECT 72.340000 37.020000 72.540000 37.220000 ;
        RECT 72.340000 37.460000 72.540000 37.660000 ;
        RECT 72.340000 37.900000 72.540000 38.100000 ;
        RECT 72.340000 49.715000 72.540000 49.915000 ;
        RECT 72.340000 50.135000 72.540000 50.335000 ;
        RECT 72.340000 50.555000 72.540000 50.755000 ;
        RECT 72.745000 34.820000 72.945000 35.020000 ;
        RECT 72.745000 35.260000 72.945000 35.460000 ;
        RECT 72.745000 35.700000 72.945000 35.900000 ;
        RECT 72.745000 36.140000 72.945000 36.340000 ;
        RECT 72.745000 36.580000 72.945000 36.780000 ;
        RECT 72.745000 37.020000 72.945000 37.220000 ;
        RECT 72.745000 37.460000 72.945000 37.660000 ;
        RECT 72.745000 37.900000 72.945000 38.100000 ;
        RECT 72.745000 49.715000 72.945000 49.915000 ;
        RECT 72.745000 50.135000 72.945000 50.335000 ;
        RECT 72.745000 50.555000 72.945000 50.755000 ;
        RECT 73.150000 34.820000 73.350000 35.020000 ;
        RECT 73.150000 35.260000 73.350000 35.460000 ;
        RECT 73.150000 35.700000 73.350000 35.900000 ;
        RECT 73.150000 36.140000 73.350000 36.340000 ;
        RECT 73.150000 36.580000 73.350000 36.780000 ;
        RECT 73.150000 37.020000 73.350000 37.220000 ;
        RECT 73.150000 37.460000 73.350000 37.660000 ;
        RECT 73.150000 37.900000 73.350000 38.100000 ;
        RECT 73.150000 49.715000 73.350000 49.915000 ;
        RECT 73.150000 50.135000 73.350000 50.335000 ;
        RECT 73.150000 50.555000 73.350000 50.755000 ;
        RECT 73.555000 34.820000 73.755000 35.020000 ;
        RECT 73.555000 35.260000 73.755000 35.460000 ;
        RECT 73.555000 35.700000 73.755000 35.900000 ;
        RECT 73.555000 36.140000 73.755000 36.340000 ;
        RECT 73.555000 36.580000 73.755000 36.780000 ;
        RECT 73.555000 37.020000 73.755000 37.220000 ;
        RECT 73.555000 37.460000 73.755000 37.660000 ;
        RECT 73.555000 37.900000 73.755000 38.100000 ;
        RECT 73.555000 49.715000 73.755000 49.915000 ;
        RECT 73.555000 50.135000 73.755000 50.335000 ;
        RECT 73.555000 50.555000 73.755000 50.755000 ;
        RECT 73.960000 34.820000 74.160000 35.020000 ;
        RECT 73.960000 35.260000 74.160000 35.460000 ;
        RECT 73.960000 35.700000 74.160000 35.900000 ;
        RECT 73.960000 36.140000 74.160000 36.340000 ;
        RECT 73.960000 36.580000 74.160000 36.780000 ;
        RECT 73.960000 37.020000 74.160000 37.220000 ;
        RECT 73.960000 37.460000 74.160000 37.660000 ;
        RECT 73.960000 37.900000 74.160000 38.100000 ;
        RECT 73.960000 49.715000 74.160000 49.915000 ;
        RECT 73.960000 50.135000 74.160000 50.335000 ;
        RECT 73.960000 50.555000 74.160000 50.755000 ;
        RECT 74.365000 34.820000 74.565000 35.020000 ;
        RECT 74.365000 35.260000 74.565000 35.460000 ;
        RECT 74.365000 35.700000 74.565000 35.900000 ;
        RECT 74.365000 36.140000 74.565000 36.340000 ;
        RECT 74.365000 36.580000 74.565000 36.780000 ;
        RECT 74.365000 37.020000 74.565000 37.220000 ;
        RECT 74.365000 37.460000 74.565000 37.660000 ;
        RECT 74.365000 37.900000 74.565000 38.100000 ;
        RECT 74.365000 49.715000 74.565000 49.915000 ;
        RECT 74.365000 50.135000 74.565000 50.335000 ;
        RECT 74.365000 50.555000 74.565000 50.755000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 75.000000  34.340000 ;
      RECT  0.000000 38.580000 75.000000  49.250000 ;
      RECT  0.000000 51.220000 75.000000 198.000000 ;
      RECT 24.800000  0.000000 50.355000 198.000000 ;
      RECT 24.800000  0.000000 50.355000 198.000000 ;
      RECT 24.800000 34.340000 50.355000  38.580000 ;
      RECT 24.800000 49.250000 50.355000  51.220000 ;
    LAYER met4 ;
      RECT  0.000000   5.885000  1.670000   6.485000 ;
      RECT  0.000000  11.935000  1.365000  12.535000 ;
      RECT  0.000000  16.785000  1.365000  17.385000 ;
      RECT  0.000000  22.835000  1.670000  23.435000 ;
      RECT  0.000000  28.885000  1.670000  29.485000 ;
      RECT  0.000000  33.735000  1.670000  34.335000 ;
      RECT  0.000000  38.585000  1.670000  39.185000 ;
      RECT  0.000000  44.635000  1.670000  45.335000 ;
      RECT  0.000000  55.135000  1.670000  55.835000 ;
      RECT  0.000000  61.085000  1.670000  61.685000 ;
      RECT  0.000000  66.935000  1.670000  67.635000 ;
      RECT  0.000000  93.400000 75.000000 173.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.670000   0.000000 73.330000  11.935000 ;
      RECT  1.670000   0.000000 73.330000  34.335000 ;
      RECT  1.670000   0.000000 73.330000  34.335000 ;
      RECT  1.670000   0.000000 73.330000  34.335000 ;
      RECT  1.670000   0.000000 73.330000  34.335000 ;
      RECT  1.670000   0.000000 73.330000  34.335000 ;
      RECT  1.670000  17.385000 73.330000  34.335000 ;
      RECT  1.670000  38.585000 73.330000  49.245000 ;
      RECT  1.670000  38.585000 73.330000  49.245000 ;
      RECT  1.670000  38.585000 73.330000  49.245000 ;
      RECT  1.670000  51.225000 73.330000  93.400000 ;
      RECT  1.670000  51.225000 73.330000 198.000000 ;
      RECT  1.670000  51.225000 73.330000 198.000000 ;
      RECT  1.670000  51.225000 73.330000 198.000000 ;
      RECT  1.670000  51.225000 73.330000 198.000000 ;
      RECT  1.670000  51.225000 73.330000 198.000000 ;
      RECT  1.670000 173.385000 73.330000 198.000000 ;
      RECT 24.775000   0.000000 50.380000  51.225000 ;
      RECT 24.775000   0.000000 50.380000 198.000000 ;
      RECT 24.775000  34.335000 50.380000  38.585000 ;
      RECT 24.775000  49.245000 50.380000  51.225000 ;
      RECT 73.330000   5.885000 75.000000   6.485000 ;
      RECT 73.330000  22.835000 75.000000  23.435000 ;
      RECT 73.330000  28.885000 75.000000  29.485000 ;
      RECT 73.330000  33.735000 75.000000  34.335000 ;
      RECT 73.330000  38.585000 75.000000  39.185000 ;
      RECT 73.330000  44.635000 75.000000  45.335000 ;
      RECT 73.330000  55.135000 75.000000  55.835000 ;
      RECT 73.330000  61.085000 75.000000  61.685000 ;
      RECT 73.330000  66.935000 75.000000  67.635000 ;
      RECT 73.635000  11.935000 75.000000  12.535000 ;
      RECT 73.635000  16.785000 75.000000  17.385000 ;
    LAYER met5 ;
      RECT 0.000000  93.785000 75.000000 172.985000 ;
      RECT 1.765000  12.235000 73.235000  17.085000 ;
      RECT 2.070000   0.000000 72.930000  12.235000 ;
      RECT 2.070000  17.085000 72.930000  93.785000 ;
      RECT 2.070000 172.985000 72.930000 198.000000 ;
  END
END sky130_fd_io__overlay_vssa_lvc


MACRO sky130_fd_io__overlay_vccd_hvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.495000 8.890000 24.395000 13.530000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 8.890000 74.290000 13.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 24.370000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.585000  8.960000  0.785000  9.160000 ;
        RECT  0.585000  9.390000  0.785000  9.590000 ;
        RECT  0.585000  9.820000  0.785000 10.020000 ;
        RECT  0.585000 10.250000  0.785000 10.450000 ;
        RECT  0.585000 10.680000  0.785000 10.880000 ;
        RECT  0.585000 11.110000  0.785000 11.310000 ;
        RECT  0.585000 11.540000  0.785000 11.740000 ;
        RECT  0.585000 11.970000  0.785000 12.170000 ;
        RECT  0.585000 12.400000  0.785000 12.600000 ;
        RECT  0.585000 12.830000  0.785000 13.030000 ;
        RECT  0.585000 13.260000  0.785000 13.460000 ;
        RECT  0.995000  8.960000  1.195000  9.160000 ;
        RECT  0.995000  9.390000  1.195000  9.590000 ;
        RECT  0.995000  9.820000  1.195000 10.020000 ;
        RECT  0.995000 10.250000  1.195000 10.450000 ;
        RECT  0.995000 10.680000  1.195000 10.880000 ;
        RECT  0.995000 11.110000  1.195000 11.310000 ;
        RECT  0.995000 11.540000  1.195000 11.740000 ;
        RECT  0.995000 11.970000  1.195000 12.170000 ;
        RECT  0.995000 12.400000  1.195000 12.600000 ;
        RECT  0.995000 12.830000  1.195000 13.030000 ;
        RECT  0.995000 13.260000  1.195000 13.460000 ;
        RECT  1.405000  8.960000  1.605000  9.160000 ;
        RECT  1.405000  9.390000  1.605000  9.590000 ;
        RECT  1.405000  9.820000  1.605000 10.020000 ;
        RECT  1.405000 10.250000  1.605000 10.450000 ;
        RECT  1.405000 10.680000  1.605000 10.880000 ;
        RECT  1.405000 11.110000  1.605000 11.310000 ;
        RECT  1.405000 11.540000  1.605000 11.740000 ;
        RECT  1.405000 11.970000  1.605000 12.170000 ;
        RECT  1.405000 12.400000  1.605000 12.600000 ;
        RECT  1.405000 12.830000  1.605000 13.030000 ;
        RECT  1.405000 13.260000  1.605000 13.460000 ;
        RECT  1.815000  8.960000  2.015000  9.160000 ;
        RECT  1.815000  9.390000  2.015000  9.590000 ;
        RECT  1.815000  9.820000  2.015000 10.020000 ;
        RECT  1.815000 10.250000  2.015000 10.450000 ;
        RECT  1.815000 10.680000  2.015000 10.880000 ;
        RECT  1.815000 11.110000  2.015000 11.310000 ;
        RECT  1.815000 11.540000  2.015000 11.740000 ;
        RECT  1.815000 11.970000  2.015000 12.170000 ;
        RECT  1.815000 12.400000  2.015000 12.600000 ;
        RECT  1.815000 12.830000  2.015000 13.030000 ;
        RECT  1.815000 13.260000  2.015000 13.460000 ;
        RECT  2.225000  8.960000  2.425000  9.160000 ;
        RECT  2.225000  9.390000  2.425000  9.590000 ;
        RECT  2.225000  9.820000  2.425000 10.020000 ;
        RECT  2.225000 10.250000  2.425000 10.450000 ;
        RECT  2.225000 10.680000  2.425000 10.880000 ;
        RECT  2.225000 11.110000  2.425000 11.310000 ;
        RECT  2.225000 11.540000  2.425000 11.740000 ;
        RECT  2.225000 11.970000  2.425000 12.170000 ;
        RECT  2.225000 12.400000  2.425000 12.600000 ;
        RECT  2.225000 12.830000  2.425000 13.030000 ;
        RECT  2.225000 13.260000  2.425000 13.460000 ;
        RECT  2.635000  8.960000  2.835000  9.160000 ;
        RECT  2.635000  9.390000  2.835000  9.590000 ;
        RECT  2.635000  9.820000  2.835000 10.020000 ;
        RECT  2.635000 10.250000  2.835000 10.450000 ;
        RECT  2.635000 10.680000  2.835000 10.880000 ;
        RECT  2.635000 11.110000  2.835000 11.310000 ;
        RECT  2.635000 11.540000  2.835000 11.740000 ;
        RECT  2.635000 11.970000  2.835000 12.170000 ;
        RECT  2.635000 12.400000  2.835000 12.600000 ;
        RECT  2.635000 12.830000  2.835000 13.030000 ;
        RECT  2.635000 13.260000  2.835000 13.460000 ;
        RECT  3.045000  8.960000  3.245000  9.160000 ;
        RECT  3.045000  9.390000  3.245000  9.590000 ;
        RECT  3.045000  9.820000  3.245000 10.020000 ;
        RECT  3.045000 10.250000  3.245000 10.450000 ;
        RECT  3.045000 10.680000  3.245000 10.880000 ;
        RECT  3.045000 11.110000  3.245000 11.310000 ;
        RECT  3.045000 11.540000  3.245000 11.740000 ;
        RECT  3.045000 11.970000  3.245000 12.170000 ;
        RECT  3.045000 12.400000  3.245000 12.600000 ;
        RECT  3.045000 12.830000  3.245000 13.030000 ;
        RECT  3.045000 13.260000  3.245000 13.460000 ;
        RECT  3.450000  8.960000  3.650000  9.160000 ;
        RECT  3.450000  9.390000  3.650000  9.590000 ;
        RECT  3.450000  9.820000  3.650000 10.020000 ;
        RECT  3.450000 10.250000  3.650000 10.450000 ;
        RECT  3.450000 10.680000  3.650000 10.880000 ;
        RECT  3.450000 11.110000  3.650000 11.310000 ;
        RECT  3.450000 11.540000  3.650000 11.740000 ;
        RECT  3.450000 11.970000  3.650000 12.170000 ;
        RECT  3.450000 12.400000  3.650000 12.600000 ;
        RECT  3.450000 12.830000  3.650000 13.030000 ;
        RECT  3.450000 13.260000  3.650000 13.460000 ;
        RECT  3.855000  8.960000  4.055000  9.160000 ;
        RECT  3.855000  9.390000  4.055000  9.590000 ;
        RECT  3.855000  9.820000  4.055000 10.020000 ;
        RECT  3.855000 10.250000  4.055000 10.450000 ;
        RECT  3.855000 10.680000  4.055000 10.880000 ;
        RECT  3.855000 11.110000  4.055000 11.310000 ;
        RECT  3.855000 11.540000  4.055000 11.740000 ;
        RECT  3.855000 11.970000  4.055000 12.170000 ;
        RECT  3.855000 12.400000  4.055000 12.600000 ;
        RECT  3.855000 12.830000  4.055000 13.030000 ;
        RECT  3.855000 13.260000  4.055000 13.460000 ;
        RECT  4.260000  8.960000  4.460000  9.160000 ;
        RECT  4.260000  9.390000  4.460000  9.590000 ;
        RECT  4.260000  9.820000  4.460000 10.020000 ;
        RECT  4.260000 10.250000  4.460000 10.450000 ;
        RECT  4.260000 10.680000  4.460000 10.880000 ;
        RECT  4.260000 11.110000  4.460000 11.310000 ;
        RECT  4.260000 11.540000  4.460000 11.740000 ;
        RECT  4.260000 11.970000  4.460000 12.170000 ;
        RECT  4.260000 12.400000  4.460000 12.600000 ;
        RECT  4.260000 12.830000  4.460000 13.030000 ;
        RECT  4.260000 13.260000  4.460000 13.460000 ;
        RECT  4.665000  8.960000  4.865000  9.160000 ;
        RECT  4.665000  9.390000  4.865000  9.590000 ;
        RECT  4.665000  9.820000  4.865000 10.020000 ;
        RECT  4.665000 10.250000  4.865000 10.450000 ;
        RECT  4.665000 10.680000  4.865000 10.880000 ;
        RECT  4.665000 11.110000  4.865000 11.310000 ;
        RECT  4.665000 11.540000  4.865000 11.740000 ;
        RECT  4.665000 11.970000  4.865000 12.170000 ;
        RECT  4.665000 12.400000  4.865000 12.600000 ;
        RECT  4.665000 12.830000  4.865000 13.030000 ;
        RECT  4.665000 13.260000  4.865000 13.460000 ;
        RECT  5.070000  8.960000  5.270000  9.160000 ;
        RECT  5.070000  9.390000  5.270000  9.590000 ;
        RECT  5.070000  9.820000  5.270000 10.020000 ;
        RECT  5.070000 10.250000  5.270000 10.450000 ;
        RECT  5.070000 10.680000  5.270000 10.880000 ;
        RECT  5.070000 11.110000  5.270000 11.310000 ;
        RECT  5.070000 11.540000  5.270000 11.740000 ;
        RECT  5.070000 11.970000  5.270000 12.170000 ;
        RECT  5.070000 12.400000  5.270000 12.600000 ;
        RECT  5.070000 12.830000  5.270000 13.030000 ;
        RECT  5.070000 13.260000  5.270000 13.460000 ;
        RECT  5.475000  8.960000  5.675000  9.160000 ;
        RECT  5.475000  9.390000  5.675000  9.590000 ;
        RECT  5.475000  9.820000  5.675000 10.020000 ;
        RECT  5.475000 10.250000  5.675000 10.450000 ;
        RECT  5.475000 10.680000  5.675000 10.880000 ;
        RECT  5.475000 11.110000  5.675000 11.310000 ;
        RECT  5.475000 11.540000  5.675000 11.740000 ;
        RECT  5.475000 11.970000  5.675000 12.170000 ;
        RECT  5.475000 12.400000  5.675000 12.600000 ;
        RECT  5.475000 12.830000  5.675000 13.030000 ;
        RECT  5.475000 13.260000  5.675000 13.460000 ;
        RECT  5.880000  8.960000  6.080000  9.160000 ;
        RECT  5.880000  9.390000  6.080000  9.590000 ;
        RECT  5.880000  9.820000  6.080000 10.020000 ;
        RECT  5.880000 10.250000  6.080000 10.450000 ;
        RECT  5.880000 10.680000  6.080000 10.880000 ;
        RECT  5.880000 11.110000  6.080000 11.310000 ;
        RECT  5.880000 11.540000  6.080000 11.740000 ;
        RECT  5.880000 11.970000  6.080000 12.170000 ;
        RECT  5.880000 12.400000  6.080000 12.600000 ;
        RECT  5.880000 12.830000  6.080000 13.030000 ;
        RECT  5.880000 13.260000  6.080000 13.460000 ;
        RECT  6.285000  8.960000  6.485000  9.160000 ;
        RECT  6.285000  9.390000  6.485000  9.590000 ;
        RECT  6.285000  9.820000  6.485000 10.020000 ;
        RECT  6.285000 10.250000  6.485000 10.450000 ;
        RECT  6.285000 10.680000  6.485000 10.880000 ;
        RECT  6.285000 11.110000  6.485000 11.310000 ;
        RECT  6.285000 11.540000  6.485000 11.740000 ;
        RECT  6.285000 11.970000  6.485000 12.170000 ;
        RECT  6.285000 12.400000  6.485000 12.600000 ;
        RECT  6.285000 12.830000  6.485000 13.030000 ;
        RECT  6.285000 13.260000  6.485000 13.460000 ;
        RECT  6.690000  8.960000  6.890000  9.160000 ;
        RECT  6.690000  9.390000  6.890000  9.590000 ;
        RECT  6.690000  9.820000  6.890000 10.020000 ;
        RECT  6.690000 10.250000  6.890000 10.450000 ;
        RECT  6.690000 10.680000  6.890000 10.880000 ;
        RECT  6.690000 11.110000  6.890000 11.310000 ;
        RECT  6.690000 11.540000  6.890000 11.740000 ;
        RECT  6.690000 11.970000  6.890000 12.170000 ;
        RECT  6.690000 12.400000  6.890000 12.600000 ;
        RECT  6.690000 12.830000  6.890000 13.030000 ;
        RECT  6.690000 13.260000  6.890000 13.460000 ;
        RECT  7.095000  8.960000  7.295000  9.160000 ;
        RECT  7.095000  9.390000  7.295000  9.590000 ;
        RECT  7.095000  9.820000  7.295000 10.020000 ;
        RECT  7.095000 10.250000  7.295000 10.450000 ;
        RECT  7.095000 10.680000  7.295000 10.880000 ;
        RECT  7.095000 11.110000  7.295000 11.310000 ;
        RECT  7.095000 11.540000  7.295000 11.740000 ;
        RECT  7.095000 11.970000  7.295000 12.170000 ;
        RECT  7.095000 12.400000  7.295000 12.600000 ;
        RECT  7.095000 12.830000  7.295000 13.030000 ;
        RECT  7.095000 13.260000  7.295000 13.460000 ;
        RECT  7.500000  8.960000  7.700000  9.160000 ;
        RECT  7.500000  9.390000  7.700000  9.590000 ;
        RECT  7.500000  9.820000  7.700000 10.020000 ;
        RECT  7.500000 10.250000  7.700000 10.450000 ;
        RECT  7.500000 10.680000  7.700000 10.880000 ;
        RECT  7.500000 11.110000  7.700000 11.310000 ;
        RECT  7.500000 11.540000  7.700000 11.740000 ;
        RECT  7.500000 11.970000  7.700000 12.170000 ;
        RECT  7.500000 12.400000  7.700000 12.600000 ;
        RECT  7.500000 12.830000  7.700000 13.030000 ;
        RECT  7.500000 13.260000  7.700000 13.460000 ;
        RECT  7.905000  8.960000  8.105000  9.160000 ;
        RECT  7.905000  9.390000  8.105000  9.590000 ;
        RECT  7.905000  9.820000  8.105000 10.020000 ;
        RECT  7.905000 10.250000  8.105000 10.450000 ;
        RECT  7.905000 10.680000  8.105000 10.880000 ;
        RECT  7.905000 11.110000  8.105000 11.310000 ;
        RECT  7.905000 11.540000  8.105000 11.740000 ;
        RECT  7.905000 11.970000  8.105000 12.170000 ;
        RECT  7.905000 12.400000  8.105000 12.600000 ;
        RECT  7.905000 12.830000  8.105000 13.030000 ;
        RECT  7.905000 13.260000  8.105000 13.460000 ;
        RECT  8.310000  8.960000  8.510000  9.160000 ;
        RECT  8.310000  9.390000  8.510000  9.590000 ;
        RECT  8.310000  9.820000  8.510000 10.020000 ;
        RECT  8.310000 10.250000  8.510000 10.450000 ;
        RECT  8.310000 10.680000  8.510000 10.880000 ;
        RECT  8.310000 11.110000  8.510000 11.310000 ;
        RECT  8.310000 11.540000  8.510000 11.740000 ;
        RECT  8.310000 11.970000  8.510000 12.170000 ;
        RECT  8.310000 12.400000  8.510000 12.600000 ;
        RECT  8.310000 12.830000  8.510000 13.030000 ;
        RECT  8.310000 13.260000  8.510000 13.460000 ;
        RECT  8.715000  8.960000  8.915000  9.160000 ;
        RECT  8.715000  9.390000  8.915000  9.590000 ;
        RECT  8.715000  9.820000  8.915000 10.020000 ;
        RECT  8.715000 10.250000  8.915000 10.450000 ;
        RECT  8.715000 10.680000  8.915000 10.880000 ;
        RECT  8.715000 11.110000  8.915000 11.310000 ;
        RECT  8.715000 11.540000  8.915000 11.740000 ;
        RECT  8.715000 11.970000  8.915000 12.170000 ;
        RECT  8.715000 12.400000  8.915000 12.600000 ;
        RECT  8.715000 12.830000  8.915000 13.030000 ;
        RECT  8.715000 13.260000  8.915000 13.460000 ;
        RECT  9.120000  8.960000  9.320000  9.160000 ;
        RECT  9.120000  9.390000  9.320000  9.590000 ;
        RECT  9.120000  9.820000  9.320000 10.020000 ;
        RECT  9.120000 10.250000  9.320000 10.450000 ;
        RECT  9.120000 10.680000  9.320000 10.880000 ;
        RECT  9.120000 11.110000  9.320000 11.310000 ;
        RECT  9.120000 11.540000  9.320000 11.740000 ;
        RECT  9.120000 11.970000  9.320000 12.170000 ;
        RECT  9.120000 12.400000  9.320000 12.600000 ;
        RECT  9.120000 12.830000  9.320000 13.030000 ;
        RECT  9.120000 13.260000  9.320000 13.460000 ;
        RECT  9.525000  8.960000  9.725000  9.160000 ;
        RECT  9.525000  9.390000  9.725000  9.590000 ;
        RECT  9.525000  9.820000  9.725000 10.020000 ;
        RECT  9.525000 10.250000  9.725000 10.450000 ;
        RECT  9.525000 10.680000  9.725000 10.880000 ;
        RECT  9.525000 11.110000  9.725000 11.310000 ;
        RECT  9.525000 11.540000  9.725000 11.740000 ;
        RECT  9.525000 11.970000  9.725000 12.170000 ;
        RECT  9.525000 12.400000  9.725000 12.600000 ;
        RECT  9.525000 12.830000  9.725000 13.030000 ;
        RECT  9.525000 13.260000  9.725000 13.460000 ;
        RECT  9.930000  8.960000 10.130000  9.160000 ;
        RECT  9.930000  9.390000 10.130000  9.590000 ;
        RECT  9.930000  9.820000 10.130000 10.020000 ;
        RECT  9.930000 10.250000 10.130000 10.450000 ;
        RECT  9.930000 10.680000 10.130000 10.880000 ;
        RECT  9.930000 11.110000 10.130000 11.310000 ;
        RECT  9.930000 11.540000 10.130000 11.740000 ;
        RECT  9.930000 11.970000 10.130000 12.170000 ;
        RECT  9.930000 12.400000 10.130000 12.600000 ;
        RECT  9.930000 12.830000 10.130000 13.030000 ;
        RECT  9.930000 13.260000 10.130000 13.460000 ;
        RECT 10.335000  8.960000 10.535000  9.160000 ;
        RECT 10.335000  9.390000 10.535000  9.590000 ;
        RECT 10.335000  9.820000 10.535000 10.020000 ;
        RECT 10.335000 10.250000 10.535000 10.450000 ;
        RECT 10.335000 10.680000 10.535000 10.880000 ;
        RECT 10.335000 11.110000 10.535000 11.310000 ;
        RECT 10.335000 11.540000 10.535000 11.740000 ;
        RECT 10.335000 11.970000 10.535000 12.170000 ;
        RECT 10.335000 12.400000 10.535000 12.600000 ;
        RECT 10.335000 12.830000 10.535000 13.030000 ;
        RECT 10.335000 13.260000 10.535000 13.460000 ;
        RECT 10.740000  8.960000 10.940000  9.160000 ;
        RECT 10.740000  9.390000 10.940000  9.590000 ;
        RECT 10.740000  9.820000 10.940000 10.020000 ;
        RECT 10.740000 10.250000 10.940000 10.450000 ;
        RECT 10.740000 10.680000 10.940000 10.880000 ;
        RECT 10.740000 11.110000 10.940000 11.310000 ;
        RECT 10.740000 11.540000 10.940000 11.740000 ;
        RECT 10.740000 11.970000 10.940000 12.170000 ;
        RECT 10.740000 12.400000 10.940000 12.600000 ;
        RECT 10.740000 12.830000 10.940000 13.030000 ;
        RECT 10.740000 13.260000 10.940000 13.460000 ;
        RECT 11.145000  8.960000 11.345000  9.160000 ;
        RECT 11.145000  9.390000 11.345000  9.590000 ;
        RECT 11.145000  9.820000 11.345000 10.020000 ;
        RECT 11.145000 10.250000 11.345000 10.450000 ;
        RECT 11.145000 10.680000 11.345000 10.880000 ;
        RECT 11.145000 11.110000 11.345000 11.310000 ;
        RECT 11.145000 11.540000 11.345000 11.740000 ;
        RECT 11.145000 11.970000 11.345000 12.170000 ;
        RECT 11.145000 12.400000 11.345000 12.600000 ;
        RECT 11.145000 12.830000 11.345000 13.030000 ;
        RECT 11.145000 13.260000 11.345000 13.460000 ;
        RECT 11.550000  8.960000 11.750000  9.160000 ;
        RECT 11.550000  9.390000 11.750000  9.590000 ;
        RECT 11.550000  9.820000 11.750000 10.020000 ;
        RECT 11.550000 10.250000 11.750000 10.450000 ;
        RECT 11.550000 10.680000 11.750000 10.880000 ;
        RECT 11.550000 11.110000 11.750000 11.310000 ;
        RECT 11.550000 11.540000 11.750000 11.740000 ;
        RECT 11.550000 11.970000 11.750000 12.170000 ;
        RECT 11.550000 12.400000 11.750000 12.600000 ;
        RECT 11.550000 12.830000 11.750000 13.030000 ;
        RECT 11.550000 13.260000 11.750000 13.460000 ;
        RECT 11.955000  8.960000 12.155000  9.160000 ;
        RECT 11.955000  9.390000 12.155000  9.590000 ;
        RECT 11.955000  9.820000 12.155000 10.020000 ;
        RECT 11.955000 10.250000 12.155000 10.450000 ;
        RECT 11.955000 10.680000 12.155000 10.880000 ;
        RECT 11.955000 11.110000 12.155000 11.310000 ;
        RECT 11.955000 11.540000 12.155000 11.740000 ;
        RECT 11.955000 11.970000 12.155000 12.170000 ;
        RECT 11.955000 12.400000 12.155000 12.600000 ;
        RECT 11.955000 12.830000 12.155000 13.030000 ;
        RECT 11.955000 13.260000 12.155000 13.460000 ;
        RECT 12.360000  8.960000 12.560000  9.160000 ;
        RECT 12.360000  9.390000 12.560000  9.590000 ;
        RECT 12.360000  9.820000 12.560000 10.020000 ;
        RECT 12.360000 10.250000 12.560000 10.450000 ;
        RECT 12.360000 10.680000 12.560000 10.880000 ;
        RECT 12.360000 11.110000 12.560000 11.310000 ;
        RECT 12.360000 11.540000 12.560000 11.740000 ;
        RECT 12.360000 11.970000 12.560000 12.170000 ;
        RECT 12.360000 12.400000 12.560000 12.600000 ;
        RECT 12.360000 12.830000 12.560000 13.030000 ;
        RECT 12.360000 13.260000 12.560000 13.460000 ;
        RECT 12.765000  8.960000 12.965000  9.160000 ;
        RECT 12.765000  9.390000 12.965000  9.590000 ;
        RECT 12.765000  9.820000 12.965000 10.020000 ;
        RECT 12.765000 10.250000 12.965000 10.450000 ;
        RECT 12.765000 10.680000 12.965000 10.880000 ;
        RECT 12.765000 11.110000 12.965000 11.310000 ;
        RECT 12.765000 11.540000 12.965000 11.740000 ;
        RECT 12.765000 11.970000 12.965000 12.170000 ;
        RECT 12.765000 12.400000 12.965000 12.600000 ;
        RECT 12.765000 12.830000 12.965000 13.030000 ;
        RECT 12.765000 13.260000 12.965000 13.460000 ;
        RECT 13.170000  8.960000 13.370000  9.160000 ;
        RECT 13.170000  9.390000 13.370000  9.590000 ;
        RECT 13.170000  9.820000 13.370000 10.020000 ;
        RECT 13.170000 10.250000 13.370000 10.450000 ;
        RECT 13.170000 10.680000 13.370000 10.880000 ;
        RECT 13.170000 11.110000 13.370000 11.310000 ;
        RECT 13.170000 11.540000 13.370000 11.740000 ;
        RECT 13.170000 11.970000 13.370000 12.170000 ;
        RECT 13.170000 12.400000 13.370000 12.600000 ;
        RECT 13.170000 12.830000 13.370000 13.030000 ;
        RECT 13.170000 13.260000 13.370000 13.460000 ;
        RECT 13.575000  8.960000 13.775000  9.160000 ;
        RECT 13.575000  9.390000 13.775000  9.590000 ;
        RECT 13.575000  9.820000 13.775000 10.020000 ;
        RECT 13.575000 10.250000 13.775000 10.450000 ;
        RECT 13.575000 10.680000 13.775000 10.880000 ;
        RECT 13.575000 11.110000 13.775000 11.310000 ;
        RECT 13.575000 11.540000 13.775000 11.740000 ;
        RECT 13.575000 11.970000 13.775000 12.170000 ;
        RECT 13.575000 12.400000 13.775000 12.600000 ;
        RECT 13.575000 12.830000 13.775000 13.030000 ;
        RECT 13.575000 13.260000 13.775000 13.460000 ;
        RECT 13.980000  8.960000 14.180000  9.160000 ;
        RECT 13.980000  9.390000 14.180000  9.590000 ;
        RECT 13.980000  9.820000 14.180000 10.020000 ;
        RECT 13.980000 10.250000 14.180000 10.450000 ;
        RECT 13.980000 10.680000 14.180000 10.880000 ;
        RECT 13.980000 11.110000 14.180000 11.310000 ;
        RECT 13.980000 11.540000 14.180000 11.740000 ;
        RECT 13.980000 11.970000 14.180000 12.170000 ;
        RECT 13.980000 12.400000 14.180000 12.600000 ;
        RECT 13.980000 12.830000 14.180000 13.030000 ;
        RECT 13.980000 13.260000 14.180000 13.460000 ;
        RECT 14.385000  8.960000 14.585000  9.160000 ;
        RECT 14.385000  9.390000 14.585000  9.590000 ;
        RECT 14.385000  9.820000 14.585000 10.020000 ;
        RECT 14.385000 10.250000 14.585000 10.450000 ;
        RECT 14.385000 10.680000 14.585000 10.880000 ;
        RECT 14.385000 11.110000 14.585000 11.310000 ;
        RECT 14.385000 11.540000 14.585000 11.740000 ;
        RECT 14.385000 11.970000 14.585000 12.170000 ;
        RECT 14.385000 12.400000 14.585000 12.600000 ;
        RECT 14.385000 12.830000 14.585000 13.030000 ;
        RECT 14.385000 13.260000 14.585000 13.460000 ;
        RECT 14.790000  8.960000 14.990000  9.160000 ;
        RECT 14.790000  9.390000 14.990000  9.590000 ;
        RECT 14.790000  9.820000 14.990000 10.020000 ;
        RECT 14.790000 10.250000 14.990000 10.450000 ;
        RECT 14.790000 10.680000 14.990000 10.880000 ;
        RECT 14.790000 11.110000 14.990000 11.310000 ;
        RECT 14.790000 11.540000 14.990000 11.740000 ;
        RECT 14.790000 11.970000 14.990000 12.170000 ;
        RECT 14.790000 12.400000 14.990000 12.600000 ;
        RECT 14.790000 12.830000 14.990000 13.030000 ;
        RECT 14.790000 13.260000 14.990000 13.460000 ;
        RECT 15.195000  8.960000 15.395000  9.160000 ;
        RECT 15.195000  9.390000 15.395000  9.590000 ;
        RECT 15.195000  9.820000 15.395000 10.020000 ;
        RECT 15.195000 10.250000 15.395000 10.450000 ;
        RECT 15.195000 10.680000 15.395000 10.880000 ;
        RECT 15.195000 11.110000 15.395000 11.310000 ;
        RECT 15.195000 11.540000 15.395000 11.740000 ;
        RECT 15.195000 11.970000 15.395000 12.170000 ;
        RECT 15.195000 12.400000 15.395000 12.600000 ;
        RECT 15.195000 12.830000 15.395000 13.030000 ;
        RECT 15.195000 13.260000 15.395000 13.460000 ;
        RECT 15.600000  8.960000 15.800000  9.160000 ;
        RECT 15.600000  9.390000 15.800000  9.590000 ;
        RECT 15.600000  9.820000 15.800000 10.020000 ;
        RECT 15.600000 10.250000 15.800000 10.450000 ;
        RECT 15.600000 10.680000 15.800000 10.880000 ;
        RECT 15.600000 11.110000 15.800000 11.310000 ;
        RECT 15.600000 11.540000 15.800000 11.740000 ;
        RECT 15.600000 11.970000 15.800000 12.170000 ;
        RECT 15.600000 12.400000 15.800000 12.600000 ;
        RECT 15.600000 12.830000 15.800000 13.030000 ;
        RECT 15.600000 13.260000 15.800000 13.460000 ;
        RECT 16.005000  8.960000 16.205000  9.160000 ;
        RECT 16.005000  9.390000 16.205000  9.590000 ;
        RECT 16.005000  9.820000 16.205000 10.020000 ;
        RECT 16.005000 10.250000 16.205000 10.450000 ;
        RECT 16.005000 10.680000 16.205000 10.880000 ;
        RECT 16.005000 11.110000 16.205000 11.310000 ;
        RECT 16.005000 11.540000 16.205000 11.740000 ;
        RECT 16.005000 11.970000 16.205000 12.170000 ;
        RECT 16.005000 12.400000 16.205000 12.600000 ;
        RECT 16.005000 12.830000 16.205000 13.030000 ;
        RECT 16.005000 13.260000 16.205000 13.460000 ;
        RECT 16.410000  8.960000 16.610000  9.160000 ;
        RECT 16.410000  9.390000 16.610000  9.590000 ;
        RECT 16.410000  9.820000 16.610000 10.020000 ;
        RECT 16.410000 10.250000 16.610000 10.450000 ;
        RECT 16.410000 10.680000 16.610000 10.880000 ;
        RECT 16.410000 11.110000 16.610000 11.310000 ;
        RECT 16.410000 11.540000 16.610000 11.740000 ;
        RECT 16.410000 11.970000 16.610000 12.170000 ;
        RECT 16.410000 12.400000 16.610000 12.600000 ;
        RECT 16.410000 12.830000 16.610000 13.030000 ;
        RECT 16.410000 13.260000 16.610000 13.460000 ;
        RECT 16.815000  8.960000 17.015000  9.160000 ;
        RECT 16.815000  9.390000 17.015000  9.590000 ;
        RECT 16.815000  9.820000 17.015000 10.020000 ;
        RECT 16.815000 10.250000 17.015000 10.450000 ;
        RECT 16.815000 10.680000 17.015000 10.880000 ;
        RECT 16.815000 11.110000 17.015000 11.310000 ;
        RECT 16.815000 11.540000 17.015000 11.740000 ;
        RECT 16.815000 11.970000 17.015000 12.170000 ;
        RECT 16.815000 12.400000 17.015000 12.600000 ;
        RECT 16.815000 12.830000 17.015000 13.030000 ;
        RECT 16.815000 13.260000 17.015000 13.460000 ;
        RECT 17.220000  8.960000 17.420000  9.160000 ;
        RECT 17.220000  9.390000 17.420000  9.590000 ;
        RECT 17.220000  9.820000 17.420000 10.020000 ;
        RECT 17.220000 10.250000 17.420000 10.450000 ;
        RECT 17.220000 10.680000 17.420000 10.880000 ;
        RECT 17.220000 11.110000 17.420000 11.310000 ;
        RECT 17.220000 11.540000 17.420000 11.740000 ;
        RECT 17.220000 11.970000 17.420000 12.170000 ;
        RECT 17.220000 12.400000 17.420000 12.600000 ;
        RECT 17.220000 12.830000 17.420000 13.030000 ;
        RECT 17.220000 13.260000 17.420000 13.460000 ;
        RECT 17.625000  8.960000 17.825000  9.160000 ;
        RECT 17.625000  9.390000 17.825000  9.590000 ;
        RECT 17.625000  9.820000 17.825000 10.020000 ;
        RECT 17.625000 10.250000 17.825000 10.450000 ;
        RECT 17.625000 10.680000 17.825000 10.880000 ;
        RECT 17.625000 11.110000 17.825000 11.310000 ;
        RECT 17.625000 11.540000 17.825000 11.740000 ;
        RECT 17.625000 11.970000 17.825000 12.170000 ;
        RECT 17.625000 12.400000 17.825000 12.600000 ;
        RECT 17.625000 12.830000 17.825000 13.030000 ;
        RECT 17.625000 13.260000 17.825000 13.460000 ;
        RECT 18.030000  8.960000 18.230000  9.160000 ;
        RECT 18.030000  9.390000 18.230000  9.590000 ;
        RECT 18.030000  9.820000 18.230000 10.020000 ;
        RECT 18.030000 10.250000 18.230000 10.450000 ;
        RECT 18.030000 10.680000 18.230000 10.880000 ;
        RECT 18.030000 11.110000 18.230000 11.310000 ;
        RECT 18.030000 11.540000 18.230000 11.740000 ;
        RECT 18.030000 11.970000 18.230000 12.170000 ;
        RECT 18.030000 12.400000 18.230000 12.600000 ;
        RECT 18.030000 12.830000 18.230000 13.030000 ;
        RECT 18.030000 13.260000 18.230000 13.460000 ;
        RECT 18.435000  8.960000 18.635000  9.160000 ;
        RECT 18.435000  9.390000 18.635000  9.590000 ;
        RECT 18.435000  9.820000 18.635000 10.020000 ;
        RECT 18.435000 10.250000 18.635000 10.450000 ;
        RECT 18.435000 10.680000 18.635000 10.880000 ;
        RECT 18.435000 11.110000 18.635000 11.310000 ;
        RECT 18.435000 11.540000 18.635000 11.740000 ;
        RECT 18.435000 11.970000 18.635000 12.170000 ;
        RECT 18.435000 12.400000 18.635000 12.600000 ;
        RECT 18.435000 12.830000 18.635000 13.030000 ;
        RECT 18.435000 13.260000 18.635000 13.460000 ;
        RECT 18.840000  8.960000 19.040000  9.160000 ;
        RECT 18.840000  9.390000 19.040000  9.590000 ;
        RECT 18.840000  9.820000 19.040000 10.020000 ;
        RECT 18.840000 10.250000 19.040000 10.450000 ;
        RECT 18.840000 10.680000 19.040000 10.880000 ;
        RECT 18.840000 11.110000 19.040000 11.310000 ;
        RECT 18.840000 11.540000 19.040000 11.740000 ;
        RECT 18.840000 11.970000 19.040000 12.170000 ;
        RECT 18.840000 12.400000 19.040000 12.600000 ;
        RECT 18.840000 12.830000 19.040000 13.030000 ;
        RECT 18.840000 13.260000 19.040000 13.460000 ;
        RECT 19.245000  8.960000 19.445000  9.160000 ;
        RECT 19.245000  9.390000 19.445000  9.590000 ;
        RECT 19.245000  9.820000 19.445000 10.020000 ;
        RECT 19.245000 10.250000 19.445000 10.450000 ;
        RECT 19.245000 10.680000 19.445000 10.880000 ;
        RECT 19.245000 11.110000 19.445000 11.310000 ;
        RECT 19.245000 11.540000 19.445000 11.740000 ;
        RECT 19.245000 11.970000 19.445000 12.170000 ;
        RECT 19.245000 12.400000 19.445000 12.600000 ;
        RECT 19.245000 12.830000 19.445000 13.030000 ;
        RECT 19.245000 13.260000 19.445000 13.460000 ;
        RECT 19.650000  8.960000 19.850000  9.160000 ;
        RECT 19.650000  9.390000 19.850000  9.590000 ;
        RECT 19.650000  9.820000 19.850000 10.020000 ;
        RECT 19.650000 10.250000 19.850000 10.450000 ;
        RECT 19.650000 10.680000 19.850000 10.880000 ;
        RECT 19.650000 11.110000 19.850000 11.310000 ;
        RECT 19.650000 11.540000 19.850000 11.740000 ;
        RECT 19.650000 11.970000 19.850000 12.170000 ;
        RECT 19.650000 12.400000 19.850000 12.600000 ;
        RECT 19.650000 12.830000 19.850000 13.030000 ;
        RECT 19.650000 13.260000 19.850000 13.460000 ;
        RECT 20.055000  8.960000 20.255000  9.160000 ;
        RECT 20.055000  9.390000 20.255000  9.590000 ;
        RECT 20.055000  9.820000 20.255000 10.020000 ;
        RECT 20.055000 10.250000 20.255000 10.450000 ;
        RECT 20.055000 10.680000 20.255000 10.880000 ;
        RECT 20.055000 11.110000 20.255000 11.310000 ;
        RECT 20.055000 11.540000 20.255000 11.740000 ;
        RECT 20.055000 11.970000 20.255000 12.170000 ;
        RECT 20.055000 12.400000 20.255000 12.600000 ;
        RECT 20.055000 12.830000 20.255000 13.030000 ;
        RECT 20.055000 13.260000 20.255000 13.460000 ;
        RECT 20.460000  8.960000 20.660000  9.160000 ;
        RECT 20.460000  9.390000 20.660000  9.590000 ;
        RECT 20.460000  9.820000 20.660000 10.020000 ;
        RECT 20.460000 10.250000 20.660000 10.450000 ;
        RECT 20.460000 10.680000 20.660000 10.880000 ;
        RECT 20.460000 11.110000 20.660000 11.310000 ;
        RECT 20.460000 11.540000 20.660000 11.740000 ;
        RECT 20.460000 11.970000 20.660000 12.170000 ;
        RECT 20.460000 12.400000 20.660000 12.600000 ;
        RECT 20.460000 12.830000 20.660000 13.030000 ;
        RECT 20.460000 13.260000 20.660000 13.460000 ;
        RECT 20.865000  8.960000 21.065000  9.160000 ;
        RECT 20.865000  9.390000 21.065000  9.590000 ;
        RECT 20.865000  9.820000 21.065000 10.020000 ;
        RECT 20.865000 10.250000 21.065000 10.450000 ;
        RECT 20.865000 10.680000 21.065000 10.880000 ;
        RECT 20.865000 11.110000 21.065000 11.310000 ;
        RECT 20.865000 11.540000 21.065000 11.740000 ;
        RECT 20.865000 11.970000 21.065000 12.170000 ;
        RECT 20.865000 12.400000 21.065000 12.600000 ;
        RECT 20.865000 12.830000 21.065000 13.030000 ;
        RECT 20.865000 13.260000 21.065000 13.460000 ;
        RECT 21.270000  8.960000 21.470000  9.160000 ;
        RECT 21.270000  9.390000 21.470000  9.590000 ;
        RECT 21.270000  9.820000 21.470000 10.020000 ;
        RECT 21.270000 10.250000 21.470000 10.450000 ;
        RECT 21.270000 10.680000 21.470000 10.880000 ;
        RECT 21.270000 11.110000 21.470000 11.310000 ;
        RECT 21.270000 11.540000 21.470000 11.740000 ;
        RECT 21.270000 11.970000 21.470000 12.170000 ;
        RECT 21.270000 12.400000 21.470000 12.600000 ;
        RECT 21.270000 12.830000 21.470000 13.030000 ;
        RECT 21.270000 13.260000 21.470000 13.460000 ;
        RECT 21.675000  8.960000 21.875000  9.160000 ;
        RECT 21.675000  9.390000 21.875000  9.590000 ;
        RECT 21.675000  9.820000 21.875000 10.020000 ;
        RECT 21.675000 10.250000 21.875000 10.450000 ;
        RECT 21.675000 10.680000 21.875000 10.880000 ;
        RECT 21.675000 11.110000 21.875000 11.310000 ;
        RECT 21.675000 11.540000 21.875000 11.740000 ;
        RECT 21.675000 11.970000 21.875000 12.170000 ;
        RECT 21.675000 12.400000 21.875000 12.600000 ;
        RECT 21.675000 12.830000 21.875000 13.030000 ;
        RECT 21.675000 13.260000 21.875000 13.460000 ;
        RECT 22.080000  8.960000 22.280000  9.160000 ;
        RECT 22.080000  9.390000 22.280000  9.590000 ;
        RECT 22.080000  9.820000 22.280000 10.020000 ;
        RECT 22.080000 10.250000 22.280000 10.450000 ;
        RECT 22.080000 10.680000 22.280000 10.880000 ;
        RECT 22.080000 11.110000 22.280000 11.310000 ;
        RECT 22.080000 11.540000 22.280000 11.740000 ;
        RECT 22.080000 11.970000 22.280000 12.170000 ;
        RECT 22.080000 12.400000 22.280000 12.600000 ;
        RECT 22.080000 12.830000 22.280000 13.030000 ;
        RECT 22.080000 13.260000 22.280000 13.460000 ;
        RECT 22.485000  8.960000 22.685000  9.160000 ;
        RECT 22.485000  9.390000 22.685000  9.590000 ;
        RECT 22.485000  9.820000 22.685000 10.020000 ;
        RECT 22.485000 10.250000 22.685000 10.450000 ;
        RECT 22.485000 10.680000 22.685000 10.880000 ;
        RECT 22.485000 11.110000 22.685000 11.310000 ;
        RECT 22.485000 11.540000 22.685000 11.740000 ;
        RECT 22.485000 11.970000 22.685000 12.170000 ;
        RECT 22.485000 12.400000 22.685000 12.600000 ;
        RECT 22.485000 12.830000 22.685000 13.030000 ;
        RECT 22.485000 13.260000 22.685000 13.460000 ;
        RECT 22.890000  8.960000 23.090000  9.160000 ;
        RECT 22.890000  9.390000 23.090000  9.590000 ;
        RECT 22.890000  9.820000 23.090000 10.020000 ;
        RECT 22.890000 10.250000 23.090000 10.450000 ;
        RECT 22.890000 10.680000 23.090000 10.880000 ;
        RECT 22.890000 11.110000 23.090000 11.310000 ;
        RECT 22.890000 11.540000 23.090000 11.740000 ;
        RECT 22.890000 11.970000 23.090000 12.170000 ;
        RECT 22.890000 12.400000 23.090000 12.600000 ;
        RECT 22.890000 12.830000 23.090000 13.030000 ;
        RECT 22.890000 13.260000 23.090000 13.460000 ;
        RECT 23.295000  8.960000 23.495000  9.160000 ;
        RECT 23.295000  9.390000 23.495000  9.590000 ;
        RECT 23.295000  9.820000 23.495000 10.020000 ;
        RECT 23.295000 10.250000 23.495000 10.450000 ;
        RECT 23.295000 10.680000 23.495000 10.880000 ;
        RECT 23.295000 11.110000 23.495000 11.310000 ;
        RECT 23.295000 11.540000 23.495000 11.740000 ;
        RECT 23.295000 11.970000 23.495000 12.170000 ;
        RECT 23.295000 12.400000 23.495000 12.600000 ;
        RECT 23.295000 12.830000 23.495000 13.030000 ;
        RECT 23.295000 13.260000 23.495000 13.460000 ;
        RECT 23.700000  8.960000 23.900000  9.160000 ;
        RECT 23.700000  9.390000 23.900000  9.590000 ;
        RECT 23.700000  9.820000 23.900000 10.020000 ;
        RECT 23.700000 10.250000 23.900000 10.450000 ;
        RECT 23.700000 10.680000 23.900000 10.880000 ;
        RECT 23.700000 11.110000 23.900000 11.310000 ;
        RECT 23.700000 11.540000 23.900000 11.740000 ;
        RECT 23.700000 11.970000 23.900000 12.170000 ;
        RECT 23.700000 12.400000 23.900000 12.600000 ;
        RECT 23.700000 12.830000 23.900000 13.030000 ;
        RECT 23.700000 13.260000 23.900000 13.460000 ;
        RECT 24.105000  8.960000 24.305000  9.160000 ;
        RECT 24.105000  9.390000 24.305000  9.590000 ;
        RECT 24.105000  9.820000 24.305000 10.020000 ;
        RECT 24.105000 10.250000 24.305000 10.450000 ;
        RECT 24.105000 10.680000 24.305000 10.880000 ;
        RECT 24.105000 11.110000 24.305000 11.310000 ;
        RECT 24.105000 11.540000 24.305000 11.740000 ;
        RECT 24.105000 11.970000 24.305000 12.170000 ;
        RECT 24.105000 12.400000 24.305000 12.600000 ;
        RECT 24.105000 12.830000 24.305000 13.030000 ;
        RECT 24.105000 13.260000 24.305000 13.460000 ;
        RECT 50.480000  8.960000 50.680000  9.160000 ;
        RECT 50.480000  9.390000 50.680000  9.590000 ;
        RECT 50.480000  9.820000 50.680000 10.020000 ;
        RECT 50.480000 10.250000 50.680000 10.450000 ;
        RECT 50.480000 10.680000 50.680000 10.880000 ;
        RECT 50.480000 11.110000 50.680000 11.310000 ;
        RECT 50.480000 11.540000 50.680000 11.740000 ;
        RECT 50.480000 11.970000 50.680000 12.170000 ;
        RECT 50.480000 12.400000 50.680000 12.600000 ;
        RECT 50.480000 12.830000 50.680000 13.030000 ;
        RECT 50.480000 13.260000 50.680000 13.460000 ;
        RECT 50.890000  8.960000 51.090000  9.160000 ;
        RECT 50.890000  9.390000 51.090000  9.590000 ;
        RECT 50.890000  9.820000 51.090000 10.020000 ;
        RECT 50.890000 10.250000 51.090000 10.450000 ;
        RECT 50.890000 10.680000 51.090000 10.880000 ;
        RECT 50.890000 11.110000 51.090000 11.310000 ;
        RECT 50.890000 11.540000 51.090000 11.740000 ;
        RECT 50.890000 11.970000 51.090000 12.170000 ;
        RECT 50.890000 12.400000 51.090000 12.600000 ;
        RECT 50.890000 12.830000 51.090000 13.030000 ;
        RECT 50.890000 13.260000 51.090000 13.460000 ;
        RECT 51.300000  8.960000 51.500000  9.160000 ;
        RECT 51.300000  9.390000 51.500000  9.590000 ;
        RECT 51.300000  9.820000 51.500000 10.020000 ;
        RECT 51.300000 10.250000 51.500000 10.450000 ;
        RECT 51.300000 10.680000 51.500000 10.880000 ;
        RECT 51.300000 11.110000 51.500000 11.310000 ;
        RECT 51.300000 11.540000 51.500000 11.740000 ;
        RECT 51.300000 11.970000 51.500000 12.170000 ;
        RECT 51.300000 12.400000 51.500000 12.600000 ;
        RECT 51.300000 12.830000 51.500000 13.030000 ;
        RECT 51.300000 13.260000 51.500000 13.460000 ;
        RECT 51.710000  8.960000 51.910000  9.160000 ;
        RECT 51.710000  9.390000 51.910000  9.590000 ;
        RECT 51.710000  9.820000 51.910000 10.020000 ;
        RECT 51.710000 10.250000 51.910000 10.450000 ;
        RECT 51.710000 10.680000 51.910000 10.880000 ;
        RECT 51.710000 11.110000 51.910000 11.310000 ;
        RECT 51.710000 11.540000 51.910000 11.740000 ;
        RECT 51.710000 11.970000 51.910000 12.170000 ;
        RECT 51.710000 12.400000 51.910000 12.600000 ;
        RECT 51.710000 12.830000 51.910000 13.030000 ;
        RECT 51.710000 13.260000 51.910000 13.460000 ;
        RECT 52.120000  8.960000 52.320000  9.160000 ;
        RECT 52.120000  9.390000 52.320000  9.590000 ;
        RECT 52.120000  9.820000 52.320000 10.020000 ;
        RECT 52.120000 10.250000 52.320000 10.450000 ;
        RECT 52.120000 10.680000 52.320000 10.880000 ;
        RECT 52.120000 11.110000 52.320000 11.310000 ;
        RECT 52.120000 11.540000 52.320000 11.740000 ;
        RECT 52.120000 11.970000 52.320000 12.170000 ;
        RECT 52.120000 12.400000 52.320000 12.600000 ;
        RECT 52.120000 12.830000 52.320000 13.030000 ;
        RECT 52.120000 13.260000 52.320000 13.460000 ;
        RECT 52.530000  8.960000 52.730000  9.160000 ;
        RECT 52.530000  9.390000 52.730000  9.590000 ;
        RECT 52.530000  9.820000 52.730000 10.020000 ;
        RECT 52.530000 10.250000 52.730000 10.450000 ;
        RECT 52.530000 10.680000 52.730000 10.880000 ;
        RECT 52.530000 11.110000 52.730000 11.310000 ;
        RECT 52.530000 11.540000 52.730000 11.740000 ;
        RECT 52.530000 11.970000 52.730000 12.170000 ;
        RECT 52.530000 12.400000 52.730000 12.600000 ;
        RECT 52.530000 12.830000 52.730000 13.030000 ;
        RECT 52.530000 13.260000 52.730000 13.460000 ;
        RECT 52.940000  8.960000 53.140000  9.160000 ;
        RECT 52.940000  9.390000 53.140000  9.590000 ;
        RECT 52.940000  9.820000 53.140000 10.020000 ;
        RECT 52.940000 10.250000 53.140000 10.450000 ;
        RECT 52.940000 10.680000 53.140000 10.880000 ;
        RECT 52.940000 11.110000 53.140000 11.310000 ;
        RECT 52.940000 11.540000 53.140000 11.740000 ;
        RECT 52.940000 11.970000 53.140000 12.170000 ;
        RECT 52.940000 12.400000 53.140000 12.600000 ;
        RECT 52.940000 12.830000 53.140000 13.030000 ;
        RECT 52.940000 13.260000 53.140000 13.460000 ;
        RECT 53.345000  8.960000 53.545000  9.160000 ;
        RECT 53.345000  9.390000 53.545000  9.590000 ;
        RECT 53.345000  9.820000 53.545000 10.020000 ;
        RECT 53.345000 10.250000 53.545000 10.450000 ;
        RECT 53.345000 10.680000 53.545000 10.880000 ;
        RECT 53.345000 11.110000 53.545000 11.310000 ;
        RECT 53.345000 11.540000 53.545000 11.740000 ;
        RECT 53.345000 11.970000 53.545000 12.170000 ;
        RECT 53.345000 12.400000 53.545000 12.600000 ;
        RECT 53.345000 12.830000 53.545000 13.030000 ;
        RECT 53.345000 13.260000 53.545000 13.460000 ;
        RECT 53.750000  8.960000 53.950000  9.160000 ;
        RECT 53.750000  9.390000 53.950000  9.590000 ;
        RECT 53.750000  9.820000 53.950000 10.020000 ;
        RECT 53.750000 10.250000 53.950000 10.450000 ;
        RECT 53.750000 10.680000 53.950000 10.880000 ;
        RECT 53.750000 11.110000 53.950000 11.310000 ;
        RECT 53.750000 11.540000 53.950000 11.740000 ;
        RECT 53.750000 11.970000 53.950000 12.170000 ;
        RECT 53.750000 12.400000 53.950000 12.600000 ;
        RECT 53.750000 12.830000 53.950000 13.030000 ;
        RECT 53.750000 13.260000 53.950000 13.460000 ;
        RECT 54.155000  8.960000 54.355000  9.160000 ;
        RECT 54.155000  9.390000 54.355000  9.590000 ;
        RECT 54.155000  9.820000 54.355000 10.020000 ;
        RECT 54.155000 10.250000 54.355000 10.450000 ;
        RECT 54.155000 10.680000 54.355000 10.880000 ;
        RECT 54.155000 11.110000 54.355000 11.310000 ;
        RECT 54.155000 11.540000 54.355000 11.740000 ;
        RECT 54.155000 11.970000 54.355000 12.170000 ;
        RECT 54.155000 12.400000 54.355000 12.600000 ;
        RECT 54.155000 12.830000 54.355000 13.030000 ;
        RECT 54.155000 13.260000 54.355000 13.460000 ;
        RECT 54.560000  8.960000 54.760000  9.160000 ;
        RECT 54.560000  9.390000 54.760000  9.590000 ;
        RECT 54.560000  9.820000 54.760000 10.020000 ;
        RECT 54.560000 10.250000 54.760000 10.450000 ;
        RECT 54.560000 10.680000 54.760000 10.880000 ;
        RECT 54.560000 11.110000 54.760000 11.310000 ;
        RECT 54.560000 11.540000 54.760000 11.740000 ;
        RECT 54.560000 11.970000 54.760000 12.170000 ;
        RECT 54.560000 12.400000 54.760000 12.600000 ;
        RECT 54.560000 12.830000 54.760000 13.030000 ;
        RECT 54.560000 13.260000 54.760000 13.460000 ;
        RECT 54.965000  8.960000 55.165000  9.160000 ;
        RECT 54.965000  9.390000 55.165000  9.590000 ;
        RECT 54.965000  9.820000 55.165000 10.020000 ;
        RECT 54.965000 10.250000 55.165000 10.450000 ;
        RECT 54.965000 10.680000 55.165000 10.880000 ;
        RECT 54.965000 11.110000 55.165000 11.310000 ;
        RECT 54.965000 11.540000 55.165000 11.740000 ;
        RECT 54.965000 11.970000 55.165000 12.170000 ;
        RECT 54.965000 12.400000 55.165000 12.600000 ;
        RECT 54.965000 12.830000 55.165000 13.030000 ;
        RECT 54.965000 13.260000 55.165000 13.460000 ;
        RECT 55.370000  8.960000 55.570000  9.160000 ;
        RECT 55.370000  9.390000 55.570000  9.590000 ;
        RECT 55.370000  9.820000 55.570000 10.020000 ;
        RECT 55.370000 10.250000 55.570000 10.450000 ;
        RECT 55.370000 10.680000 55.570000 10.880000 ;
        RECT 55.370000 11.110000 55.570000 11.310000 ;
        RECT 55.370000 11.540000 55.570000 11.740000 ;
        RECT 55.370000 11.970000 55.570000 12.170000 ;
        RECT 55.370000 12.400000 55.570000 12.600000 ;
        RECT 55.370000 12.830000 55.570000 13.030000 ;
        RECT 55.370000 13.260000 55.570000 13.460000 ;
        RECT 55.775000  8.960000 55.975000  9.160000 ;
        RECT 55.775000  9.390000 55.975000  9.590000 ;
        RECT 55.775000  9.820000 55.975000 10.020000 ;
        RECT 55.775000 10.250000 55.975000 10.450000 ;
        RECT 55.775000 10.680000 55.975000 10.880000 ;
        RECT 55.775000 11.110000 55.975000 11.310000 ;
        RECT 55.775000 11.540000 55.975000 11.740000 ;
        RECT 55.775000 11.970000 55.975000 12.170000 ;
        RECT 55.775000 12.400000 55.975000 12.600000 ;
        RECT 55.775000 12.830000 55.975000 13.030000 ;
        RECT 55.775000 13.260000 55.975000 13.460000 ;
        RECT 56.180000  8.960000 56.380000  9.160000 ;
        RECT 56.180000  9.390000 56.380000  9.590000 ;
        RECT 56.180000  9.820000 56.380000 10.020000 ;
        RECT 56.180000 10.250000 56.380000 10.450000 ;
        RECT 56.180000 10.680000 56.380000 10.880000 ;
        RECT 56.180000 11.110000 56.380000 11.310000 ;
        RECT 56.180000 11.540000 56.380000 11.740000 ;
        RECT 56.180000 11.970000 56.380000 12.170000 ;
        RECT 56.180000 12.400000 56.380000 12.600000 ;
        RECT 56.180000 12.830000 56.380000 13.030000 ;
        RECT 56.180000 13.260000 56.380000 13.460000 ;
        RECT 56.585000  8.960000 56.785000  9.160000 ;
        RECT 56.585000  9.390000 56.785000  9.590000 ;
        RECT 56.585000  9.820000 56.785000 10.020000 ;
        RECT 56.585000 10.250000 56.785000 10.450000 ;
        RECT 56.585000 10.680000 56.785000 10.880000 ;
        RECT 56.585000 11.110000 56.785000 11.310000 ;
        RECT 56.585000 11.540000 56.785000 11.740000 ;
        RECT 56.585000 11.970000 56.785000 12.170000 ;
        RECT 56.585000 12.400000 56.785000 12.600000 ;
        RECT 56.585000 12.830000 56.785000 13.030000 ;
        RECT 56.585000 13.260000 56.785000 13.460000 ;
        RECT 56.990000  8.960000 57.190000  9.160000 ;
        RECT 56.990000  9.390000 57.190000  9.590000 ;
        RECT 56.990000  9.820000 57.190000 10.020000 ;
        RECT 56.990000 10.250000 57.190000 10.450000 ;
        RECT 56.990000 10.680000 57.190000 10.880000 ;
        RECT 56.990000 11.110000 57.190000 11.310000 ;
        RECT 56.990000 11.540000 57.190000 11.740000 ;
        RECT 56.990000 11.970000 57.190000 12.170000 ;
        RECT 56.990000 12.400000 57.190000 12.600000 ;
        RECT 56.990000 12.830000 57.190000 13.030000 ;
        RECT 56.990000 13.260000 57.190000 13.460000 ;
        RECT 57.395000  8.960000 57.595000  9.160000 ;
        RECT 57.395000  9.390000 57.595000  9.590000 ;
        RECT 57.395000  9.820000 57.595000 10.020000 ;
        RECT 57.395000 10.250000 57.595000 10.450000 ;
        RECT 57.395000 10.680000 57.595000 10.880000 ;
        RECT 57.395000 11.110000 57.595000 11.310000 ;
        RECT 57.395000 11.540000 57.595000 11.740000 ;
        RECT 57.395000 11.970000 57.595000 12.170000 ;
        RECT 57.395000 12.400000 57.595000 12.600000 ;
        RECT 57.395000 12.830000 57.595000 13.030000 ;
        RECT 57.395000 13.260000 57.595000 13.460000 ;
        RECT 57.800000  8.960000 58.000000  9.160000 ;
        RECT 57.800000  9.390000 58.000000  9.590000 ;
        RECT 57.800000  9.820000 58.000000 10.020000 ;
        RECT 57.800000 10.250000 58.000000 10.450000 ;
        RECT 57.800000 10.680000 58.000000 10.880000 ;
        RECT 57.800000 11.110000 58.000000 11.310000 ;
        RECT 57.800000 11.540000 58.000000 11.740000 ;
        RECT 57.800000 11.970000 58.000000 12.170000 ;
        RECT 57.800000 12.400000 58.000000 12.600000 ;
        RECT 57.800000 12.830000 58.000000 13.030000 ;
        RECT 57.800000 13.260000 58.000000 13.460000 ;
        RECT 58.205000  8.960000 58.405000  9.160000 ;
        RECT 58.205000  9.390000 58.405000  9.590000 ;
        RECT 58.205000  9.820000 58.405000 10.020000 ;
        RECT 58.205000 10.250000 58.405000 10.450000 ;
        RECT 58.205000 10.680000 58.405000 10.880000 ;
        RECT 58.205000 11.110000 58.405000 11.310000 ;
        RECT 58.205000 11.540000 58.405000 11.740000 ;
        RECT 58.205000 11.970000 58.405000 12.170000 ;
        RECT 58.205000 12.400000 58.405000 12.600000 ;
        RECT 58.205000 12.830000 58.405000 13.030000 ;
        RECT 58.205000 13.260000 58.405000 13.460000 ;
        RECT 58.610000  8.960000 58.810000  9.160000 ;
        RECT 58.610000  9.390000 58.810000  9.590000 ;
        RECT 58.610000  9.820000 58.810000 10.020000 ;
        RECT 58.610000 10.250000 58.810000 10.450000 ;
        RECT 58.610000 10.680000 58.810000 10.880000 ;
        RECT 58.610000 11.110000 58.810000 11.310000 ;
        RECT 58.610000 11.540000 58.810000 11.740000 ;
        RECT 58.610000 11.970000 58.810000 12.170000 ;
        RECT 58.610000 12.400000 58.810000 12.600000 ;
        RECT 58.610000 12.830000 58.810000 13.030000 ;
        RECT 58.610000 13.260000 58.810000 13.460000 ;
        RECT 59.015000  8.960000 59.215000  9.160000 ;
        RECT 59.015000  9.390000 59.215000  9.590000 ;
        RECT 59.015000  9.820000 59.215000 10.020000 ;
        RECT 59.015000 10.250000 59.215000 10.450000 ;
        RECT 59.015000 10.680000 59.215000 10.880000 ;
        RECT 59.015000 11.110000 59.215000 11.310000 ;
        RECT 59.015000 11.540000 59.215000 11.740000 ;
        RECT 59.015000 11.970000 59.215000 12.170000 ;
        RECT 59.015000 12.400000 59.215000 12.600000 ;
        RECT 59.015000 12.830000 59.215000 13.030000 ;
        RECT 59.015000 13.260000 59.215000 13.460000 ;
        RECT 59.420000  8.960000 59.620000  9.160000 ;
        RECT 59.420000  9.390000 59.620000  9.590000 ;
        RECT 59.420000  9.820000 59.620000 10.020000 ;
        RECT 59.420000 10.250000 59.620000 10.450000 ;
        RECT 59.420000 10.680000 59.620000 10.880000 ;
        RECT 59.420000 11.110000 59.620000 11.310000 ;
        RECT 59.420000 11.540000 59.620000 11.740000 ;
        RECT 59.420000 11.970000 59.620000 12.170000 ;
        RECT 59.420000 12.400000 59.620000 12.600000 ;
        RECT 59.420000 12.830000 59.620000 13.030000 ;
        RECT 59.420000 13.260000 59.620000 13.460000 ;
        RECT 59.825000  8.960000 60.025000  9.160000 ;
        RECT 59.825000  9.390000 60.025000  9.590000 ;
        RECT 59.825000  9.820000 60.025000 10.020000 ;
        RECT 59.825000 10.250000 60.025000 10.450000 ;
        RECT 59.825000 10.680000 60.025000 10.880000 ;
        RECT 59.825000 11.110000 60.025000 11.310000 ;
        RECT 59.825000 11.540000 60.025000 11.740000 ;
        RECT 59.825000 11.970000 60.025000 12.170000 ;
        RECT 59.825000 12.400000 60.025000 12.600000 ;
        RECT 59.825000 12.830000 60.025000 13.030000 ;
        RECT 59.825000 13.260000 60.025000 13.460000 ;
        RECT 60.230000  8.960000 60.430000  9.160000 ;
        RECT 60.230000  9.390000 60.430000  9.590000 ;
        RECT 60.230000  9.820000 60.430000 10.020000 ;
        RECT 60.230000 10.250000 60.430000 10.450000 ;
        RECT 60.230000 10.680000 60.430000 10.880000 ;
        RECT 60.230000 11.110000 60.430000 11.310000 ;
        RECT 60.230000 11.540000 60.430000 11.740000 ;
        RECT 60.230000 11.970000 60.430000 12.170000 ;
        RECT 60.230000 12.400000 60.430000 12.600000 ;
        RECT 60.230000 12.830000 60.430000 13.030000 ;
        RECT 60.230000 13.260000 60.430000 13.460000 ;
        RECT 60.635000  8.960000 60.835000  9.160000 ;
        RECT 60.635000  9.390000 60.835000  9.590000 ;
        RECT 60.635000  9.820000 60.835000 10.020000 ;
        RECT 60.635000 10.250000 60.835000 10.450000 ;
        RECT 60.635000 10.680000 60.835000 10.880000 ;
        RECT 60.635000 11.110000 60.835000 11.310000 ;
        RECT 60.635000 11.540000 60.835000 11.740000 ;
        RECT 60.635000 11.970000 60.835000 12.170000 ;
        RECT 60.635000 12.400000 60.835000 12.600000 ;
        RECT 60.635000 12.830000 60.835000 13.030000 ;
        RECT 60.635000 13.260000 60.835000 13.460000 ;
        RECT 61.040000  8.960000 61.240000  9.160000 ;
        RECT 61.040000  9.390000 61.240000  9.590000 ;
        RECT 61.040000  9.820000 61.240000 10.020000 ;
        RECT 61.040000 10.250000 61.240000 10.450000 ;
        RECT 61.040000 10.680000 61.240000 10.880000 ;
        RECT 61.040000 11.110000 61.240000 11.310000 ;
        RECT 61.040000 11.540000 61.240000 11.740000 ;
        RECT 61.040000 11.970000 61.240000 12.170000 ;
        RECT 61.040000 12.400000 61.240000 12.600000 ;
        RECT 61.040000 12.830000 61.240000 13.030000 ;
        RECT 61.040000 13.260000 61.240000 13.460000 ;
        RECT 61.445000  8.960000 61.645000  9.160000 ;
        RECT 61.445000  9.390000 61.645000  9.590000 ;
        RECT 61.445000  9.820000 61.645000 10.020000 ;
        RECT 61.445000 10.250000 61.645000 10.450000 ;
        RECT 61.445000 10.680000 61.645000 10.880000 ;
        RECT 61.445000 11.110000 61.645000 11.310000 ;
        RECT 61.445000 11.540000 61.645000 11.740000 ;
        RECT 61.445000 11.970000 61.645000 12.170000 ;
        RECT 61.445000 12.400000 61.645000 12.600000 ;
        RECT 61.445000 12.830000 61.645000 13.030000 ;
        RECT 61.445000 13.260000 61.645000 13.460000 ;
        RECT 61.850000  8.960000 62.050000  9.160000 ;
        RECT 61.850000  9.390000 62.050000  9.590000 ;
        RECT 61.850000  9.820000 62.050000 10.020000 ;
        RECT 61.850000 10.250000 62.050000 10.450000 ;
        RECT 61.850000 10.680000 62.050000 10.880000 ;
        RECT 61.850000 11.110000 62.050000 11.310000 ;
        RECT 61.850000 11.540000 62.050000 11.740000 ;
        RECT 61.850000 11.970000 62.050000 12.170000 ;
        RECT 61.850000 12.400000 62.050000 12.600000 ;
        RECT 61.850000 12.830000 62.050000 13.030000 ;
        RECT 61.850000 13.260000 62.050000 13.460000 ;
        RECT 62.255000  8.960000 62.455000  9.160000 ;
        RECT 62.255000  9.390000 62.455000  9.590000 ;
        RECT 62.255000  9.820000 62.455000 10.020000 ;
        RECT 62.255000 10.250000 62.455000 10.450000 ;
        RECT 62.255000 10.680000 62.455000 10.880000 ;
        RECT 62.255000 11.110000 62.455000 11.310000 ;
        RECT 62.255000 11.540000 62.455000 11.740000 ;
        RECT 62.255000 11.970000 62.455000 12.170000 ;
        RECT 62.255000 12.400000 62.455000 12.600000 ;
        RECT 62.255000 12.830000 62.455000 13.030000 ;
        RECT 62.255000 13.260000 62.455000 13.460000 ;
        RECT 62.660000  8.960000 62.860000  9.160000 ;
        RECT 62.660000  9.390000 62.860000  9.590000 ;
        RECT 62.660000  9.820000 62.860000 10.020000 ;
        RECT 62.660000 10.250000 62.860000 10.450000 ;
        RECT 62.660000 10.680000 62.860000 10.880000 ;
        RECT 62.660000 11.110000 62.860000 11.310000 ;
        RECT 62.660000 11.540000 62.860000 11.740000 ;
        RECT 62.660000 11.970000 62.860000 12.170000 ;
        RECT 62.660000 12.400000 62.860000 12.600000 ;
        RECT 62.660000 12.830000 62.860000 13.030000 ;
        RECT 62.660000 13.260000 62.860000 13.460000 ;
        RECT 63.065000  8.960000 63.265000  9.160000 ;
        RECT 63.065000  9.390000 63.265000  9.590000 ;
        RECT 63.065000  9.820000 63.265000 10.020000 ;
        RECT 63.065000 10.250000 63.265000 10.450000 ;
        RECT 63.065000 10.680000 63.265000 10.880000 ;
        RECT 63.065000 11.110000 63.265000 11.310000 ;
        RECT 63.065000 11.540000 63.265000 11.740000 ;
        RECT 63.065000 11.970000 63.265000 12.170000 ;
        RECT 63.065000 12.400000 63.265000 12.600000 ;
        RECT 63.065000 12.830000 63.265000 13.030000 ;
        RECT 63.065000 13.260000 63.265000 13.460000 ;
        RECT 63.470000  8.960000 63.670000  9.160000 ;
        RECT 63.470000  9.390000 63.670000  9.590000 ;
        RECT 63.470000  9.820000 63.670000 10.020000 ;
        RECT 63.470000 10.250000 63.670000 10.450000 ;
        RECT 63.470000 10.680000 63.670000 10.880000 ;
        RECT 63.470000 11.110000 63.670000 11.310000 ;
        RECT 63.470000 11.540000 63.670000 11.740000 ;
        RECT 63.470000 11.970000 63.670000 12.170000 ;
        RECT 63.470000 12.400000 63.670000 12.600000 ;
        RECT 63.470000 12.830000 63.670000 13.030000 ;
        RECT 63.470000 13.260000 63.670000 13.460000 ;
        RECT 63.875000  8.960000 64.075000  9.160000 ;
        RECT 63.875000  9.390000 64.075000  9.590000 ;
        RECT 63.875000  9.820000 64.075000 10.020000 ;
        RECT 63.875000 10.250000 64.075000 10.450000 ;
        RECT 63.875000 10.680000 64.075000 10.880000 ;
        RECT 63.875000 11.110000 64.075000 11.310000 ;
        RECT 63.875000 11.540000 64.075000 11.740000 ;
        RECT 63.875000 11.970000 64.075000 12.170000 ;
        RECT 63.875000 12.400000 64.075000 12.600000 ;
        RECT 63.875000 12.830000 64.075000 13.030000 ;
        RECT 63.875000 13.260000 64.075000 13.460000 ;
        RECT 64.280000  8.960000 64.480000  9.160000 ;
        RECT 64.280000  9.390000 64.480000  9.590000 ;
        RECT 64.280000  9.820000 64.480000 10.020000 ;
        RECT 64.280000 10.250000 64.480000 10.450000 ;
        RECT 64.280000 10.680000 64.480000 10.880000 ;
        RECT 64.280000 11.110000 64.480000 11.310000 ;
        RECT 64.280000 11.540000 64.480000 11.740000 ;
        RECT 64.280000 11.970000 64.480000 12.170000 ;
        RECT 64.280000 12.400000 64.480000 12.600000 ;
        RECT 64.280000 12.830000 64.480000 13.030000 ;
        RECT 64.280000 13.260000 64.480000 13.460000 ;
        RECT 64.685000  8.960000 64.885000  9.160000 ;
        RECT 64.685000  9.390000 64.885000  9.590000 ;
        RECT 64.685000  9.820000 64.885000 10.020000 ;
        RECT 64.685000 10.250000 64.885000 10.450000 ;
        RECT 64.685000 10.680000 64.885000 10.880000 ;
        RECT 64.685000 11.110000 64.885000 11.310000 ;
        RECT 64.685000 11.540000 64.885000 11.740000 ;
        RECT 64.685000 11.970000 64.885000 12.170000 ;
        RECT 64.685000 12.400000 64.885000 12.600000 ;
        RECT 64.685000 12.830000 64.885000 13.030000 ;
        RECT 64.685000 13.260000 64.885000 13.460000 ;
        RECT 65.090000  8.960000 65.290000  9.160000 ;
        RECT 65.090000  9.390000 65.290000  9.590000 ;
        RECT 65.090000  9.820000 65.290000 10.020000 ;
        RECT 65.090000 10.250000 65.290000 10.450000 ;
        RECT 65.090000 10.680000 65.290000 10.880000 ;
        RECT 65.090000 11.110000 65.290000 11.310000 ;
        RECT 65.090000 11.540000 65.290000 11.740000 ;
        RECT 65.090000 11.970000 65.290000 12.170000 ;
        RECT 65.090000 12.400000 65.290000 12.600000 ;
        RECT 65.090000 12.830000 65.290000 13.030000 ;
        RECT 65.090000 13.260000 65.290000 13.460000 ;
        RECT 65.495000  8.960000 65.695000  9.160000 ;
        RECT 65.495000  9.390000 65.695000  9.590000 ;
        RECT 65.495000  9.820000 65.695000 10.020000 ;
        RECT 65.495000 10.250000 65.695000 10.450000 ;
        RECT 65.495000 10.680000 65.695000 10.880000 ;
        RECT 65.495000 11.110000 65.695000 11.310000 ;
        RECT 65.495000 11.540000 65.695000 11.740000 ;
        RECT 65.495000 11.970000 65.695000 12.170000 ;
        RECT 65.495000 12.400000 65.695000 12.600000 ;
        RECT 65.495000 12.830000 65.695000 13.030000 ;
        RECT 65.495000 13.260000 65.695000 13.460000 ;
        RECT 65.900000  8.960000 66.100000  9.160000 ;
        RECT 65.900000  9.390000 66.100000  9.590000 ;
        RECT 65.900000  9.820000 66.100000 10.020000 ;
        RECT 65.900000 10.250000 66.100000 10.450000 ;
        RECT 65.900000 10.680000 66.100000 10.880000 ;
        RECT 65.900000 11.110000 66.100000 11.310000 ;
        RECT 65.900000 11.540000 66.100000 11.740000 ;
        RECT 65.900000 11.970000 66.100000 12.170000 ;
        RECT 65.900000 12.400000 66.100000 12.600000 ;
        RECT 65.900000 12.830000 66.100000 13.030000 ;
        RECT 65.900000 13.260000 66.100000 13.460000 ;
        RECT 66.305000  8.960000 66.505000  9.160000 ;
        RECT 66.305000  9.390000 66.505000  9.590000 ;
        RECT 66.305000  9.820000 66.505000 10.020000 ;
        RECT 66.305000 10.250000 66.505000 10.450000 ;
        RECT 66.305000 10.680000 66.505000 10.880000 ;
        RECT 66.305000 11.110000 66.505000 11.310000 ;
        RECT 66.305000 11.540000 66.505000 11.740000 ;
        RECT 66.305000 11.970000 66.505000 12.170000 ;
        RECT 66.305000 12.400000 66.505000 12.600000 ;
        RECT 66.305000 12.830000 66.505000 13.030000 ;
        RECT 66.305000 13.260000 66.505000 13.460000 ;
        RECT 66.710000  8.960000 66.910000  9.160000 ;
        RECT 66.710000  9.390000 66.910000  9.590000 ;
        RECT 66.710000  9.820000 66.910000 10.020000 ;
        RECT 66.710000 10.250000 66.910000 10.450000 ;
        RECT 66.710000 10.680000 66.910000 10.880000 ;
        RECT 66.710000 11.110000 66.910000 11.310000 ;
        RECT 66.710000 11.540000 66.910000 11.740000 ;
        RECT 66.710000 11.970000 66.910000 12.170000 ;
        RECT 66.710000 12.400000 66.910000 12.600000 ;
        RECT 66.710000 12.830000 66.910000 13.030000 ;
        RECT 66.710000 13.260000 66.910000 13.460000 ;
        RECT 67.115000  8.960000 67.315000  9.160000 ;
        RECT 67.115000  9.390000 67.315000  9.590000 ;
        RECT 67.115000  9.820000 67.315000 10.020000 ;
        RECT 67.115000 10.250000 67.315000 10.450000 ;
        RECT 67.115000 10.680000 67.315000 10.880000 ;
        RECT 67.115000 11.110000 67.315000 11.310000 ;
        RECT 67.115000 11.540000 67.315000 11.740000 ;
        RECT 67.115000 11.970000 67.315000 12.170000 ;
        RECT 67.115000 12.400000 67.315000 12.600000 ;
        RECT 67.115000 12.830000 67.315000 13.030000 ;
        RECT 67.115000 13.260000 67.315000 13.460000 ;
        RECT 67.520000  8.960000 67.720000  9.160000 ;
        RECT 67.520000  9.390000 67.720000  9.590000 ;
        RECT 67.520000  9.820000 67.720000 10.020000 ;
        RECT 67.520000 10.250000 67.720000 10.450000 ;
        RECT 67.520000 10.680000 67.720000 10.880000 ;
        RECT 67.520000 11.110000 67.720000 11.310000 ;
        RECT 67.520000 11.540000 67.720000 11.740000 ;
        RECT 67.520000 11.970000 67.720000 12.170000 ;
        RECT 67.520000 12.400000 67.720000 12.600000 ;
        RECT 67.520000 12.830000 67.720000 13.030000 ;
        RECT 67.520000 13.260000 67.720000 13.460000 ;
        RECT 67.925000  8.960000 68.125000  9.160000 ;
        RECT 67.925000  9.390000 68.125000  9.590000 ;
        RECT 67.925000  9.820000 68.125000 10.020000 ;
        RECT 67.925000 10.250000 68.125000 10.450000 ;
        RECT 67.925000 10.680000 68.125000 10.880000 ;
        RECT 67.925000 11.110000 68.125000 11.310000 ;
        RECT 67.925000 11.540000 68.125000 11.740000 ;
        RECT 67.925000 11.970000 68.125000 12.170000 ;
        RECT 67.925000 12.400000 68.125000 12.600000 ;
        RECT 67.925000 12.830000 68.125000 13.030000 ;
        RECT 67.925000 13.260000 68.125000 13.460000 ;
        RECT 68.330000  8.960000 68.530000  9.160000 ;
        RECT 68.330000  9.390000 68.530000  9.590000 ;
        RECT 68.330000  9.820000 68.530000 10.020000 ;
        RECT 68.330000 10.250000 68.530000 10.450000 ;
        RECT 68.330000 10.680000 68.530000 10.880000 ;
        RECT 68.330000 11.110000 68.530000 11.310000 ;
        RECT 68.330000 11.540000 68.530000 11.740000 ;
        RECT 68.330000 11.970000 68.530000 12.170000 ;
        RECT 68.330000 12.400000 68.530000 12.600000 ;
        RECT 68.330000 12.830000 68.530000 13.030000 ;
        RECT 68.330000 13.260000 68.530000 13.460000 ;
        RECT 68.735000  8.960000 68.935000  9.160000 ;
        RECT 68.735000  9.390000 68.935000  9.590000 ;
        RECT 68.735000  9.820000 68.935000 10.020000 ;
        RECT 68.735000 10.250000 68.935000 10.450000 ;
        RECT 68.735000 10.680000 68.935000 10.880000 ;
        RECT 68.735000 11.110000 68.935000 11.310000 ;
        RECT 68.735000 11.540000 68.935000 11.740000 ;
        RECT 68.735000 11.970000 68.935000 12.170000 ;
        RECT 68.735000 12.400000 68.935000 12.600000 ;
        RECT 68.735000 12.830000 68.935000 13.030000 ;
        RECT 68.735000 13.260000 68.935000 13.460000 ;
        RECT 69.140000  8.960000 69.340000  9.160000 ;
        RECT 69.140000  9.390000 69.340000  9.590000 ;
        RECT 69.140000  9.820000 69.340000 10.020000 ;
        RECT 69.140000 10.250000 69.340000 10.450000 ;
        RECT 69.140000 10.680000 69.340000 10.880000 ;
        RECT 69.140000 11.110000 69.340000 11.310000 ;
        RECT 69.140000 11.540000 69.340000 11.740000 ;
        RECT 69.140000 11.970000 69.340000 12.170000 ;
        RECT 69.140000 12.400000 69.340000 12.600000 ;
        RECT 69.140000 12.830000 69.340000 13.030000 ;
        RECT 69.140000 13.260000 69.340000 13.460000 ;
        RECT 69.545000  8.960000 69.745000  9.160000 ;
        RECT 69.545000  9.390000 69.745000  9.590000 ;
        RECT 69.545000  9.820000 69.745000 10.020000 ;
        RECT 69.545000 10.250000 69.745000 10.450000 ;
        RECT 69.545000 10.680000 69.745000 10.880000 ;
        RECT 69.545000 11.110000 69.745000 11.310000 ;
        RECT 69.545000 11.540000 69.745000 11.740000 ;
        RECT 69.545000 11.970000 69.745000 12.170000 ;
        RECT 69.545000 12.400000 69.745000 12.600000 ;
        RECT 69.545000 12.830000 69.745000 13.030000 ;
        RECT 69.545000 13.260000 69.745000 13.460000 ;
        RECT 69.950000  8.960000 70.150000  9.160000 ;
        RECT 69.950000  9.390000 70.150000  9.590000 ;
        RECT 69.950000  9.820000 70.150000 10.020000 ;
        RECT 69.950000 10.250000 70.150000 10.450000 ;
        RECT 69.950000 10.680000 70.150000 10.880000 ;
        RECT 69.950000 11.110000 70.150000 11.310000 ;
        RECT 69.950000 11.540000 70.150000 11.740000 ;
        RECT 69.950000 11.970000 70.150000 12.170000 ;
        RECT 69.950000 12.400000 70.150000 12.600000 ;
        RECT 69.950000 12.830000 70.150000 13.030000 ;
        RECT 69.950000 13.260000 70.150000 13.460000 ;
        RECT 70.355000  8.960000 70.555000  9.160000 ;
        RECT 70.355000  9.390000 70.555000  9.590000 ;
        RECT 70.355000  9.820000 70.555000 10.020000 ;
        RECT 70.355000 10.250000 70.555000 10.450000 ;
        RECT 70.355000 10.680000 70.555000 10.880000 ;
        RECT 70.355000 11.110000 70.555000 11.310000 ;
        RECT 70.355000 11.540000 70.555000 11.740000 ;
        RECT 70.355000 11.970000 70.555000 12.170000 ;
        RECT 70.355000 12.400000 70.555000 12.600000 ;
        RECT 70.355000 12.830000 70.555000 13.030000 ;
        RECT 70.355000 13.260000 70.555000 13.460000 ;
        RECT 70.760000  8.960000 70.960000  9.160000 ;
        RECT 70.760000  9.390000 70.960000  9.590000 ;
        RECT 70.760000  9.820000 70.960000 10.020000 ;
        RECT 70.760000 10.250000 70.960000 10.450000 ;
        RECT 70.760000 10.680000 70.960000 10.880000 ;
        RECT 70.760000 11.110000 70.960000 11.310000 ;
        RECT 70.760000 11.540000 70.960000 11.740000 ;
        RECT 70.760000 11.970000 70.960000 12.170000 ;
        RECT 70.760000 12.400000 70.960000 12.600000 ;
        RECT 70.760000 12.830000 70.960000 13.030000 ;
        RECT 70.760000 13.260000 70.960000 13.460000 ;
        RECT 71.165000  8.960000 71.365000  9.160000 ;
        RECT 71.165000  9.390000 71.365000  9.590000 ;
        RECT 71.165000  9.820000 71.365000 10.020000 ;
        RECT 71.165000 10.250000 71.365000 10.450000 ;
        RECT 71.165000 10.680000 71.365000 10.880000 ;
        RECT 71.165000 11.110000 71.365000 11.310000 ;
        RECT 71.165000 11.540000 71.365000 11.740000 ;
        RECT 71.165000 11.970000 71.365000 12.170000 ;
        RECT 71.165000 12.400000 71.365000 12.600000 ;
        RECT 71.165000 12.830000 71.365000 13.030000 ;
        RECT 71.165000 13.260000 71.365000 13.460000 ;
        RECT 71.570000  8.960000 71.770000  9.160000 ;
        RECT 71.570000  9.390000 71.770000  9.590000 ;
        RECT 71.570000  9.820000 71.770000 10.020000 ;
        RECT 71.570000 10.250000 71.770000 10.450000 ;
        RECT 71.570000 10.680000 71.770000 10.880000 ;
        RECT 71.570000 11.110000 71.770000 11.310000 ;
        RECT 71.570000 11.540000 71.770000 11.740000 ;
        RECT 71.570000 11.970000 71.770000 12.170000 ;
        RECT 71.570000 12.400000 71.770000 12.600000 ;
        RECT 71.570000 12.830000 71.770000 13.030000 ;
        RECT 71.570000 13.260000 71.770000 13.460000 ;
        RECT 71.975000  8.960000 72.175000  9.160000 ;
        RECT 71.975000  9.390000 72.175000  9.590000 ;
        RECT 71.975000  9.820000 72.175000 10.020000 ;
        RECT 71.975000 10.250000 72.175000 10.450000 ;
        RECT 71.975000 10.680000 72.175000 10.880000 ;
        RECT 71.975000 11.110000 72.175000 11.310000 ;
        RECT 71.975000 11.540000 72.175000 11.740000 ;
        RECT 71.975000 11.970000 72.175000 12.170000 ;
        RECT 71.975000 12.400000 72.175000 12.600000 ;
        RECT 71.975000 12.830000 72.175000 13.030000 ;
        RECT 71.975000 13.260000 72.175000 13.460000 ;
        RECT 72.380000  8.960000 72.580000  9.160000 ;
        RECT 72.380000  9.390000 72.580000  9.590000 ;
        RECT 72.380000  9.820000 72.580000 10.020000 ;
        RECT 72.380000 10.250000 72.580000 10.450000 ;
        RECT 72.380000 10.680000 72.580000 10.880000 ;
        RECT 72.380000 11.110000 72.580000 11.310000 ;
        RECT 72.380000 11.540000 72.580000 11.740000 ;
        RECT 72.380000 11.970000 72.580000 12.170000 ;
        RECT 72.380000 12.400000 72.580000 12.600000 ;
        RECT 72.380000 12.830000 72.580000 13.030000 ;
        RECT 72.380000 13.260000 72.580000 13.460000 ;
        RECT 72.785000  8.960000 72.985000  9.160000 ;
        RECT 72.785000  9.390000 72.985000  9.590000 ;
        RECT 72.785000  9.820000 72.985000 10.020000 ;
        RECT 72.785000 10.250000 72.985000 10.450000 ;
        RECT 72.785000 10.680000 72.985000 10.880000 ;
        RECT 72.785000 11.110000 72.985000 11.310000 ;
        RECT 72.785000 11.540000 72.985000 11.740000 ;
        RECT 72.785000 11.970000 72.985000 12.170000 ;
        RECT 72.785000 12.400000 72.985000 12.600000 ;
        RECT 72.785000 12.830000 72.985000 13.030000 ;
        RECT 72.785000 13.260000 72.985000 13.460000 ;
        RECT 73.190000  8.960000 73.390000  9.160000 ;
        RECT 73.190000  9.390000 73.390000  9.590000 ;
        RECT 73.190000  9.820000 73.390000 10.020000 ;
        RECT 73.190000 10.250000 73.390000 10.450000 ;
        RECT 73.190000 10.680000 73.390000 10.880000 ;
        RECT 73.190000 11.110000 73.390000 11.310000 ;
        RECT 73.190000 11.540000 73.390000 11.740000 ;
        RECT 73.190000 11.970000 73.390000 12.170000 ;
        RECT 73.190000 12.400000 73.390000 12.600000 ;
        RECT 73.190000 12.830000 73.390000 13.030000 ;
        RECT 73.190000 13.260000 73.390000 13.460000 ;
        RECT 73.595000  8.960000 73.795000  9.160000 ;
        RECT 73.595000  9.390000 73.795000  9.590000 ;
        RECT 73.595000  9.820000 73.795000 10.020000 ;
        RECT 73.595000 10.250000 73.795000 10.450000 ;
        RECT 73.595000 10.680000 73.795000 10.880000 ;
        RECT 73.595000 11.110000 73.795000 11.310000 ;
        RECT 73.595000 11.540000 73.795000 11.740000 ;
        RECT 73.595000 11.970000 73.795000 12.170000 ;
        RECT 73.595000 12.400000 73.795000 12.600000 ;
        RECT 73.595000 12.830000 73.795000 13.030000 ;
        RECT 73.595000 13.260000 73.795000 13.460000 ;
        RECT 74.000000  8.960000 74.200000  9.160000 ;
        RECT 74.000000  9.390000 74.200000  9.590000 ;
        RECT 74.000000  9.820000 74.200000 10.020000 ;
        RECT 74.000000 10.250000 74.200000 10.450000 ;
        RECT 74.000000 10.680000 74.200000 10.880000 ;
        RECT 74.000000 11.110000 74.200000 11.310000 ;
        RECT 74.000000 11.540000 74.200000 11.740000 ;
        RECT 74.000000 11.970000 74.200000 12.170000 ;
        RECT 74.000000 12.400000 74.200000 12.600000 ;
        RECT 74.000000 12.830000 74.200000 13.030000 ;
        RECT 74.000000 13.260000 74.200000 13.460000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
  END
END sky130_fd_io__overlay_vccd_hvc


MACRO sky130_fd_io__overlay_vdda_hvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.495000 14.940000 24.395000 18.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 14.940000 74.290000 18.380000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 24.370000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.585000 15.020000  0.785000 15.220000 ;
        RECT  0.585000 15.460000  0.785000 15.660000 ;
        RECT  0.585000 15.900000  0.785000 16.100000 ;
        RECT  0.585000 16.340000  0.785000 16.540000 ;
        RECT  0.585000 16.780000  0.785000 16.980000 ;
        RECT  0.585000 17.220000  0.785000 17.420000 ;
        RECT  0.585000 17.660000  0.785000 17.860000 ;
        RECT  0.585000 18.100000  0.785000 18.300000 ;
        RECT  0.995000 15.020000  1.195000 15.220000 ;
        RECT  0.995000 15.460000  1.195000 15.660000 ;
        RECT  0.995000 15.900000  1.195000 16.100000 ;
        RECT  0.995000 16.340000  1.195000 16.540000 ;
        RECT  0.995000 16.780000  1.195000 16.980000 ;
        RECT  0.995000 17.220000  1.195000 17.420000 ;
        RECT  0.995000 17.660000  1.195000 17.860000 ;
        RECT  0.995000 18.100000  1.195000 18.300000 ;
        RECT  1.405000 15.020000  1.605000 15.220000 ;
        RECT  1.405000 15.460000  1.605000 15.660000 ;
        RECT  1.405000 15.900000  1.605000 16.100000 ;
        RECT  1.405000 16.340000  1.605000 16.540000 ;
        RECT  1.405000 16.780000  1.605000 16.980000 ;
        RECT  1.405000 17.220000  1.605000 17.420000 ;
        RECT  1.405000 17.660000  1.605000 17.860000 ;
        RECT  1.405000 18.100000  1.605000 18.300000 ;
        RECT  1.815000 15.020000  2.015000 15.220000 ;
        RECT  1.815000 15.460000  2.015000 15.660000 ;
        RECT  1.815000 15.900000  2.015000 16.100000 ;
        RECT  1.815000 16.340000  2.015000 16.540000 ;
        RECT  1.815000 16.780000  2.015000 16.980000 ;
        RECT  1.815000 17.220000  2.015000 17.420000 ;
        RECT  1.815000 17.660000  2.015000 17.860000 ;
        RECT  1.815000 18.100000  2.015000 18.300000 ;
        RECT  2.225000 15.020000  2.425000 15.220000 ;
        RECT  2.225000 15.460000  2.425000 15.660000 ;
        RECT  2.225000 15.900000  2.425000 16.100000 ;
        RECT  2.225000 16.340000  2.425000 16.540000 ;
        RECT  2.225000 16.780000  2.425000 16.980000 ;
        RECT  2.225000 17.220000  2.425000 17.420000 ;
        RECT  2.225000 17.660000  2.425000 17.860000 ;
        RECT  2.225000 18.100000  2.425000 18.300000 ;
        RECT  2.635000 15.020000  2.835000 15.220000 ;
        RECT  2.635000 15.460000  2.835000 15.660000 ;
        RECT  2.635000 15.900000  2.835000 16.100000 ;
        RECT  2.635000 16.340000  2.835000 16.540000 ;
        RECT  2.635000 16.780000  2.835000 16.980000 ;
        RECT  2.635000 17.220000  2.835000 17.420000 ;
        RECT  2.635000 17.660000  2.835000 17.860000 ;
        RECT  2.635000 18.100000  2.835000 18.300000 ;
        RECT  3.045000 15.020000  3.245000 15.220000 ;
        RECT  3.045000 15.460000  3.245000 15.660000 ;
        RECT  3.045000 15.900000  3.245000 16.100000 ;
        RECT  3.045000 16.340000  3.245000 16.540000 ;
        RECT  3.045000 16.780000  3.245000 16.980000 ;
        RECT  3.045000 17.220000  3.245000 17.420000 ;
        RECT  3.045000 17.660000  3.245000 17.860000 ;
        RECT  3.045000 18.100000  3.245000 18.300000 ;
        RECT  3.450000 15.020000  3.650000 15.220000 ;
        RECT  3.450000 15.460000  3.650000 15.660000 ;
        RECT  3.450000 15.900000  3.650000 16.100000 ;
        RECT  3.450000 16.340000  3.650000 16.540000 ;
        RECT  3.450000 16.780000  3.650000 16.980000 ;
        RECT  3.450000 17.220000  3.650000 17.420000 ;
        RECT  3.450000 17.660000  3.650000 17.860000 ;
        RECT  3.450000 18.100000  3.650000 18.300000 ;
        RECT  3.855000 15.020000  4.055000 15.220000 ;
        RECT  3.855000 15.460000  4.055000 15.660000 ;
        RECT  3.855000 15.900000  4.055000 16.100000 ;
        RECT  3.855000 16.340000  4.055000 16.540000 ;
        RECT  3.855000 16.780000  4.055000 16.980000 ;
        RECT  3.855000 17.220000  4.055000 17.420000 ;
        RECT  3.855000 17.660000  4.055000 17.860000 ;
        RECT  3.855000 18.100000  4.055000 18.300000 ;
        RECT  4.260000 15.020000  4.460000 15.220000 ;
        RECT  4.260000 15.460000  4.460000 15.660000 ;
        RECT  4.260000 15.900000  4.460000 16.100000 ;
        RECT  4.260000 16.340000  4.460000 16.540000 ;
        RECT  4.260000 16.780000  4.460000 16.980000 ;
        RECT  4.260000 17.220000  4.460000 17.420000 ;
        RECT  4.260000 17.660000  4.460000 17.860000 ;
        RECT  4.260000 18.100000  4.460000 18.300000 ;
        RECT  4.665000 15.020000  4.865000 15.220000 ;
        RECT  4.665000 15.460000  4.865000 15.660000 ;
        RECT  4.665000 15.900000  4.865000 16.100000 ;
        RECT  4.665000 16.340000  4.865000 16.540000 ;
        RECT  4.665000 16.780000  4.865000 16.980000 ;
        RECT  4.665000 17.220000  4.865000 17.420000 ;
        RECT  4.665000 17.660000  4.865000 17.860000 ;
        RECT  4.665000 18.100000  4.865000 18.300000 ;
        RECT  5.070000 15.020000  5.270000 15.220000 ;
        RECT  5.070000 15.460000  5.270000 15.660000 ;
        RECT  5.070000 15.900000  5.270000 16.100000 ;
        RECT  5.070000 16.340000  5.270000 16.540000 ;
        RECT  5.070000 16.780000  5.270000 16.980000 ;
        RECT  5.070000 17.220000  5.270000 17.420000 ;
        RECT  5.070000 17.660000  5.270000 17.860000 ;
        RECT  5.070000 18.100000  5.270000 18.300000 ;
        RECT  5.475000 15.020000  5.675000 15.220000 ;
        RECT  5.475000 15.460000  5.675000 15.660000 ;
        RECT  5.475000 15.900000  5.675000 16.100000 ;
        RECT  5.475000 16.340000  5.675000 16.540000 ;
        RECT  5.475000 16.780000  5.675000 16.980000 ;
        RECT  5.475000 17.220000  5.675000 17.420000 ;
        RECT  5.475000 17.660000  5.675000 17.860000 ;
        RECT  5.475000 18.100000  5.675000 18.300000 ;
        RECT  5.880000 15.020000  6.080000 15.220000 ;
        RECT  5.880000 15.460000  6.080000 15.660000 ;
        RECT  5.880000 15.900000  6.080000 16.100000 ;
        RECT  5.880000 16.340000  6.080000 16.540000 ;
        RECT  5.880000 16.780000  6.080000 16.980000 ;
        RECT  5.880000 17.220000  6.080000 17.420000 ;
        RECT  5.880000 17.660000  6.080000 17.860000 ;
        RECT  5.880000 18.100000  6.080000 18.300000 ;
        RECT  6.285000 15.020000  6.485000 15.220000 ;
        RECT  6.285000 15.460000  6.485000 15.660000 ;
        RECT  6.285000 15.900000  6.485000 16.100000 ;
        RECT  6.285000 16.340000  6.485000 16.540000 ;
        RECT  6.285000 16.780000  6.485000 16.980000 ;
        RECT  6.285000 17.220000  6.485000 17.420000 ;
        RECT  6.285000 17.660000  6.485000 17.860000 ;
        RECT  6.285000 18.100000  6.485000 18.300000 ;
        RECT  6.690000 15.020000  6.890000 15.220000 ;
        RECT  6.690000 15.460000  6.890000 15.660000 ;
        RECT  6.690000 15.900000  6.890000 16.100000 ;
        RECT  6.690000 16.340000  6.890000 16.540000 ;
        RECT  6.690000 16.780000  6.890000 16.980000 ;
        RECT  6.690000 17.220000  6.890000 17.420000 ;
        RECT  6.690000 17.660000  6.890000 17.860000 ;
        RECT  6.690000 18.100000  6.890000 18.300000 ;
        RECT  7.095000 15.020000  7.295000 15.220000 ;
        RECT  7.095000 15.460000  7.295000 15.660000 ;
        RECT  7.095000 15.900000  7.295000 16.100000 ;
        RECT  7.095000 16.340000  7.295000 16.540000 ;
        RECT  7.095000 16.780000  7.295000 16.980000 ;
        RECT  7.095000 17.220000  7.295000 17.420000 ;
        RECT  7.095000 17.660000  7.295000 17.860000 ;
        RECT  7.095000 18.100000  7.295000 18.300000 ;
        RECT  7.500000 15.020000  7.700000 15.220000 ;
        RECT  7.500000 15.460000  7.700000 15.660000 ;
        RECT  7.500000 15.900000  7.700000 16.100000 ;
        RECT  7.500000 16.340000  7.700000 16.540000 ;
        RECT  7.500000 16.780000  7.700000 16.980000 ;
        RECT  7.500000 17.220000  7.700000 17.420000 ;
        RECT  7.500000 17.660000  7.700000 17.860000 ;
        RECT  7.500000 18.100000  7.700000 18.300000 ;
        RECT  7.905000 15.020000  8.105000 15.220000 ;
        RECT  7.905000 15.460000  8.105000 15.660000 ;
        RECT  7.905000 15.900000  8.105000 16.100000 ;
        RECT  7.905000 16.340000  8.105000 16.540000 ;
        RECT  7.905000 16.780000  8.105000 16.980000 ;
        RECT  7.905000 17.220000  8.105000 17.420000 ;
        RECT  7.905000 17.660000  8.105000 17.860000 ;
        RECT  7.905000 18.100000  8.105000 18.300000 ;
        RECT  8.310000 15.020000  8.510000 15.220000 ;
        RECT  8.310000 15.460000  8.510000 15.660000 ;
        RECT  8.310000 15.900000  8.510000 16.100000 ;
        RECT  8.310000 16.340000  8.510000 16.540000 ;
        RECT  8.310000 16.780000  8.510000 16.980000 ;
        RECT  8.310000 17.220000  8.510000 17.420000 ;
        RECT  8.310000 17.660000  8.510000 17.860000 ;
        RECT  8.310000 18.100000  8.510000 18.300000 ;
        RECT  8.715000 15.020000  8.915000 15.220000 ;
        RECT  8.715000 15.460000  8.915000 15.660000 ;
        RECT  8.715000 15.900000  8.915000 16.100000 ;
        RECT  8.715000 16.340000  8.915000 16.540000 ;
        RECT  8.715000 16.780000  8.915000 16.980000 ;
        RECT  8.715000 17.220000  8.915000 17.420000 ;
        RECT  8.715000 17.660000  8.915000 17.860000 ;
        RECT  8.715000 18.100000  8.915000 18.300000 ;
        RECT  9.120000 15.020000  9.320000 15.220000 ;
        RECT  9.120000 15.460000  9.320000 15.660000 ;
        RECT  9.120000 15.900000  9.320000 16.100000 ;
        RECT  9.120000 16.340000  9.320000 16.540000 ;
        RECT  9.120000 16.780000  9.320000 16.980000 ;
        RECT  9.120000 17.220000  9.320000 17.420000 ;
        RECT  9.120000 17.660000  9.320000 17.860000 ;
        RECT  9.120000 18.100000  9.320000 18.300000 ;
        RECT  9.525000 15.020000  9.725000 15.220000 ;
        RECT  9.525000 15.460000  9.725000 15.660000 ;
        RECT  9.525000 15.900000  9.725000 16.100000 ;
        RECT  9.525000 16.340000  9.725000 16.540000 ;
        RECT  9.525000 16.780000  9.725000 16.980000 ;
        RECT  9.525000 17.220000  9.725000 17.420000 ;
        RECT  9.525000 17.660000  9.725000 17.860000 ;
        RECT  9.525000 18.100000  9.725000 18.300000 ;
        RECT  9.930000 15.020000 10.130000 15.220000 ;
        RECT  9.930000 15.460000 10.130000 15.660000 ;
        RECT  9.930000 15.900000 10.130000 16.100000 ;
        RECT  9.930000 16.340000 10.130000 16.540000 ;
        RECT  9.930000 16.780000 10.130000 16.980000 ;
        RECT  9.930000 17.220000 10.130000 17.420000 ;
        RECT  9.930000 17.660000 10.130000 17.860000 ;
        RECT  9.930000 18.100000 10.130000 18.300000 ;
        RECT 10.335000 15.020000 10.535000 15.220000 ;
        RECT 10.335000 15.460000 10.535000 15.660000 ;
        RECT 10.335000 15.900000 10.535000 16.100000 ;
        RECT 10.335000 16.340000 10.535000 16.540000 ;
        RECT 10.335000 16.780000 10.535000 16.980000 ;
        RECT 10.335000 17.220000 10.535000 17.420000 ;
        RECT 10.335000 17.660000 10.535000 17.860000 ;
        RECT 10.335000 18.100000 10.535000 18.300000 ;
        RECT 10.740000 15.020000 10.940000 15.220000 ;
        RECT 10.740000 15.460000 10.940000 15.660000 ;
        RECT 10.740000 15.900000 10.940000 16.100000 ;
        RECT 10.740000 16.340000 10.940000 16.540000 ;
        RECT 10.740000 16.780000 10.940000 16.980000 ;
        RECT 10.740000 17.220000 10.940000 17.420000 ;
        RECT 10.740000 17.660000 10.940000 17.860000 ;
        RECT 10.740000 18.100000 10.940000 18.300000 ;
        RECT 11.145000 15.020000 11.345000 15.220000 ;
        RECT 11.145000 15.460000 11.345000 15.660000 ;
        RECT 11.145000 15.900000 11.345000 16.100000 ;
        RECT 11.145000 16.340000 11.345000 16.540000 ;
        RECT 11.145000 16.780000 11.345000 16.980000 ;
        RECT 11.145000 17.220000 11.345000 17.420000 ;
        RECT 11.145000 17.660000 11.345000 17.860000 ;
        RECT 11.145000 18.100000 11.345000 18.300000 ;
        RECT 11.550000 15.020000 11.750000 15.220000 ;
        RECT 11.550000 15.460000 11.750000 15.660000 ;
        RECT 11.550000 15.900000 11.750000 16.100000 ;
        RECT 11.550000 16.340000 11.750000 16.540000 ;
        RECT 11.550000 16.780000 11.750000 16.980000 ;
        RECT 11.550000 17.220000 11.750000 17.420000 ;
        RECT 11.550000 17.660000 11.750000 17.860000 ;
        RECT 11.550000 18.100000 11.750000 18.300000 ;
        RECT 11.955000 15.020000 12.155000 15.220000 ;
        RECT 11.955000 15.460000 12.155000 15.660000 ;
        RECT 11.955000 15.900000 12.155000 16.100000 ;
        RECT 11.955000 16.340000 12.155000 16.540000 ;
        RECT 11.955000 16.780000 12.155000 16.980000 ;
        RECT 11.955000 17.220000 12.155000 17.420000 ;
        RECT 11.955000 17.660000 12.155000 17.860000 ;
        RECT 11.955000 18.100000 12.155000 18.300000 ;
        RECT 12.360000 15.020000 12.560000 15.220000 ;
        RECT 12.360000 15.460000 12.560000 15.660000 ;
        RECT 12.360000 15.900000 12.560000 16.100000 ;
        RECT 12.360000 16.340000 12.560000 16.540000 ;
        RECT 12.360000 16.780000 12.560000 16.980000 ;
        RECT 12.360000 17.220000 12.560000 17.420000 ;
        RECT 12.360000 17.660000 12.560000 17.860000 ;
        RECT 12.360000 18.100000 12.560000 18.300000 ;
        RECT 12.765000 15.020000 12.965000 15.220000 ;
        RECT 12.765000 15.460000 12.965000 15.660000 ;
        RECT 12.765000 15.900000 12.965000 16.100000 ;
        RECT 12.765000 16.340000 12.965000 16.540000 ;
        RECT 12.765000 16.780000 12.965000 16.980000 ;
        RECT 12.765000 17.220000 12.965000 17.420000 ;
        RECT 12.765000 17.660000 12.965000 17.860000 ;
        RECT 12.765000 18.100000 12.965000 18.300000 ;
        RECT 13.170000 15.020000 13.370000 15.220000 ;
        RECT 13.170000 15.460000 13.370000 15.660000 ;
        RECT 13.170000 15.900000 13.370000 16.100000 ;
        RECT 13.170000 16.340000 13.370000 16.540000 ;
        RECT 13.170000 16.780000 13.370000 16.980000 ;
        RECT 13.170000 17.220000 13.370000 17.420000 ;
        RECT 13.170000 17.660000 13.370000 17.860000 ;
        RECT 13.170000 18.100000 13.370000 18.300000 ;
        RECT 13.575000 15.020000 13.775000 15.220000 ;
        RECT 13.575000 15.460000 13.775000 15.660000 ;
        RECT 13.575000 15.900000 13.775000 16.100000 ;
        RECT 13.575000 16.340000 13.775000 16.540000 ;
        RECT 13.575000 16.780000 13.775000 16.980000 ;
        RECT 13.575000 17.220000 13.775000 17.420000 ;
        RECT 13.575000 17.660000 13.775000 17.860000 ;
        RECT 13.575000 18.100000 13.775000 18.300000 ;
        RECT 13.980000 15.020000 14.180000 15.220000 ;
        RECT 13.980000 15.460000 14.180000 15.660000 ;
        RECT 13.980000 15.900000 14.180000 16.100000 ;
        RECT 13.980000 16.340000 14.180000 16.540000 ;
        RECT 13.980000 16.780000 14.180000 16.980000 ;
        RECT 13.980000 17.220000 14.180000 17.420000 ;
        RECT 13.980000 17.660000 14.180000 17.860000 ;
        RECT 13.980000 18.100000 14.180000 18.300000 ;
        RECT 14.385000 15.020000 14.585000 15.220000 ;
        RECT 14.385000 15.460000 14.585000 15.660000 ;
        RECT 14.385000 15.900000 14.585000 16.100000 ;
        RECT 14.385000 16.340000 14.585000 16.540000 ;
        RECT 14.385000 16.780000 14.585000 16.980000 ;
        RECT 14.385000 17.220000 14.585000 17.420000 ;
        RECT 14.385000 17.660000 14.585000 17.860000 ;
        RECT 14.385000 18.100000 14.585000 18.300000 ;
        RECT 14.790000 15.020000 14.990000 15.220000 ;
        RECT 14.790000 15.460000 14.990000 15.660000 ;
        RECT 14.790000 15.900000 14.990000 16.100000 ;
        RECT 14.790000 16.340000 14.990000 16.540000 ;
        RECT 14.790000 16.780000 14.990000 16.980000 ;
        RECT 14.790000 17.220000 14.990000 17.420000 ;
        RECT 14.790000 17.660000 14.990000 17.860000 ;
        RECT 14.790000 18.100000 14.990000 18.300000 ;
        RECT 15.195000 15.020000 15.395000 15.220000 ;
        RECT 15.195000 15.460000 15.395000 15.660000 ;
        RECT 15.195000 15.900000 15.395000 16.100000 ;
        RECT 15.195000 16.340000 15.395000 16.540000 ;
        RECT 15.195000 16.780000 15.395000 16.980000 ;
        RECT 15.195000 17.220000 15.395000 17.420000 ;
        RECT 15.195000 17.660000 15.395000 17.860000 ;
        RECT 15.195000 18.100000 15.395000 18.300000 ;
        RECT 15.600000 15.020000 15.800000 15.220000 ;
        RECT 15.600000 15.460000 15.800000 15.660000 ;
        RECT 15.600000 15.900000 15.800000 16.100000 ;
        RECT 15.600000 16.340000 15.800000 16.540000 ;
        RECT 15.600000 16.780000 15.800000 16.980000 ;
        RECT 15.600000 17.220000 15.800000 17.420000 ;
        RECT 15.600000 17.660000 15.800000 17.860000 ;
        RECT 15.600000 18.100000 15.800000 18.300000 ;
        RECT 16.005000 15.020000 16.205000 15.220000 ;
        RECT 16.005000 15.460000 16.205000 15.660000 ;
        RECT 16.005000 15.900000 16.205000 16.100000 ;
        RECT 16.005000 16.340000 16.205000 16.540000 ;
        RECT 16.005000 16.780000 16.205000 16.980000 ;
        RECT 16.005000 17.220000 16.205000 17.420000 ;
        RECT 16.005000 17.660000 16.205000 17.860000 ;
        RECT 16.005000 18.100000 16.205000 18.300000 ;
        RECT 16.410000 15.020000 16.610000 15.220000 ;
        RECT 16.410000 15.460000 16.610000 15.660000 ;
        RECT 16.410000 15.900000 16.610000 16.100000 ;
        RECT 16.410000 16.340000 16.610000 16.540000 ;
        RECT 16.410000 16.780000 16.610000 16.980000 ;
        RECT 16.410000 17.220000 16.610000 17.420000 ;
        RECT 16.410000 17.660000 16.610000 17.860000 ;
        RECT 16.410000 18.100000 16.610000 18.300000 ;
        RECT 16.815000 15.020000 17.015000 15.220000 ;
        RECT 16.815000 15.460000 17.015000 15.660000 ;
        RECT 16.815000 15.900000 17.015000 16.100000 ;
        RECT 16.815000 16.340000 17.015000 16.540000 ;
        RECT 16.815000 16.780000 17.015000 16.980000 ;
        RECT 16.815000 17.220000 17.015000 17.420000 ;
        RECT 16.815000 17.660000 17.015000 17.860000 ;
        RECT 16.815000 18.100000 17.015000 18.300000 ;
        RECT 17.220000 15.020000 17.420000 15.220000 ;
        RECT 17.220000 15.460000 17.420000 15.660000 ;
        RECT 17.220000 15.900000 17.420000 16.100000 ;
        RECT 17.220000 16.340000 17.420000 16.540000 ;
        RECT 17.220000 16.780000 17.420000 16.980000 ;
        RECT 17.220000 17.220000 17.420000 17.420000 ;
        RECT 17.220000 17.660000 17.420000 17.860000 ;
        RECT 17.220000 18.100000 17.420000 18.300000 ;
        RECT 17.625000 15.020000 17.825000 15.220000 ;
        RECT 17.625000 15.460000 17.825000 15.660000 ;
        RECT 17.625000 15.900000 17.825000 16.100000 ;
        RECT 17.625000 16.340000 17.825000 16.540000 ;
        RECT 17.625000 16.780000 17.825000 16.980000 ;
        RECT 17.625000 17.220000 17.825000 17.420000 ;
        RECT 17.625000 17.660000 17.825000 17.860000 ;
        RECT 17.625000 18.100000 17.825000 18.300000 ;
        RECT 18.030000 15.020000 18.230000 15.220000 ;
        RECT 18.030000 15.460000 18.230000 15.660000 ;
        RECT 18.030000 15.900000 18.230000 16.100000 ;
        RECT 18.030000 16.340000 18.230000 16.540000 ;
        RECT 18.030000 16.780000 18.230000 16.980000 ;
        RECT 18.030000 17.220000 18.230000 17.420000 ;
        RECT 18.030000 17.660000 18.230000 17.860000 ;
        RECT 18.030000 18.100000 18.230000 18.300000 ;
        RECT 18.435000 15.020000 18.635000 15.220000 ;
        RECT 18.435000 15.460000 18.635000 15.660000 ;
        RECT 18.435000 15.900000 18.635000 16.100000 ;
        RECT 18.435000 16.340000 18.635000 16.540000 ;
        RECT 18.435000 16.780000 18.635000 16.980000 ;
        RECT 18.435000 17.220000 18.635000 17.420000 ;
        RECT 18.435000 17.660000 18.635000 17.860000 ;
        RECT 18.435000 18.100000 18.635000 18.300000 ;
        RECT 18.840000 15.020000 19.040000 15.220000 ;
        RECT 18.840000 15.460000 19.040000 15.660000 ;
        RECT 18.840000 15.900000 19.040000 16.100000 ;
        RECT 18.840000 16.340000 19.040000 16.540000 ;
        RECT 18.840000 16.780000 19.040000 16.980000 ;
        RECT 18.840000 17.220000 19.040000 17.420000 ;
        RECT 18.840000 17.660000 19.040000 17.860000 ;
        RECT 18.840000 18.100000 19.040000 18.300000 ;
        RECT 19.245000 15.020000 19.445000 15.220000 ;
        RECT 19.245000 15.460000 19.445000 15.660000 ;
        RECT 19.245000 15.900000 19.445000 16.100000 ;
        RECT 19.245000 16.340000 19.445000 16.540000 ;
        RECT 19.245000 16.780000 19.445000 16.980000 ;
        RECT 19.245000 17.220000 19.445000 17.420000 ;
        RECT 19.245000 17.660000 19.445000 17.860000 ;
        RECT 19.245000 18.100000 19.445000 18.300000 ;
        RECT 19.650000 15.020000 19.850000 15.220000 ;
        RECT 19.650000 15.460000 19.850000 15.660000 ;
        RECT 19.650000 15.900000 19.850000 16.100000 ;
        RECT 19.650000 16.340000 19.850000 16.540000 ;
        RECT 19.650000 16.780000 19.850000 16.980000 ;
        RECT 19.650000 17.220000 19.850000 17.420000 ;
        RECT 19.650000 17.660000 19.850000 17.860000 ;
        RECT 19.650000 18.100000 19.850000 18.300000 ;
        RECT 20.055000 15.020000 20.255000 15.220000 ;
        RECT 20.055000 15.460000 20.255000 15.660000 ;
        RECT 20.055000 15.900000 20.255000 16.100000 ;
        RECT 20.055000 16.340000 20.255000 16.540000 ;
        RECT 20.055000 16.780000 20.255000 16.980000 ;
        RECT 20.055000 17.220000 20.255000 17.420000 ;
        RECT 20.055000 17.660000 20.255000 17.860000 ;
        RECT 20.055000 18.100000 20.255000 18.300000 ;
        RECT 20.460000 15.020000 20.660000 15.220000 ;
        RECT 20.460000 15.460000 20.660000 15.660000 ;
        RECT 20.460000 15.900000 20.660000 16.100000 ;
        RECT 20.460000 16.340000 20.660000 16.540000 ;
        RECT 20.460000 16.780000 20.660000 16.980000 ;
        RECT 20.460000 17.220000 20.660000 17.420000 ;
        RECT 20.460000 17.660000 20.660000 17.860000 ;
        RECT 20.460000 18.100000 20.660000 18.300000 ;
        RECT 20.865000 15.020000 21.065000 15.220000 ;
        RECT 20.865000 15.460000 21.065000 15.660000 ;
        RECT 20.865000 15.900000 21.065000 16.100000 ;
        RECT 20.865000 16.340000 21.065000 16.540000 ;
        RECT 20.865000 16.780000 21.065000 16.980000 ;
        RECT 20.865000 17.220000 21.065000 17.420000 ;
        RECT 20.865000 17.660000 21.065000 17.860000 ;
        RECT 20.865000 18.100000 21.065000 18.300000 ;
        RECT 21.270000 15.020000 21.470000 15.220000 ;
        RECT 21.270000 15.460000 21.470000 15.660000 ;
        RECT 21.270000 15.900000 21.470000 16.100000 ;
        RECT 21.270000 16.340000 21.470000 16.540000 ;
        RECT 21.270000 16.780000 21.470000 16.980000 ;
        RECT 21.270000 17.220000 21.470000 17.420000 ;
        RECT 21.270000 17.660000 21.470000 17.860000 ;
        RECT 21.270000 18.100000 21.470000 18.300000 ;
        RECT 21.675000 15.020000 21.875000 15.220000 ;
        RECT 21.675000 15.460000 21.875000 15.660000 ;
        RECT 21.675000 15.900000 21.875000 16.100000 ;
        RECT 21.675000 16.340000 21.875000 16.540000 ;
        RECT 21.675000 16.780000 21.875000 16.980000 ;
        RECT 21.675000 17.220000 21.875000 17.420000 ;
        RECT 21.675000 17.660000 21.875000 17.860000 ;
        RECT 21.675000 18.100000 21.875000 18.300000 ;
        RECT 22.080000 15.020000 22.280000 15.220000 ;
        RECT 22.080000 15.460000 22.280000 15.660000 ;
        RECT 22.080000 15.900000 22.280000 16.100000 ;
        RECT 22.080000 16.340000 22.280000 16.540000 ;
        RECT 22.080000 16.780000 22.280000 16.980000 ;
        RECT 22.080000 17.220000 22.280000 17.420000 ;
        RECT 22.080000 17.660000 22.280000 17.860000 ;
        RECT 22.080000 18.100000 22.280000 18.300000 ;
        RECT 22.485000 15.020000 22.685000 15.220000 ;
        RECT 22.485000 15.460000 22.685000 15.660000 ;
        RECT 22.485000 15.900000 22.685000 16.100000 ;
        RECT 22.485000 16.340000 22.685000 16.540000 ;
        RECT 22.485000 16.780000 22.685000 16.980000 ;
        RECT 22.485000 17.220000 22.685000 17.420000 ;
        RECT 22.485000 17.660000 22.685000 17.860000 ;
        RECT 22.485000 18.100000 22.685000 18.300000 ;
        RECT 22.890000 15.020000 23.090000 15.220000 ;
        RECT 22.890000 15.460000 23.090000 15.660000 ;
        RECT 22.890000 15.900000 23.090000 16.100000 ;
        RECT 22.890000 16.340000 23.090000 16.540000 ;
        RECT 22.890000 16.780000 23.090000 16.980000 ;
        RECT 22.890000 17.220000 23.090000 17.420000 ;
        RECT 22.890000 17.660000 23.090000 17.860000 ;
        RECT 22.890000 18.100000 23.090000 18.300000 ;
        RECT 23.295000 15.020000 23.495000 15.220000 ;
        RECT 23.295000 15.460000 23.495000 15.660000 ;
        RECT 23.295000 15.900000 23.495000 16.100000 ;
        RECT 23.295000 16.340000 23.495000 16.540000 ;
        RECT 23.295000 16.780000 23.495000 16.980000 ;
        RECT 23.295000 17.220000 23.495000 17.420000 ;
        RECT 23.295000 17.660000 23.495000 17.860000 ;
        RECT 23.295000 18.100000 23.495000 18.300000 ;
        RECT 23.700000 15.020000 23.900000 15.220000 ;
        RECT 23.700000 15.460000 23.900000 15.660000 ;
        RECT 23.700000 15.900000 23.900000 16.100000 ;
        RECT 23.700000 16.340000 23.900000 16.540000 ;
        RECT 23.700000 16.780000 23.900000 16.980000 ;
        RECT 23.700000 17.220000 23.900000 17.420000 ;
        RECT 23.700000 17.660000 23.900000 17.860000 ;
        RECT 23.700000 18.100000 23.900000 18.300000 ;
        RECT 24.105000 15.020000 24.305000 15.220000 ;
        RECT 24.105000 15.460000 24.305000 15.660000 ;
        RECT 24.105000 15.900000 24.305000 16.100000 ;
        RECT 24.105000 16.340000 24.305000 16.540000 ;
        RECT 24.105000 16.780000 24.305000 16.980000 ;
        RECT 24.105000 17.220000 24.305000 17.420000 ;
        RECT 24.105000 17.660000 24.305000 17.860000 ;
        RECT 24.105000 18.100000 24.305000 18.300000 ;
        RECT 50.480000 15.020000 50.680000 15.220000 ;
        RECT 50.480000 15.460000 50.680000 15.660000 ;
        RECT 50.480000 15.900000 50.680000 16.100000 ;
        RECT 50.480000 16.340000 50.680000 16.540000 ;
        RECT 50.480000 16.780000 50.680000 16.980000 ;
        RECT 50.480000 17.220000 50.680000 17.420000 ;
        RECT 50.480000 17.660000 50.680000 17.860000 ;
        RECT 50.480000 18.100000 50.680000 18.300000 ;
        RECT 50.890000 15.020000 51.090000 15.220000 ;
        RECT 50.890000 15.460000 51.090000 15.660000 ;
        RECT 50.890000 15.900000 51.090000 16.100000 ;
        RECT 50.890000 16.340000 51.090000 16.540000 ;
        RECT 50.890000 16.780000 51.090000 16.980000 ;
        RECT 50.890000 17.220000 51.090000 17.420000 ;
        RECT 50.890000 17.660000 51.090000 17.860000 ;
        RECT 50.890000 18.100000 51.090000 18.300000 ;
        RECT 51.300000 15.020000 51.500000 15.220000 ;
        RECT 51.300000 15.460000 51.500000 15.660000 ;
        RECT 51.300000 15.900000 51.500000 16.100000 ;
        RECT 51.300000 16.340000 51.500000 16.540000 ;
        RECT 51.300000 16.780000 51.500000 16.980000 ;
        RECT 51.300000 17.220000 51.500000 17.420000 ;
        RECT 51.300000 17.660000 51.500000 17.860000 ;
        RECT 51.300000 18.100000 51.500000 18.300000 ;
        RECT 51.710000 15.020000 51.910000 15.220000 ;
        RECT 51.710000 15.460000 51.910000 15.660000 ;
        RECT 51.710000 15.900000 51.910000 16.100000 ;
        RECT 51.710000 16.340000 51.910000 16.540000 ;
        RECT 51.710000 16.780000 51.910000 16.980000 ;
        RECT 51.710000 17.220000 51.910000 17.420000 ;
        RECT 51.710000 17.660000 51.910000 17.860000 ;
        RECT 51.710000 18.100000 51.910000 18.300000 ;
        RECT 52.120000 15.020000 52.320000 15.220000 ;
        RECT 52.120000 15.460000 52.320000 15.660000 ;
        RECT 52.120000 15.900000 52.320000 16.100000 ;
        RECT 52.120000 16.340000 52.320000 16.540000 ;
        RECT 52.120000 16.780000 52.320000 16.980000 ;
        RECT 52.120000 17.220000 52.320000 17.420000 ;
        RECT 52.120000 17.660000 52.320000 17.860000 ;
        RECT 52.120000 18.100000 52.320000 18.300000 ;
        RECT 52.530000 15.020000 52.730000 15.220000 ;
        RECT 52.530000 15.460000 52.730000 15.660000 ;
        RECT 52.530000 15.900000 52.730000 16.100000 ;
        RECT 52.530000 16.340000 52.730000 16.540000 ;
        RECT 52.530000 16.780000 52.730000 16.980000 ;
        RECT 52.530000 17.220000 52.730000 17.420000 ;
        RECT 52.530000 17.660000 52.730000 17.860000 ;
        RECT 52.530000 18.100000 52.730000 18.300000 ;
        RECT 52.940000 15.020000 53.140000 15.220000 ;
        RECT 52.940000 15.460000 53.140000 15.660000 ;
        RECT 52.940000 15.900000 53.140000 16.100000 ;
        RECT 52.940000 16.340000 53.140000 16.540000 ;
        RECT 52.940000 16.780000 53.140000 16.980000 ;
        RECT 52.940000 17.220000 53.140000 17.420000 ;
        RECT 52.940000 17.660000 53.140000 17.860000 ;
        RECT 52.940000 18.100000 53.140000 18.300000 ;
        RECT 53.345000 15.020000 53.545000 15.220000 ;
        RECT 53.345000 15.460000 53.545000 15.660000 ;
        RECT 53.345000 15.900000 53.545000 16.100000 ;
        RECT 53.345000 16.340000 53.545000 16.540000 ;
        RECT 53.345000 16.780000 53.545000 16.980000 ;
        RECT 53.345000 17.220000 53.545000 17.420000 ;
        RECT 53.345000 17.660000 53.545000 17.860000 ;
        RECT 53.345000 18.100000 53.545000 18.300000 ;
        RECT 53.750000 15.020000 53.950000 15.220000 ;
        RECT 53.750000 15.460000 53.950000 15.660000 ;
        RECT 53.750000 15.900000 53.950000 16.100000 ;
        RECT 53.750000 16.340000 53.950000 16.540000 ;
        RECT 53.750000 16.780000 53.950000 16.980000 ;
        RECT 53.750000 17.220000 53.950000 17.420000 ;
        RECT 53.750000 17.660000 53.950000 17.860000 ;
        RECT 53.750000 18.100000 53.950000 18.300000 ;
        RECT 54.155000 15.020000 54.355000 15.220000 ;
        RECT 54.155000 15.460000 54.355000 15.660000 ;
        RECT 54.155000 15.900000 54.355000 16.100000 ;
        RECT 54.155000 16.340000 54.355000 16.540000 ;
        RECT 54.155000 16.780000 54.355000 16.980000 ;
        RECT 54.155000 17.220000 54.355000 17.420000 ;
        RECT 54.155000 17.660000 54.355000 17.860000 ;
        RECT 54.155000 18.100000 54.355000 18.300000 ;
        RECT 54.560000 15.020000 54.760000 15.220000 ;
        RECT 54.560000 15.460000 54.760000 15.660000 ;
        RECT 54.560000 15.900000 54.760000 16.100000 ;
        RECT 54.560000 16.340000 54.760000 16.540000 ;
        RECT 54.560000 16.780000 54.760000 16.980000 ;
        RECT 54.560000 17.220000 54.760000 17.420000 ;
        RECT 54.560000 17.660000 54.760000 17.860000 ;
        RECT 54.560000 18.100000 54.760000 18.300000 ;
        RECT 54.965000 15.020000 55.165000 15.220000 ;
        RECT 54.965000 15.460000 55.165000 15.660000 ;
        RECT 54.965000 15.900000 55.165000 16.100000 ;
        RECT 54.965000 16.340000 55.165000 16.540000 ;
        RECT 54.965000 16.780000 55.165000 16.980000 ;
        RECT 54.965000 17.220000 55.165000 17.420000 ;
        RECT 54.965000 17.660000 55.165000 17.860000 ;
        RECT 54.965000 18.100000 55.165000 18.300000 ;
        RECT 55.370000 15.020000 55.570000 15.220000 ;
        RECT 55.370000 15.460000 55.570000 15.660000 ;
        RECT 55.370000 15.900000 55.570000 16.100000 ;
        RECT 55.370000 16.340000 55.570000 16.540000 ;
        RECT 55.370000 16.780000 55.570000 16.980000 ;
        RECT 55.370000 17.220000 55.570000 17.420000 ;
        RECT 55.370000 17.660000 55.570000 17.860000 ;
        RECT 55.370000 18.100000 55.570000 18.300000 ;
        RECT 55.775000 15.020000 55.975000 15.220000 ;
        RECT 55.775000 15.460000 55.975000 15.660000 ;
        RECT 55.775000 15.900000 55.975000 16.100000 ;
        RECT 55.775000 16.340000 55.975000 16.540000 ;
        RECT 55.775000 16.780000 55.975000 16.980000 ;
        RECT 55.775000 17.220000 55.975000 17.420000 ;
        RECT 55.775000 17.660000 55.975000 17.860000 ;
        RECT 55.775000 18.100000 55.975000 18.300000 ;
        RECT 56.180000 15.020000 56.380000 15.220000 ;
        RECT 56.180000 15.460000 56.380000 15.660000 ;
        RECT 56.180000 15.900000 56.380000 16.100000 ;
        RECT 56.180000 16.340000 56.380000 16.540000 ;
        RECT 56.180000 16.780000 56.380000 16.980000 ;
        RECT 56.180000 17.220000 56.380000 17.420000 ;
        RECT 56.180000 17.660000 56.380000 17.860000 ;
        RECT 56.180000 18.100000 56.380000 18.300000 ;
        RECT 56.585000 15.020000 56.785000 15.220000 ;
        RECT 56.585000 15.460000 56.785000 15.660000 ;
        RECT 56.585000 15.900000 56.785000 16.100000 ;
        RECT 56.585000 16.340000 56.785000 16.540000 ;
        RECT 56.585000 16.780000 56.785000 16.980000 ;
        RECT 56.585000 17.220000 56.785000 17.420000 ;
        RECT 56.585000 17.660000 56.785000 17.860000 ;
        RECT 56.585000 18.100000 56.785000 18.300000 ;
        RECT 56.990000 15.020000 57.190000 15.220000 ;
        RECT 56.990000 15.460000 57.190000 15.660000 ;
        RECT 56.990000 15.900000 57.190000 16.100000 ;
        RECT 56.990000 16.340000 57.190000 16.540000 ;
        RECT 56.990000 16.780000 57.190000 16.980000 ;
        RECT 56.990000 17.220000 57.190000 17.420000 ;
        RECT 56.990000 17.660000 57.190000 17.860000 ;
        RECT 56.990000 18.100000 57.190000 18.300000 ;
        RECT 57.395000 15.020000 57.595000 15.220000 ;
        RECT 57.395000 15.460000 57.595000 15.660000 ;
        RECT 57.395000 15.900000 57.595000 16.100000 ;
        RECT 57.395000 16.340000 57.595000 16.540000 ;
        RECT 57.395000 16.780000 57.595000 16.980000 ;
        RECT 57.395000 17.220000 57.595000 17.420000 ;
        RECT 57.395000 17.660000 57.595000 17.860000 ;
        RECT 57.395000 18.100000 57.595000 18.300000 ;
        RECT 57.800000 15.020000 58.000000 15.220000 ;
        RECT 57.800000 15.460000 58.000000 15.660000 ;
        RECT 57.800000 15.900000 58.000000 16.100000 ;
        RECT 57.800000 16.340000 58.000000 16.540000 ;
        RECT 57.800000 16.780000 58.000000 16.980000 ;
        RECT 57.800000 17.220000 58.000000 17.420000 ;
        RECT 57.800000 17.660000 58.000000 17.860000 ;
        RECT 57.800000 18.100000 58.000000 18.300000 ;
        RECT 58.205000 15.020000 58.405000 15.220000 ;
        RECT 58.205000 15.460000 58.405000 15.660000 ;
        RECT 58.205000 15.900000 58.405000 16.100000 ;
        RECT 58.205000 16.340000 58.405000 16.540000 ;
        RECT 58.205000 16.780000 58.405000 16.980000 ;
        RECT 58.205000 17.220000 58.405000 17.420000 ;
        RECT 58.205000 17.660000 58.405000 17.860000 ;
        RECT 58.205000 18.100000 58.405000 18.300000 ;
        RECT 58.610000 15.020000 58.810000 15.220000 ;
        RECT 58.610000 15.460000 58.810000 15.660000 ;
        RECT 58.610000 15.900000 58.810000 16.100000 ;
        RECT 58.610000 16.340000 58.810000 16.540000 ;
        RECT 58.610000 16.780000 58.810000 16.980000 ;
        RECT 58.610000 17.220000 58.810000 17.420000 ;
        RECT 58.610000 17.660000 58.810000 17.860000 ;
        RECT 58.610000 18.100000 58.810000 18.300000 ;
        RECT 59.015000 15.020000 59.215000 15.220000 ;
        RECT 59.015000 15.460000 59.215000 15.660000 ;
        RECT 59.015000 15.900000 59.215000 16.100000 ;
        RECT 59.015000 16.340000 59.215000 16.540000 ;
        RECT 59.015000 16.780000 59.215000 16.980000 ;
        RECT 59.015000 17.220000 59.215000 17.420000 ;
        RECT 59.015000 17.660000 59.215000 17.860000 ;
        RECT 59.015000 18.100000 59.215000 18.300000 ;
        RECT 59.420000 15.020000 59.620000 15.220000 ;
        RECT 59.420000 15.460000 59.620000 15.660000 ;
        RECT 59.420000 15.900000 59.620000 16.100000 ;
        RECT 59.420000 16.340000 59.620000 16.540000 ;
        RECT 59.420000 16.780000 59.620000 16.980000 ;
        RECT 59.420000 17.220000 59.620000 17.420000 ;
        RECT 59.420000 17.660000 59.620000 17.860000 ;
        RECT 59.420000 18.100000 59.620000 18.300000 ;
        RECT 59.825000 15.020000 60.025000 15.220000 ;
        RECT 59.825000 15.460000 60.025000 15.660000 ;
        RECT 59.825000 15.900000 60.025000 16.100000 ;
        RECT 59.825000 16.340000 60.025000 16.540000 ;
        RECT 59.825000 16.780000 60.025000 16.980000 ;
        RECT 59.825000 17.220000 60.025000 17.420000 ;
        RECT 59.825000 17.660000 60.025000 17.860000 ;
        RECT 59.825000 18.100000 60.025000 18.300000 ;
        RECT 60.230000 15.020000 60.430000 15.220000 ;
        RECT 60.230000 15.460000 60.430000 15.660000 ;
        RECT 60.230000 15.900000 60.430000 16.100000 ;
        RECT 60.230000 16.340000 60.430000 16.540000 ;
        RECT 60.230000 16.780000 60.430000 16.980000 ;
        RECT 60.230000 17.220000 60.430000 17.420000 ;
        RECT 60.230000 17.660000 60.430000 17.860000 ;
        RECT 60.230000 18.100000 60.430000 18.300000 ;
        RECT 60.635000 15.020000 60.835000 15.220000 ;
        RECT 60.635000 15.460000 60.835000 15.660000 ;
        RECT 60.635000 15.900000 60.835000 16.100000 ;
        RECT 60.635000 16.340000 60.835000 16.540000 ;
        RECT 60.635000 16.780000 60.835000 16.980000 ;
        RECT 60.635000 17.220000 60.835000 17.420000 ;
        RECT 60.635000 17.660000 60.835000 17.860000 ;
        RECT 60.635000 18.100000 60.835000 18.300000 ;
        RECT 61.040000 15.020000 61.240000 15.220000 ;
        RECT 61.040000 15.460000 61.240000 15.660000 ;
        RECT 61.040000 15.900000 61.240000 16.100000 ;
        RECT 61.040000 16.340000 61.240000 16.540000 ;
        RECT 61.040000 16.780000 61.240000 16.980000 ;
        RECT 61.040000 17.220000 61.240000 17.420000 ;
        RECT 61.040000 17.660000 61.240000 17.860000 ;
        RECT 61.040000 18.100000 61.240000 18.300000 ;
        RECT 61.445000 15.020000 61.645000 15.220000 ;
        RECT 61.445000 15.460000 61.645000 15.660000 ;
        RECT 61.445000 15.900000 61.645000 16.100000 ;
        RECT 61.445000 16.340000 61.645000 16.540000 ;
        RECT 61.445000 16.780000 61.645000 16.980000 ;
        RECT 61.445000 17.220000 61.645000 17.420000 ;
        RECT 61.445000 17.660000 61.645000 17.860000 ;
        RECT 61.445000 18.100000 61.645000 18.300000 ;
        RECT 61.850000 15.020000 62.050000 15.220000 ;
        RECT 61.850000 15.460000 62.050000 15.660000 ;
        RECT 61.850000 15.900000 62.050000 16.100000 ;
        RECT 61.850000 16.340000 62.050000 16.540000 ;
        RECT 61.850000 16.780000 62.050000 16.980000 ;
        RECT 61.850000 17.220000 62.050000 17.420000 ;
        RECT 61.850000 17.660000 62.050000 17.860000 ;
        RECT 61.850000 18.100000 62.050000 18.300000 ;
        RECT 62.255000 15.020000 62.455000 15.220000 ;
        RECT 62.255000 15.460000 62.455000 15.660000 ;
        RECT 62.255000 15.900000 62.455000 16.100000 ;
        RECT 62.255000 16.340000 62.455000 16.540000 ;
        RECT 62.255000 16.780000 62.455000 16.980000 ;
        RECT 62.255000 17.220000 62.455000 17.420000 ;
        RECT 62.255000 17.660000 62.455000 17.860000 ;
        RECT 62.255000 18.100000 62.455000 18.300000 ;
        RECT 62.660000 15.020000 62.860000 15.220000 ;
        RECT 62.660000 15.460000 62.860000 15.660000 ;
        RECT 62.660000 15.900000 62.860000 16.100000 ;
        RECT 62.660000 16.340000 62.860000 16.540000 ;
        RECT 62.660000 16.780000 62.860000 16.980000 ;
        RECT 62.660000 17.220000 62.860000 17.420000 ;
        RECT 62.660000 17.660000 62.860000 17.860000 ;
        RECT 62.660000 18.100000 62.860000 18.300000 ;
        RECT 63.065000 15.020000 63.265000 15.220000 ;
        RECT 63.065000 15.460000 63.265000 15.660000 ;
        RECT 63.065000 15.900000 63.265000 16.100000 ;
        RECT 63.065000 16.340000 63.265000 16.540000 ;
        RECT 63.065000 16.780000 63.265000 16.980000 ;
        RECT 63.065000 17.220000 63.265000 17.420000 ;
        RECT 63.065000 17.660000 63.265000 17.860000 ;
        RECT 63.065000 18.100000 63.265000 18.300000 ;
        RECT 63.470000 15.020000 63.670000 15.220000 ;
        RECT 63.470000 15.460000 63.670000 15.660000 ;
        RECT 63.470000 15.900000 63.670000 16.100000 ;
        RECT 63.470000 16.340000 63.670000 16.540000 ;
        RECT 63.470000 16.780000 63.670000 16.980000 ;
        RECT 63.470000 17.220000 63.670000 17.420000 ;
        RECT 63.470000 17.660000 63.670000 17.860000 ;
        RECT 63.470000 18.100000 63.670000 18.300000 ;
        RECT 63.875000 15.020000 64.075000 15.220000 ;
        RECT 63.875000 15.460000 64.075000 15.660000 ;
        RECT 63.875000 15.900000 64.075000 16.100000 ;
        RECT 63.875000 16.340000 64.075000 16.540000 ;
        RECT 63.875000 16.780000 64.075000 16.980000 ;
        RECT 63.875000 17.220000 64.075000 17.420000 ;
        RECT 63.875000 17.660000 64.075000 17.860000 ;
        RECT 63.875000 18.100000 64.075000 18.300000 ;
        RECT 64.280000 15.020000 64.480000 15.220000 ;
        RECT 64.280000 15.460000 64.480000 15.660000 ;
        RECT 64.280000 15.900000 64.480000 16.100000 ;
        RECT 64.280000 16.340000 64.480000 16.540000 ;
        RECT 64.280000 16.780000 64.480000 16.980000 ;
        RECT 64.280000 17.220000 64.480000 17.420000 ;
        RECT 64.280000 17.660000 64.480000 17.860000 ;
        RECT 64.280000 18.100000 64.480000 18.300000 ;
        RECT 64.685000 15.020000 64.885000 15.220000 ;
        RECT 64.685000 15.460000 64.885000 15.660000 ;
        RECT 64.685000 15.900000 64.885000 16.100000 ;
        RECT 64.685000 16.340000 64.885000 16.540000 ;
        RECT 64.685000 16.780000 64.885000 16.980000 ;
        RECT 64.685000 17.220000 64.885000 17.420000 ;
        RECT 64.685000 17.660000 64.885000 17.860000 ;
        RECT 64.685000 18.100000 64.885000 18.300000 ;
        RECT 65.090000 15.020000 65.290000 15.220000 ;
        RECT 65.090000 15.460000 65.290000 15.660000 ;
        RECT 65.090000 15.900000 65.290000 16.100000 ;
        RECT 65.090000 16.340000 65.290000 16.540000 ;
        RECT 65.090000 16.780000 65.290000 16.980000 ;
        RECT 65.090000 17.220000 65.290000 17.420000 ;
        RECT 65.090000 17.660000 65.290000 17.860000 ;
        RECT 65.090000 18.100000 65.290000 18.300000 ;
        RECT 65.495000 15.020000 65.695000 15.220000 ;
        RECT 65.495000 15.460000 65.695000 15.660000 ;
        RECT 65.495000 15.900000 65.695000 16.100000 ;
        RECT 65.495000 16.340000 65.695000 16.540000 ;
        RECT 65.495000 16.780000 65.695000 16.980000 ;
        RECT 65.495000 17.220000 65.695000 17.420000 ;
        RECT 65.495000 17.660000 65.695000 17.860000 ;
        RECT 65.495000 18.100000 65.695000 18.300000 ;
        RECT 65.900000 15.020000 66.100000 15.220000 ;
        RECT 65.900000 15.460000 66.100000 15.660000 ;
        RECT 65.900000 15.900000 66.100000 16.100000 ;
        RECT 65.900000 16.340000 66.100000 16.540000 ;
        RECT 65.900000 16.780000 66.100000 16.980000 ;
        RECT 65.900000 17.220000 66.100000 17.420000 ;
        RECT 65.900000 17.660000 66.100000 17.860000 ;
        RECT 65.900000 18.100000 66.100000 18.300000 ;
        RECT 66.305000 15.020000 66.505000 15.220000 ;
        RECT 66.305000 15.460000 66.505000 15.660000 ;
        RECT 66.305000 15.900000 66.505000 16.100000 ;
        RECT 66.305000 16.340000 66.505000 16.540000 ;
        RECT 66.305000 16.780000 66.505000 16.980000 ;
        RECT 66.305000 17.220000 66.505000 17.420000 ;
        RECT 66.305000 17.660000 66.505000 17.860000 ;
        RECT 66.305000 18.100000 66.505000 18.300000 ;
        RECT 66.710000 15.020000 66.910000 15.220000 ;
        RECT 66.710000 15.460000 66.910000 15.660000 ;
        RECT 66.710000 15.900000 66.910000 16.100000 ;
        RECT 66.710000 16.340000 66.910000 16.540000 ;
        RECT 66.710000 16.780000 66.910000 16.980000 ;
        RECT 66.710000 17.220000 66.910000 17.420000 ;
        RECT 66.710000 17.660000 66.910000 17.860000 ;
        RECT 66.710000 18.100000 66.910000 18.300000 ;
        RECT 67.115000 15.020000 67.315000 15.220000 ;
        RECT 67.115000 15.460000 67.315000 15.660000 ;
        RECT 67.115000 15.900000 67.315000 16.100000 ;
        RECT 67.115000 16.340000 67.315000 16.540000 ;
        RECT 67.115000 16.780000 67.315000 16.980000 ;
        RECT 67.115000 17.220000 67.315000 17.420000 ;
        RECT 67.115000 17.660000 67.315000 17.860000 ;
        RECT 67.115000 18.100000 67.315000 18.300000 ;
        RECT 67.520000 15.020000 67.720000 15.220000 ;
        RECT 67.520000 15.460000 67.720000 15.660000 ;
        RECT 67.520000 15.900000 67.720000 16.100000 ;
        RECT 67.520000 16.340000 67.720000 16.540000 ;
        RECT 67.520000 16.780000 67.720000 16.980000 ;
        RECT 67.520000 17.220000 67.720000 17.420000 ;
        RECT 67.520000 17.660000 67.720000 17.860000 ;
        RECT 67.520000 18.100000 67.720000 18.300000 ;
        RECT 67.925000 15.020000 68.125000 15.220000 ;
        RECT 67.925000 15.460000 68.125000 15.660000 ;
        RECT 67.925000 15.900000 68.125000 16.100000 ;
        RECT 67.925000 16.340000 68.125000 16.540000 ;
        RECT 67.925000 16.780000 68.125000 16.980000 ;
        RECT 67.925000 17.220000 68.125000 17.420000 ;
        RECT 67.925000 17.660000 68.125000 17.860000 ;
        RECT 67.925000 18.100000 68.125000 18.300000 ;
        RECT 68.330000 15.020000 68.530000 15.220000 ;
        RECT 68.330000 15.460000 68.530000 15.660000 ;
        RECT 68.330000 15.900000 68.530000 16.100000 ;
        RECT 68.330000 16.340000 68.530000 16.540000 ;
        RECT 68.330000 16.780000 68.530000 16.980000 ;
        RECT 68.330000 17.220000 68.530000 17.420000 ;
        RECT 68.330000 17.660000 68.530000 17.860000 ;
        RECT 68.330000 18.100000 68.530000 18.300000 ;
        RECT 68.735000 15.020000 68.935000 15.220000 ;
        RECT 68.735000 15.460000 68.935000 15.660000 ;
        RECT 68.735000 15.900000 68.935000 16.100000 ;
        RECT 68.735000 16.340000 68.935000 16.540000 ;
        RECT 68.735000 16.780000 68.935000 16.980000 ;
        RECT 68.735000 17.220000 68.935000 17.420000 ;
        RECT 68.735000 17.660000 68.935000 17.860000 ;
        RECT 68.735000 18.100000 68.935000 18.300000 ;
        RECT 69.140000 15.020000 69.340000 15.220000 ;
        RECT 69.140000 15.460000 69.340000 15.660000 ;
        RECT 69.140000 15.900000 69.340000 16.100000 ;
        RECT 69.140000 16.340000 69.340000 16.540000 ;
        RECT 69.140000 16.780000 69.340000 16.980000 ;
        RECT 69.140000 17.220000 69.340000 17.420000 ;
        RECT 69.140000 17.660000 69.340000 17.860000 ;
        RECT 69.140000 18.100000 69.340000 18.300000 ;
        RECT 69.545000 15.020000 69.745000 15.220000 ;
        RECT 69.545000 15.460000 69.745000 15.660000 ;
        RECT 69.545000 15.900000 69.745000 16.100000 ;
        RECT 69.545000 16.340000 69.745000 16.540000 ;
        RECT 69.545000 16.780000 69.745000 16.980000 ;
        RECT 69.545000 17.220000 69.745000 17.420000 ;
        RECT 69.545000 17.660000 69.745000 17.860000 ;
        RECT 69.545000 18.100000 69.745000 18.300000 ;
        RECT 69.950000 15.020000 70.150000 15.220000 ;
        RECT 69.950000 15.460000 70.150000 15.660000 ;
        RECT 69.950000 15.900000 70.150000 16.100000 ;
        RECT 69.950000 16.340000 70.150000 16.540000 ;
        RECT 69.950000 16.780000 70.150000 16.980000 ;
        RECT 69.950000 17.220000 70.150000 17.420000 ;
        RECT 69.950000 17.660000 70.150000 17.860000 ;
        RECT 69.950000 18.100000 70.150000 18.300000 ;
        RECT 70.355000 15.020000 70.555000 15.220000 ;
        RECT 70.355000 15.460000 70.555000 15.660000 ;
        RECT 70.355000 15.900000 70.555000 16.100000 ;
        RECT 70.355000 16.340000 70.555000 16.540000 ;
        RECT 70.355000 16.780000 70.555000 16.980000 ;
        RECT 70.355000 17.220000 70.555000 17.420000 ;
        RECT 70.355000 17.660000 70.555000 17.860000 ;
        RECT 70.355000 18.100000 70.555000 18.300000 ;
        RECT 70.760000 15.020000 70.960000 15.220000 ;
        RECT 70.760000 15.460000 70.960000 15.660000 ;
        RECT 70.760000 15.900000 70.960000 16.100000 ;
        RECT 70.760000 16.340000 70.960000 16.540000 ;
        RECT 70.760000 16.780000 70.960000 16.980000 ;
        RECT 70.760000 17.220000 70.960000 17.420000 ;
        RECT 70.760000 17.660000 70.960000 17.860000 ;
        RECT 70.760000 18.100000 70.960000 18.300000 ;
        RECT 71.165000 15.020000 71.365000 15.220000 ;
        RECT 71.165000 15.460000 71.365000 15.660000 ;
        RECT 71.165000 15.900000 71.365000 16.100000 ;
        RECT 71.165000 16.340000 71.365000 16.540000 ;
        RECT 71.165000 16.780000 71.365000 16.980000 ;
        RECT 71.165000 17.220000 71.365000 17.420000 ;
        RECT 71.165000 17.660000 71.365000 17.860000 ;
        RECT 71.165000 18.100000 71.365000 18.300000 ;
        RECT 71.570000 15.020000 71.770000 15.220000 ;
        RECT 71.570000 15.460000 71.770000 15.660000 ;
        RECT 71.570000 15.900000 71.770000 16.100000 ;
        RECT 71.570000 16.340000 71.770000 16.540000 ;
        RECT 71.570000 16.780000 71.770000 16.980000 ;
        RECT 71.570000 17.220000 71.770000 17.420000 ;
        RECT 71.570000 17.660000 71.770000 17.860000 ;
        RECT 71.570000 18.100000 71.770000 18.300000 ;
        RECT 71.975000 15.020000 72.175000 15.220000 ;
        RECT 71.975000 15.460000 72.175000 15.660000 ;
        RECT 71.975000 15.900000 72.175000 16.100000 ;
        RECT 71.975000 16.340000 72.175000 16.540000 ;
        RECT 71.975000 16.780000 72.175000 16.980000 ;
        RECT 71.975000 17.220000 72.175000 17.420000 ;
        RECT 71.975000 17.660000 72.175000 17.860000 ;
        RECT 71.975000 18.100000 72.175000 18.300000 ;
        RECT 72.380000 15.020000 72.580000 15.220000 ;
        RECT 72.380000 15.460000 72.580000 15.660000 ;
        RECT 72.380000 15.900000 72.580000 16.100000 ;
        RECT 72.380000 16.340000 72.580000 16.540000 ;
        RECT 72.380000 16.780000 72.580000 16.980000 ;
        RECT 72.380000 17.220000 72.580000 17.420000 ;
        RECT 72.380000 17.660000 72.580000 17.860000 ;
        RECT 72.380000 18.100000 72.580000 18.300000 ;
        RECT 72.785000 15.020000 72.985000 15.220000 ;
        RECT 72.785000 15.460000 72.985000 15.660000 ;
        RECT 72.785000 15.900000 72.985000 16.100000 ;
        RECT 72.785000 16.340000 72.985000 16.540000 ;
        RECT 72.785000 16.780000 72.985000 16.980000 ;
        RECT 72.785000 17.220000 72.985000 17.420000 ;
        RECT 72.785000 17.660000 72.985000 17.860000 ;
        RECT 72.785000 18.100000 72.985000 18.300000 ;
        RECT 73.190000 15.020000 73.390000 15.220000 ;
        RECT 73.190000 15.460000 73.390000 15.660000 ;
        RECT 73.190000 15.900000 73.390000 16.100000 ;
        RECT 73.190000 16.340000 73.390000 16.540000 ;
        RECT 73.190000 16.780000 73.390000 16.980000 ;
        RECT 73.190000 17.220000 73.390000 17.420000 ;
        RECT 73.190000 17.660000 73.390000 17.860000 ;
        RECT 73.190000 18.100000 73.390000 18.300000 ;
        RECT 73.595000 15.020000 73.795000 15.220000 ;
        RECT 73.595000 15.460000 73.795000 15.660000 ;
        RECT 73.595000 15.900000 73.795000 16.100000 ;
        RECT 73.595000 16.340000 73.795000 16.540000 ;
        RECT 73.595000 16.780000 73.795000 16.980000 ;
        RECT 73.595000 17.220000 73.795000 17.420000 ;
        RECT 73.595000 17.660000 73.795000 17.860000 ;
        RECT 73.595000 18.100000 73.795000 18.300000 ;
        RECT 74.000000 15.020000 74.200000 15.220000 ;
        RECT 74.000000 15.460000 74.200000 15.660000 ;
        RECT 74.000000 15.900000 74.200000 16.100000 ;
        RECT 74.000000 16.340000 74.200000 16.540000 ;
        RECT 74.000000 16.780000 74.200000 16.980000 ;
        RECT 74.000000 17.220000 74.200000 17.420000 ;
        RECT 74.000000 17.660000 74.200000 17.860000 ;
        RECT 74.000000 18.100000 74.200000 18.300000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 75.000000  14.540000 ;
      RECT  0.000000 18.780000 75.000000 200.000000 ;
      RECT 24.795000 14.540000 49.990000  18.780000 ;
      RECT 74.690000 14.540000 75.000000  18.780000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000  13.935000  1.670000  14.535000 ;
      RECT  0.000000  18.785000  1.670000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.670000   0.000000 73.330000  14.535000 ;
      RECT  1.670000  18.785000 73.330000  95.400000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT 24.770000  14.535000 50.015000  18.785000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  13.935000 75.000000  14.535000 ;
      RECT 73.330000  18.785000 75.000000  19.385000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
    LAYER met5 ;
      RECT 0.000000   0.000000 75.000000   1.335000 ;
      RECT 0.000000  95.785000 75.000000 174.985000 ;
      RECT 1.765000  14.235000 73.235000  19.085000 ;
      RECT 2.070000   1.335000 72.930000  14.235000 ;
      RECT 2.070000  19.085000 72.930000  95.785000 ;
      RECT 2.070000 174.985000 72.930000 200.000000 ;
  END
END sky130_fd_io__overlay_vdda_hvc


MACRO sky130_fd_io__top_power_lvc_wpad
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN P_PAD
    ANTENNAPARTIALMETALSIDEAREA  243.2170 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 31.695000 162.765000 52.340000 167.120000 ;
    END
  END P_PAD
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 17.630000 5.115000 53.535000 9.540000 ;
        RECT 17.635000 5.110000 53.535000 5.115000 ;
        RECT 17.705000 5.040000 53.535000 5.110000 ;
        RECT 17.775000 4.970000 53.535000 5.040000 ;
        RECT 17.845000 4.900000 53.535000 4.970000 ;
        RECT 17.915000 4.830000 53.535000 4.900000 ;
        RECT 17.985000 4.760000 53.535000 4.830000 ;
        RECT 18.055000 4.690000 53.535000 4.760000 ;
        RECT 18.125000 4.620000 53.535000 4.690000 ;
        RECT 18.195000 4.550000 53.535000 4.620000 ;
        RECT 18.265000 4.480000 53.535000 4.550000 ;
        RECT 18.335000 4.410000 53.535000 4.480000 ;
        RECT 18.405000 4.340000 53.535000 4.410000 ;
        RECT 18.475000 4.270000 53.535000 4.340000 ;
        RECT 18.545000 4.200000 53.535000 4.270000 ;
        RECT 18.615000 4.130000 53.535000 4.200000 ;
        RECT 18.685000 4.060000 53.535000 4.130000 ;
        RECT 18.755000 3.990000 53.535000 4.060000 ;
        RECT 18.825000 3.920000 53.535000 3.990000 ;
        RECT 18.895000 3.850000 53.535000 3.920000 ;
        RECT 18.965000 3.780000 53.535000 3.850000 ;
        RECT 19.035000 3.710000 53.535000 3.780000 ;
        RECT 19.105000 3.640000 53.535000 3.710000 ;
        RECT 19.175000 3.570000 53.535000 3.640000 ;
        RECT 19.245000 3.500000 53.535000 3.570000 ;
        RECT 19.315000 3.430000 53.535000 3.500000 ;
        RECT 19.385000 3.360000 53.535000 3.430000 ;
        RECT 19.455000 3.290000 53.535000 3.360000 ;
        RECT 19.525000 3.220000 53.535000 3.290000 ;
        RECT 19.595000 3.150000 53.535000 3.220000 ;
        RECT 19.665000 3.080000 53.535000 3.150000 ;
        RECT 19.735000 3.010000 53.535000 3.080000 ;
        RECT 19.805000 2.940000 53.535000 3.010000 ;
        RECT 19.875000 2.870000 53.535000 2.940000 ;
        RECT 19.945000 2.800000 53.535000 2.870000 ;
        RECT 20.015000 2.730000 53.535000 2.800000 ;
        RECT 20.085000 2.660000 53.535000 2.730000 ;
        RECT 20.155000 2.590000 53.535000 2.660000 ;
        RECT 20.225000 2.520000 53.535000 2.590000 ;
        RECT 20.295000 2.450000 53.535000 2.520000 ;
        RECT 20.365000 2.380000 53.535000 2.450000 ;
        RECT 20.435000 2.310000 53.535000 2.380000 ;
        RECT 20.505000 2.240000 53.535000 2.310000 ;
        RECT 20.575000 2.170000 53.535000 2.240000 ;
        RECT 20.645000 2.100000 53.535000 2.170000 ;
        RECT 20.715000 2.030000 53.535000 2.100000 ;
        RECT 20.785000 1.960000 53.535000 2.030000 ;
        RECT 20.855000 1.890000 53.535000 1.960000 ;
        RECT 20.925000 0.000000 53.535000 1.820000 ;
        RECT 20.925000 1.820000 53.535000 1.890000 ;
    END
  END BDY2_B2B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 15.605000  94.310000 23.935000  94.460000 ;
        RECT 15.605000  94.460000 23.785000  94.610000 ;
        RECT 15.605000  94.610000 23.635000  94.760000 ;
        RECT 15.605000  94.760000 23.485000  94.910000 ;
        RECT 15.605000  94.910000 23.335000  95.060000 ;
        RECT 15.605000  95.060000 23.185000  95.210000 ;
        RECT 15.605000  95.210000 23.035000  95.360000 ;
        RECT 15.605000  95.360000 22.885000  95.510000 ;
        RECT 15.605000  95.510000 22.735000  95.660000 ;
        RECT 15.605000  95.660000 22.585000  95.810000 ;
        RECT 15.605000  95.810000 22.435000  95.960000 ;
        RECT 15.605000  95.960000 22.285000  96.110000 ;
        RECT 15.605000  96.110000 22.135000  96.260000 ;
        RECT 15.605000  96.260000 21.985000  96.410000 ;
        RECT 15.605000  96.410000 21.835000  96.560000 ;
        RECT 15.605000  96.560000 21.685000  96.710000 ;
        RECT 15.605000  96.710000 21.605000  96.790000 ;
        RECT 15.605000  96.790000 21.605000 167.100000 ;
        RECT 15.605000 167.100000 21.605000 167.250000 ;
        RECT 15.605000 167.250000 21.755000 167.400000 ;
        RECT 15.605000 167.400000 21.905000 167.550000 ;
        RECT 15.605000 167.550000 22.055000 167.700000 ;
        RECT 15.605000 167.700000 22.205000 167.850000 ;
        RECT 15.605000 167.850000 22.355000 168.000000 ;
        RECT 15.605000 168.000000 22.505000 168.150000 ;
        RECT 15.605000 168.150000 22.655000 168.300000 ;
        RECT 15.605000 168.300000 22.805000 168.450000 ;
        RECT 15.605000 168.450000 22.955000 168.600000 ;
        RECT 15.605000 168.600000 23.105000 168.750000 ;
        RECT 15.605000 168.750000 23.255000 168.900000 ;
        RECT 15.605000 168.900000 23.405000 169.050000 ;
        RECT 15.605000 169.050000 23.555000 169.200000 ;
        RECT 15.605000 169.200000 23.705000 169.350000 ;
        RECT 15.605000 169.350000 23.855000 169.500000 ;
        RECT 15.605000 169.500000 24.005000 169.650000 ;
        RECT 15.605000 169.650000 24.155000 169.800000 ;
        RECT 15.605000 169.800000 24.305000 169.950000 ;
        RECT 15.605000 169.950000 24.455000 170.100000 ;
        RECT 15.605000 170.100000 24.605000 170.250000 ;
        RECT 15.605000 170.250000 24.755000 170.400000 ;
        RECT 15.605000 170.400000 24.905000 170.550000 ;
        RECT 15.605000 170.550000 25.055000 170.610000 ;
        RECT 15.605000 170.610000 25.115000 189.515000 ;
        RECT 15.715000  94.200000 24.085000  94.310000 ;
        RECT 15.865000  94.050000 24.195000  94.200000 ;
        RECT 16.015000  93.900000 24.345000  94.050000 ;
        RECT 16.165000  93.750000 24.495000  93.900000 ;
        RECT 16.315000  93.600000 24.645000  93.750000 ;
        RECT 16.465000  93.450000 24.795000  93.600000 ;
        RECT 16.615000  93.300000 24.945000  93.450000 ;
        RECT 16.765000  93.150000 25.095000  93.300000 ;
        RECT 16.915000  93.000000 25.245000  93.150000 ;
        RECT 17.065000  92.850000 25.395000  93.000000 ;
        RECT 17.215000  92.700000 25.545000  92.850000 ;
        RECT 17.365000  92.550000 25.695000  92.700000 ;
        RECT 17.515000  92.400000 25.845000  92.550000 ;
        RECT 17.665000  92.250000 25.995000  92.400000 ;
        RECT 17.815000  92.100000 26.145000  92.250000 ;
        RECT 17.965000  91.950000 26.295000  92.100000 ;
        RECT 18.115000  91.800000 26.445000  91.950000 ;
        RECT 18.265000  91.650000 26.595000  91.800000 ;
        RECT 18.415000  91.500000 26.745000  91.650000 ;
        RECT 18.565000  91.350000 26.895000  91.500000 ;
        RECT 18.715000  91.200000 27.045000  91.350000 ;
        RECT 18.865000  91.050000 27.195000  91.200000 ;
        RECT 19.015000  90.900000 27.345000  91.050000 ;
        RECT 19.165000  90.750000 27.495000  90.900000 ;
        RECT 19.315000  90.600000 27.645000  90.750000 ;
        RECT 19.465000  90.450000 27.795000  90.600000 ;
        RECT 19.615000  90.300000 27.945000  90.450000 ;
        RECT 19.765000  90.150000 28.095000  90.300000 ;
        RECT 19.915000  90.000000 28.245000  90.150000 ;
        RECT 20.065000  89.850000 28.395000  90.000000 ;
        RECT 20.215000  89.700000 28.545000  89.850000 ;
        RECT 20.365000  89.550000 28.695000  89.700000 ;
        RECT 20.515000  89.400000 28.845000  89.550000 ;
        RECT 20.665000  89.250000 28.995000  89.400000 ;
        RECT 20.815000  89.100000 29.145000  89.250000 ;
        RECT 20.965000  88.950000 29.295000  89.100000 ;
        RECT 21.115000  88.800000 29.445000  88.950000 ;
        RECT 21.265000  88.650000 29.595000  88.800000 ;
        RECT 21.415000  88.500000 29.745000  88.650000 ;
        RECT 21.565000  88.350000 29.895000  88.500000 ;
        RECT 21.715000  88.200000 30.045000  88.350000 ;
        RECT 21.865000  88.050000 30.195000  88.200000 ;
        RECT 22.015000  87.900000 30.345000  88.050000 ;
        RECT 22.165000  87.750000 30.495000  87.900000 ;
        RECT 22.315000  87.600000 30.645000  87.750000 ;
        RECT 22.465000  87.450000 30.795000  87.600000 ;
        RECT 22.615000  87.300000 30.945000  87.450000 ;
        RECT 22.765000  87.150000 31.095000  87.300000 ;
        RECT 22.915000  87.000000 31.245000  87.150000 ;
        RECT 23.065000  86.850000 31.395000  87.000000 ;
        RECT 23.215000  86.700000 31.545000  86.850000 ;
        RECT 23.365000  86.550000 31.695000  86.700000 ;
        RECT 23.515000  86.400000 31.845000  86.550000 ;
        RECT 23.665000  86.250000 31.995000  86.400000 ;
        RECT 23.670000  86.245000 32.145000  86.250000 ;
        RECT 23.760000  86.155000 32.145000  86.245000 ;
        RECT 23.850000  84.650000 32.165000  84.670000 ;
        RECT 23.850000  84.670000 32.145000  84.690000 ;
        RECT 23.850000  84.690000 32.145000  86.065000 ;
        RECT 23.850000  86.065000 32.145000  86.155000 ;
        RECT 23.920000  84.580000 32.185000  84.650000 ;
        RECT 24.070000  84.430000 32.255000  84.580000 ;
        RECT 24.220000  84.280000 32.405000  84.430000 ;
        RECT 24.370000  84.130000 32.555000  84.280000 ;
        RECT 24.520000  83.980000 32.705000  84.130000 ;
        RECT 24.650000  83.850000 48.870000  83.980000 ;
        RECT 24.800000  83.700000 48.870000  83.850000 ;
        RECT 24.950000  83.550000 48.870000  83.700000 ;
        RECT 25.100000  83.400000 48.870000  83.550000 ;
        RECT 25.250000  83.250000 48.870000  83.400000 ;
        RECT 25.400000  83.100000 48.870000  83.250000 ;
        RECT 25.550000  82.950000 48.870000  83.100000 ;
        RECT 25.700000  82.800000 48.870000  82.950000 ;
        RECT 25.850000  82.650000 48.870000  82.800000 ;
        RECT 26.000000   0.000000 36.880000  71.105000 ;
        RECT 26.000000  71.105000 36.880000  71.255000 ;
        RECT 26.000000  71.255000 37.030000  71.405000 ;
        RECT 26.000000  71.405000 37.180000  71.555000 ;
        RECT 26.000000  71.555000 37.330000  71.705000 ;
        RECT 26.000000  71.705000 37.480000  71.855000 ;
        RECT 26.000000  71.855000 37.630000  72.005000 ;
        RECT 26.000000  72.005000 37.780000  72.155000 ;
        RECT 26.000000  72.155000 37.930000  72.305000 ;
        RECT 26.000000  72.305000 38.080000  72.455000 ;
        RECT 26.000000  72.455000 38.230000  72.605000 ;
        RECT 26.000000  72.605000 38.380000  72.755000 ;
        RECT 26.000000  72.755000 38.530000  72.905000 ;
        RECT 26.000000  72.905000 38.680000  73.055000 ;
        RECT 26.000000  73.055000 38.830000  73.205000 ;
        RECT 26.000000  73.205000 38.980000  73.355000 ;
        RECT 26.000000  73.355000 39.130000  73.505000 ;
        RECT 26.000000  73.505000 39.280000  73.655000 ;
        RECT 26.000000  73.655000 39.430000  73.805000 ;
        RECT 26.000000  73.805000 39.580000  73.955000 ;
        RECT 26.000000  73.955000 39.730000  74.105000 ;
        RECT 26.000000  74.105000 39.880000  74.255000 ;
        RECT 26.000000  74.255000 40.030000  74.405000 ;
        RECT 26.000000  74.405000 40.180000  74.555000 ;
        RECT 26.000000  74.555000 40.330000  74.705000 ;
        RECT 26.000000  74.705000 40.480000  74.740000 ;
        RECT 26.000000  74.740000 46.795000  74.890000 ;
        RECT 26.000000  74.890000 46.945000  75.040000 ;
        RECT 26.000000  75.040000 47.095000  75.190000 ;
        RECT 26.000000  75.190000 47.245000  75.340000 ;
        RECT 26.000000  75.340000 47.395000  75.490000 ;
        RECT 26.000000  75.490000 47.545000  75.640000 ;
        RECT 26.000000  75.640000 47.695000  75.790000 ;
        RECT 26.000000  75.790000 47.845000  75.940000 ;
        RECT 26.000000  75.940000 47.995000  76.090000 ;
        RECT 26.000000  76.090000 48.145000  76.240000 ;
        RECT 26.000000  76.240000 48.295000  76.390000 ;
        RECT 26.000000  76.390000 48.445000  76.540000 ;
        RECT 26.000000  76.540000 48.595000  76.690000 ;
        RECT 26.000000  76.690000 48.745000  76.815000 ;
        RECT 26.000000  76.815000 48.870000  82.500000 ;
        RECT 26.000000  82.500000 48.870000  82.650000 ;
        RECT 26.035000  94.500000 32.035000 162.570000 ;
        RECT 26.035000 162.570000 32.035000 162.720000 ;
        RECT 26.035000 162.720000 32.185000 162.870000 ;
        RECT 26.035000 162.870000 32.335000 163.020000 ;
        RECT 26.035000 163.020000 32.485000 163.170000 ;
        RECT 26.035000 163.170000 32.635000 163.320000 ;
        RECT 26.035000 163.320000 32.785000 163.470000 ;
        RECT 26.035000 163.470000 32.935000 163.620000 ;
        RECT 26.035000 163.620000 33.085000 163.770000 ;
        RECT 26.035000 163.770000 33.235000 163.920000 ;
        RECT 26.035000 163.920000 33.385000 164.070000 ;
        RECT 26.035000 164.070000 33.535000 164.220000 ;
        RECT 26.035000 164.220000 33.685000 164.370000 ;
        RECT 26.035000 164.370000 33.835000 164.520000 ;
        RECT 26.035000 164.520000 33.985000 164.670000 ;
        RECT 26.035000 164.670000 34.135000 164.820000 ;
        RECT 26.035000 164.820000 34.285000 164.970000 ;
        RECT 26.035000 164.970000 34.435000 165.120000 ;
        RECT 26.035000 165.120000 34.585000 165.270000 ;
        RECT 26.035000 165.270000 34.735000 165.420000 ;
        RECT 26.035000 165.420000 34.885000 165.570000 ;
        RECT 26.035000 165.570000 35.035000 165.720000 ;
        RECT 26.035000 165.720000 35.185000 165.870000 ;
        RECT 26.035000 165.870000 35.335000 166.020000 ;
        RECT 26.035000 166.020000 35.485000 166.170000 ;
        RECT 26.035000 166.170000 35.635000 166.320000 ;
        RECT 26.035000 166.320000 35.785000 166.470000 ;
        RECT 26.035000 166.470000 35.935000 166.620000 ;
        RECT 26.035000 166.620000 36.085000 166.770000 ;
        RECT 26.035000 166.770000 36.235000 166.920000 ;
        RECT 26.035000 166.920000 36.385000 167.070000 ;
        RECT 26.035000 167.070000 36.535000 167.220000 ;
        RECT 26.035000 167.220000 36.685000 167.370000 ;
        RECT 26.035000 167.370000 36.835000 167.460000 ;
        RECT 26.035000 167.460000 36.925000 189.515000 ;
        RECT 26.095000  94.440000 32.035000  94.500000 ;
        RECT 26.245000  94.290000 32.035000  94.440000 ;
        RECT 26.395000  94.140000 32.035000  94.290000 ;
        RECT 26.545000  93.990000 32.035000  94.140000 ;
        RECT 26.695000  93.840000 32.035000  93.990000 ;
        RECT 26.845000  93.690000 32.035000  93.840000 ;
        RECT 26.995000  93.540000 32.035000  93.690000 ;
        RECT 27.145000  93.390000 32.035000  93.540000 ;
        RECT 27.160000  93.375000 32.035000  93.390000 ;
        RECT 27.310000  93.225000 32.050000  93.375000 ;
        RECT 27.460000  93.075000 32.200000  93.225000 ;
        RECT 27.610000  92.925000 32.350000  93.075000 ;
        RECT 27.760000  92.775000 32.500000  92.925000 ;
        RECT 27.910000  92.625000 32.650000  92.775000 ;
        RECT 28.060000  92.475000 32.800000  92.625000 ;
        RECT 28.210000  92.325000 32.950000  92.475000 ;
        RECT 28.360000  92.175000 33.100000  92.325000 ;
        RECT 28.510000  92.025000 33.250000  92.175000 ;
        RECT 28.660000  91.875000 33.400000  92.025000 ;
        RECT 28.810000  91.725000 33.550000  91.875000 ;
        RECT 28.960000  91.575000 33.700000  91.725000 ;
        RECT 29.110000  91.425000 33.850000  91.575000 ;
        RECT 29.260000  91.275000 34.000000  91.425000 ;
        RECT 29.410000  91.125000 34.150000  91.275000 ;
        RECT 29.560000  90.975000 34.300000  91.125000 ;
        RECT 29.710000  90.825000 34.450000  90.975000 ;
        RECT 29.860000  90.675000 34.600000  90.825000 ;
        RECT 30.010000  90.525000 34.750000  90.675000 ;
        RECT 30.160000  90.375000 34.900000  90.525000 ;
        RECT 30.175000  90.360000 42.385000  90.375000 ;
        RECT 30.325000  90.210000 42.235000  90.360000 ;
        RECT 30.475000  90.060000 42.085000  90.210000 ;
        RECT 30.625000  89.910000 41.935000  90.060000 ;
        RECT 30.775000  89.760000 41.785000  89.910000 ;
        RECT 30.925000  89.610000 41.635000  89.760000 ;
        RECT 31.075000  89.460000 41.485000  89.610000 ;
        RECT 31.225000  89.310000 41.335000  89.460000 ;
        RECT 31.375000  89.160000 41.185000  89.310000 ;
        RECT 31.525000  89.010000 41.035000  89.160000 ;
        RECT 31.675000  88.860000 40.885000  89.010000 ;
        RECT 31.825000  88.710000 40.735000  88.860000 ;
        RECT 31.975000  88.560000 40.585000  88.710000 ;
        RECT 32.125000  88.410000 40.435000  88.560000 ;
        RECT 32.275000  88.260000 40.285000  88.410000 ;
        RECT 32.425000  88.110000 40.135000  88.260000 ;
        RECT 32.575000  87.960000 39.985000  88.110000 ;
        RECT 32.725000  87.810000 39.835000  87.960000 ;
        RECT 32.875000  87.660000 39.685000  87.810000 ;
        RECT 33.025000  87.510000 39.535000  87.660000 ;
        RECT 33.175000  87.360000 39.385000  87.510000 ;
        RECT 33.305000  87.230000 39.385000  87.360000 ;
        RECT 33.455000  87.080000 39.385000  87.230000 ;
        RECT 33.605000  86.930000 39.385000  87.080000 ;
        RECT 33.755000  86.780000 39.385000  86.930000 ;
        RECT 33.905000  86.630000 39.385000  86.780000 ;
        RECT 33.945000  83.980000 39.945000  84.130000 ;
        RECT 34.055000  86.480000 39.385000  86.630000 ;
        RECT 34.095000  84.130000 39.795000  84.280000 ;
        RECT 34.205000  86.330000 39.385000  86.480000 ;
        RECT 34.245000  84.280000 39.645000  84.430000 ;
        RECT 34.355000  86.180000 39.385000  86.330000 ;
        RECT 34.395000  84.430000 39.495000  84.580000 ;
        RECT 34.505000  84.580000 39.385000  84.690000 ;
        RECT 34.505000  84.690000 39.385000  86.030000 ;
        RECT 34.505000  86.030000 39.385000  86.180000 ;
        RECT 37.945000  90.375000 42.400000  90.525000 ;
        RECT 37.945000 169.025000 48.835000 189.515000 ;
        RECT 38.035000 168.935000 48.835000 169.025000 ;
        RECT 38.095000  90.525000 42.550000  90.675000 ;
        RECT 38.185000 168.785000 48.835000 168.935000 ;
        RECT 38.245000  90.675000 42.700000  90.825000 ;
        RECT 38.335000 168.635000 48.835000 168.785000 ;
        RECT 38.395000  90.825000 42.850000  90.975000 ;
        RECT 38.485000 168.485000 48.835000 168.635000 ;
        RECT 38.545000  90.975000 43.000000  91.125000 ;
        RECT 38.635000 168.335000 48.835000 168.485000 ;
        RECT 38.695000  91.125000 43.150000  91.275000 ;
        RECT 38.785000 168.185000 48.835000 168.335000 ;
        RECT 38.845000  91.275000 43.300000  91.425000 ;
        RECT 38.935000 168.035000 48.835000 168.185000 ;
        RECT 38.995000  91.425000 43.450000  91.575000 ;
        RECT 39.085000 167.885000 48.835000 168.035000 ;
        RECT 39.145000  91.575000 43.600000  91.725000 ;
        RECT 39.235000 167.735000 48.835000 167.885000 ;
        RECT 39.295000  91.725000 43.750000  91.875000 ;
        RECT 39.385000 167.585000 48.835000 167.735000 ;
        RECT 39.445000  91.875000 43.900000  92.025000 ;
        RECT 39.535000 167.435000 48.835000 167.585000 ;
        RECT 39.595000  92.025000 44.050000  92.175000 ;
        RECT 39.685000 167.285000 48.835000 167.435000 ;
        RECT 39.745000  92.175000 44.200000  92.325000 ;
        RECT 39.835000 167.135000 48.835000 167.285000 ;
        RECT 39.895000  92.325000 44.350000  92.475000 ;
        RECT 39.985000 166.985000 48.835000 167.135000 ;
        RECT 40.045000  92.475000 44.500000  92.625000 ;
        RECT 40.135000 166.835000 48.835000 166.985000 ;
        RECT 40.195000  92.625000 44.650000  92.775000 ;
        RECT 40.285000 166.685000 48.835000 166.835000 ;
        RECT 40.345000  92.775000 44.800000  92.925000 ;
        RECT 40.435000 166.535000 48.835000 166.685000 ;
        RECT 40.495000  92.925000 44.950000  93.075000 ;
        RECT 40.585000 166.385000 48.835000 166.535000 ;
        RECT 40.645000  93.075000 45.100000  93.225000 ;
        RECT 40.735000 166.235000 48.835000 166.385000 ;
        RECT 40.795000  93.225000 45.250000  93.375000 ;
        RECT 40.885000 166.085000 48.835000 166.235000 ;
        RECT 40.945000  93.375000 45.400000  93.525000 ;
        RECT 41.035000 165.935000 48.835000 166.085000 ;
        RECT 41.050000  83.980000 48.870000  84.130000 ;
        RECT 41.095000  93.525000 45.550000  93.675000 ;
        RECT 41.185000 165.785000 48.835000 165.935000 ;
        RECT 41.200000  84.130000 48.870000  84.280000 ;
        RECT 41.245000  93.675000 45.700000  93.825000 ;
        RECT 41.335000 165.635000 48.835000 165.785000 ;
        RECT 41.350000  84.280000 48.870000  84.430000 ;
        RECT 41.395000  93.825000 45.850000  93.975000 ;
        RECT 41.485000 165.485000 48.835000 165.635000 ;
        RECT 41.500000  84.430000 48.870000  84.580000 ;
        RECT 41.545000  93.975000 46.000000  94.125000 ;
        RECT 41.610000  84.580000 48.870000  84.690000 ;
        RECT 41.610000  84.690000 48.870000  84.810000 ;
        RECT 41.610000  84.810000 48.870000  84.960000 ;
        RECT 41.610000  84.960000 49.020000  85.110000 ;
        RECT 41.610000  85.110000 49.170000  85.260000 ;
        RECT 41.610000  85.260000 49.320000  85.410000 ;
        RECT 41.610000  85.410000 49.470000  85.560000 ;
        RECT 41.610000  85.560000 49.620000  85.710000 ;
        RECT 41.610000  85.710000 49.770000  85.860000 ;
        RECT 41.610000  85.860000 49.920000  86.010000 ;
        RECT 41.610000  86.010000 50.070000  86.160000 ;
        RECT 41.610000  86.160000 50.220000  86.310000 ;
        RECT 41.610000  86.310000 50.370000  86.460000 ;
        RECT 41.610000  86.460000 50.520000  86.610000 ;
        RECT 41.610000  86.610000 50.670000  86.760000 ;
        RECT 41.610000  86.760000 50.820000  86.910000 ;
        RECT 41.610000  86.910000 50.970000  86.960000 ;
        RECT 41.610000  86.960000 51.020000  87.445000 ;
        RECT 41.635000 165.335000 48.835000 165.485000 ;
        RECT 41.695000  94.125000 46.150000  94.275000 ;
        RECT 41.760000  87.445000 51.020000  87.595000 ;
        RECT 41.785000 165.185000 48.835000 165.335000 ;
        RECT 41.845000  94.275000 46.300000  94.425000 ;
        RECT 41.910000  87.595000 51.020000  87.745000 ;
        RECT 41.935000 165.035000 48.835000 165.185000 ;
        RECT 41.995000  94.425000 46.450000  94.575000 ;
        RECT 42.060000  87.745000 51.020000  87.895000 ;
        RECT 42.085000 164.885000 48.835000 165.035000 ;
        RECT 42.145000  94.575000 46.600000  94.725000 ;
        RECT 42.210000  87.895000 51.020000  88.045000 ;
        RECT 42.235000 164.735000 48.835000 164.885000 ;
        RECT 42.295000  94.725000 46.750000  94.875000 ;
        RECT 42.360000  88.045000 51.020000  88.195000 ;
        RECT 42.385000 164.585000 48.835000 164.735000 ;
        RECT 42.445000  94.875000 46.900000  95.025000 ;
        RECT 42.510000  88.195000 51.020000  88.345000 ;
        RECT 42.535000 164.435000 48.835000 164.585000 ;
        RECT 42.540000  88.345000 51.020000  88.375000 ;
        RECT 42.595000  95.025000 47.050000  95.175000 ;
        RECT 42.685000 164.285000 48.835000 164.435000 ;
        RECT 42.690000  88.375000 51.020000  88.525000 ;
        RECT 42.745000  95.175000 47.200000  95.325000 ;
        RECT 42.835000  95.325000 47.350000  95.415000 ;
        RECT 42.835000  95.415000 47.440000  95.565000 ;
        RECT 42.835000  95.565000 47.590000  95.715000 ;
        RECT 42.835000  95.715000 47.740000  95.865000 ;
        RECT 42.835000  95.865000 47.890000  96.015000 ;
        RECT 42.835000  96.015000 48.040000  96.165000 ;
        RECT 42.835000  96.165000 48.190000  96.315000 ;
        RECT 42.835000  96.315000 48.340000  96.465000 ;
        RECT 42.835000  96.465000 48.490000  96.615000 ;
        RECT 42.835000  96.615000 48.640000  96.765000 ;
        RECT 42.835000  96.765000 48.790000  96.810000 ;
        RECT 42.835000  96.810000 48.835000 164.135000 ;
        RECT 42.835000 164.135000 48.835000 164.285000 ;
        RECT 42.840000  88.525000 51.170000  88.675000 ;
        RECT 42.990000  88.675000 51.320000  88.825000 ;
        RECT 43.140000  88.825000 51.470000  88.975000 ;
        RECT 43.290000  88.975000 51.620000  89.125000 ;
        RECT 43.440000  89.125000 51.770000  89.275000 ;
        RECT 43.590000  89.275000 51.920000  89.425000 ;
        RECT 43.740000  89.425000 52.070000  89.575000 ;
        RECT 43.890000  89.575000 52.220000  89.725000 ;
        RECT 44.040000  89.725000 52.370000  89.875000 ;
        RECT 44.190000  89.875000 52.520000  90.025000 ;
        RECT 44.340000  90.025000 52.670000  90.175000 ;
        RECT 44.490000  90.175000 52.820000  90.325000 ;
        RECT 44.640000  90.325000 52.970000  90.475000 ;
        RECT 44.790000  90.475000 53.120000  90.625000 ;
        RECT 44.940000  90.625000 53.270000  90.775000 ;
        RECT 45.090000  90.775000 53.420000  90.925000 ;
        RECT 45.240000  90.925000 53.570000  91.075000 ;
        RECT 45.390000  91.075000 53.720000  91.225000 ;
        RECT 45.540000  91.225000 53.870000  91.375000 ;
        RECT 45.690000  91.375000 54.020000  91.525000 ;
        RECT 45.840000  91.525000 54.170000  91.675000 ;
        RECT 45.990000  91.675000 54.320000  91.825000 ;
        RECT 46.140000  91.825000 54.470000  91.975000 ;
        RECT 46.290000  91.975000 54.620000  92.125000 ;
        RECT 46.440000  92.125000 54.770000  92.275000 ;
        RECT 46.590000  92.275000 54.920000  92.425000 ;
        RECT 46.740000  92.425000 55.070000  92.575000 ;
        RECT 46.890000  92.575000 55.220000  92.725000 ;
        RECT 47.040000  92.725000 55.370000  92.875000 ;
        RECT 47.190000  92.875000 55.520000  93.025000 ;
        RECT 47.340000  93.025000 55.670000  93.175000 ;
        RECT 47.490000  93.175000 55.820000  93.325000 ;
        RECT 47.640000  93.325000 55.970000  93.475000 ;
        RECT 47.790000  93.475000 56.120000  93.625000 ;
        RECT 47.940000  93.625000 56.270000  93.775000 ;
        RECT 48.090000  93.775000 56.420000  93.925000 ;
        RECT 48.240000  93.925000 56.570000  94.075000 ;
        RECT 48.390000  94.075000 56.720000  94.225000 ;
        RECT 48.540000  94.225000 56.870000  94.375000 ;
        RECT 48.690000  94.375000 57.020000  94.525000 ;
        RECT 48.840000  94.525000 57.170000  94.675000 ;
        RECT 48.990000  94.675000 57.320000  94.825000 ;
        RECT 49.140000  94.825000 57.470000  94.975000 ;
        RECT 49.290000  94.975000 57.620000  95.125000 ;
        RECT 49.440000  95.125000 57.770000  95.275000 ;
        RECT 49.590000  95.275000 57.920000  95.425000 ;
        RECT 49.740000  95.425000 58.070000  95.575000 ;
        RECT 49.870000 168.920000 60.330000 189.515000 ;
        RECT 49.890000  95.575000 58.220000  95.725000 ;
        RECT 49.980000 168.810000 60.330000 168.920000 ;
        RECT 50.040000  95.725000 58.370000  95.875000 ;
        RECT 50.130000 168.660000 60.330000 168.810000 ;
        RECT 50.190000  95.875000 58.520000  96.025000 ;
        RECT 50.280000 168.510000 60.330000 168.660000 ;
        RECT 50.340000  96.025000 58.670000  96.175000 ;
        RECT 50.430000 168.360000 60.330000 168.510000 ;
        RECT 50.490000  96.175000 58.820000  96.325000 ;
        RECT 50.580000 168.210000 60.330000 168.360000 ;
        RECT 50.640000  96.325000 58.970000  96.475000 ;
        RECT 50.730000 168.060000 60.330000 168.210000 ;
        RECT 50.790000  96.475000 59.120000  96.625000 ;
        RECT 50.880000 167.910000 60.330000 168.060000 ;
        RECT 50.940000  96.625000 59.270000  96.775000 ;
        RECT 51.030000 167.760000 60.330000 167.910000 ;
        RECT 51.090000  96.775000 59.420000  96.925000 ;
        RECT 51.180000 167.610000 60.330000 167.760000 ;
        RECT 51.240000  96.925000 59.570000  97.075000 ;
        RECT 51.330000 167.460000 60.330000 167.610000 ;
        RECT 51.390000  97.075000 59.720000  97.225000 ;
        RECT 51.480000 167.310000 60.330000 167.460000 ;
        RECT 51.540000  97.225000 59.870000  97.375000 ;
        RECT 51.630000 167.160000 60.330000 167.310000 ;
        RECT 51.690000  97.375000 60.020000  97.525000 ;
        RECT 51.780000 167.010000 60.330000 167.160000 ;
        RECT 51.840000  97.525000 60.170000  97.675000 ;
        RECT 51.850000  97.675000 60.320000  97.685000 ;
        RECT 51.930000 166.860000 60.330000 167.010000 ;
        RECT 52.000000  97.685000 60.330000  97.835000 ;
        RECT 52.080000 166.710000 60.330000 166.860000 ;
        RECT 52.150000  97.835000 60.330000  97.985000 ;
        RECT 52.230000 166.560000 60.330000 166.710000 ;
        RECT 52.300000  97.985000 60.330000  98.135000 ;
        RECT 52.380000 166.410000 60.330000 166.560000 ;
        RECT 52.450000  98.135000 60.330000  98.285000 ;
        RECT 52.530000 166.260000 60.330000 166.410000 ;
        RECT 52.600000  98.285000 60.330000  98.435000 ;
        RECT 52.680000 166.110000 60.330000 166.260000 ;
        RECT 52.750000  98.435000 60.330000  98.585000 ;
        RECT 52.830000 165.960000 60.330000 166.110000 ;
        RECT 52.900000  98.585000 60.330000  98.735000 ;
        RECT 52.980000 165.810000 60.330000 165.960000 ;
        RECT 53.050000  98.735000 60.330000  98.885000 ;
        RECT 53.130000 165.660000 60.330000 165.810000 ;
        RECT 53.200000  98.885000 60.330000  99.035000 ;
        RECT 53.280000 165.510000 60.330000 165.660000 ;
        RECT 53.350000  99.035000 60.330000  99.185000 ;
        RECT 53.430000 165.360000 60.330000 165.510000 ;
        RECT 53.500000  99.185000 60.330000  99.335000 ;
        RECT 53.580000 165.210000 60.330000 165.360000 ;
        RECT 53.650000  99.335000 60.330000  99.485000 ;
        RECT 53.730000 165.060000 60.330000 165.210000 ;
        RECT 53.800000  99.485000 60.330000  99.635000 ;
        RECT 53.880000 164.910000 60.330000 165.060000 ;
        RECT 53.950000  99.635000 60.330000  99.785000 ;
        RECT 54.030000 164.760000 60.330000 164.910000 ;
        RECT 54.100000  99.785000 60.330000  99.935000 ;
        RECT 54.180000 164.610000 60.330000 164.760000 ;
        RECT 54.250000  99.935000 60.330000 100.085000 ;
        RECT 54.330000 100.085000 60.330000 100.165000 ;
        RECT 54.330000 100.165000 60.330000 164.460000 ;
        RECT 54.330000 164.460000 60.330000 164.610000 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380000 0.000000 49.255000 69.490000 ;
    END
  END DRN_LVC2
  PIN OGC_LVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 26.210000 0.000000 27.700000 0.170000 ;
    END
  END OGC_LVC
  PIN P_CORE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.500000  0.000000 24.500000  82.660000 ;
        RECT 0.500000 82.660000 24.350000  82.810000 ;
        RECT 0.500000 82.810000 24.200000  82.960000 ;
        RECT 0.500000 82.960000 24.050000  83.110000 ;
        RECT 0.500000 83.110000 23.900000  83.260000 ;
        RECT 0.500000 83.260000 23.750000  83.410000 ;
        RECT 0.500000 83.410000 23.600000  83.560000 ;
        RECT 0.500000 83.560000 23.450000  83.710000 ;
        RECT 0.500000 83.710000 23.300000  83.860000 ;
        RECT 0.500000 83.860000 23.150000  84.010000 ;
        RECT 0.500000 84.010000 23.000000  84.160000 ;
        RECT 0.500000 84.160000 22.850000  84.310000 ;
        RECT 0.500000 84.310000 22.700000  84.460000 ;
        RECT 0.500000 84.460000 22.550000  84.610000 ;
        RECT 0.500000 84.610000 22.400000  84.760000 ;
        RECT 0.500000 84.760000 22.250000  84.910000 ;
        RECT 0.500000 84.910000 22.100000  85.060000 ;
        RECT 0.500000 85.060000 21.950000  85.210000 ;
        RECT 0.500000 85.210000 21.800000  85.360000 ;
        RECT 0.500000 85.360000 21.650000  85.510000 ;
        RECT 0.500000 85.510000 21.500000  85.660000 ;
        RECT 0.500000 85.660000 21.350000  85.810000 ;
        RECT 0.500000 85.810000 21.200000  85.960000 ;
        RECT 0.500000 85.960000 21.050000  86.110000 ;
        RECT 0.500000 86.110000 20.900000  86.260000 ;
        RECT 0.500000 86.260000 20.750000  86.410000 ;
        RECT 0.500000 86.410000 20.600000  86.560000 ;
        RECT 0.500000 86.560000 20.450000  86.710000 ;
        RECT 0.500000 86.710000 20.300000  86.860000 ;
        RECT 0.500000 86.860000 20.150000  87.010000 ;
        RECT 0.500000 87.010000 20.000000  87.160000 ;
        RECT 0.500000 87.160000 19.850000  87.310000 ;
        RECT 0.500000 87.310000 19.700000  87.460000 ;
        RECT 0.500000 87.460000 19.550000  87.610000 ;
        RECT 0.500000 87.610000 19.400000  87.760000 ;
        RECT 0.500000 87.760000 19.250000  87.910000 ;
        RECT 0.500000 87.910000 19.100000  88.060000 ;
        RECT 0.500000 88.060000 18.950000  88.210000 ;
        RECT 0.500000 88.210000 18.800000  88.360000 ;
        RECT 0.500000 88.360000 18.650000  88.510000 ;
        RECT 0.500000 88.510000 18.500000  88.660000 ;
        RECT 0.500000 88.660000 18.350000  88.810000 ;
        RECT 0.500000 88.810000 18.200000  88.960000 ;
        RECT 0.500000 88.960000 18.050000  89.110000 ;
        RECT 0.500000 89.110000 17.900000  89.260000 ;
        RECT 0.500000 89.260000 17.750000  89.410000 ;
        RECT 0.500000 89.410000 17.600000  89.560000 ;
        RECT 0.500000 89.560000 17.450000  89.710000 ;
        RECT 0.500000 89.710000 17.300000  89.860000 ;
        RECT 0.500000 89.860000 17.150000  90.010000 ;
        RECT 0.500000 90.010000 17.000000  90.160000 ;
        RECT 0.500000 90.160000 16.850000  90.310000 ;
        RECT 0.500000 90.310000 16.700000  90.460000 ;
        RECT 0.500000 90.460000 16.550000  90.610000 ;
        RECT 0.500000 90.610000 16.400000  90.760000 ;
        RECT 0.500000 90.760000 16.250000  90.910000 ;
        RECT 0.500000 90.910000 16.100000  91.060000 ;
        RECT 0.500000 91.060000 15.950000  91.210000 ;
        RECT 0.500000 91.210000 15.800000  91.360000 ;
        RECT 0.500000 91.360000 15.650000  91.510000 ;
        RECT 0.500000 91.510000 15.500000  91.660000 ;
        RECT 0.500000 91.660000 15.350000  91.810000 ;
        RECT 0.500000 91.810000 15.200000  91.960000 ;
        RECT 0.500000 91.960000 15.050000  92.110000 ;
        RECT 0.500000 92.110000 14.900000  92.260000 ;
        RECT 0.500000 92.260000 14.750000  92.410000 ;
        RECT 0.500000 92.410000 14.600000  92.560000 ;
        RECT 0.500000 92.560000 14.450000  92.710000 ;
        RECT 0.500000 92.710000 14.300000  92.860000 ;
        RECT 0.500000 92.860000 14.150000  93.010000 ;
        RECT 0.500000 93.010000 14.000000  93.160000 ;
        RECT 0.500000 93.160000 13.850000  93.310000 ;
        RECT 0.500000 93.310000 13.700000  93.460000 ;
        RECT 0.500000 93.460000 13.550000  93.610000 ;
        RECT 0.500000 93.610000 13.400000  93.760000 ;
        RECT 0.500000 93.760000 13.250000  93.910000 ;
        RECT 0.500000 93.910000 13.100000  94.060000 ;
        RECT 0.500000 94.060000 12.950000  94.210000 ;
        RECT 0.500000 94.210000 12.900000  94.260000 ;
        RECT 0.500000 94.260000 12.900000 171.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000  0.000000 74.700000  84.465000 ;
        RECT 50.905000 84.465000 74.700000  84.615000 ;
        RECT 51.055000 84.615000 74.700000  84.765000 ;
        RECT 51.205000 84.765000 74.700000  84.915000 ;
        RECT 51.355000 84.915000 74.700000  85.065000 ;
        RECT 51.505000 85.065000 74.700000  85.215000 ;
        RECT 51.655000 85.215000 74.700000  85.365000 ;
        RECT 51.805000 85.365000 74.700000  85.515000 ;
        RECT 51.955000 85.515000 74.700000  85.665000 ;
        RECT 52.105000 85.665000 74.700000  85.815000 ;
        RECT 52.255000 85.815000 74.700000  85.965000 ;
        RECT 52.405000 85.965000 74.700000  86.115000 ;
        RECT 52.555000 86.115000 74.700000  86.265000 ;
        RECT 52.705000 86.265000 74.700000  86.415000 ;
        RECT 52.855000 86.415000 74.700000  86.565000 ;
        RECT 53.005000 86.565000 74.700000  86.715000 ;
        RECT 53.155000 86.715000 74.700000  86.865000 ;
        RECT 53.305000 86.865000 74.700000  87.015000 ;
        RECT 53.455000 87.015000 74.700000  87.165000 ;
        RECT 53.605000 87.165000 74.700000  87.315000 ;
        RECT 53.755000 87.315000 74.700000  87.465000 ;
        RECT 53.905000 87.465000 74.700000  87.615000 ;
        RECT 54.055000 87.615000 74.700000  87.765000 ;
        RECT 54.205000 87.765000 74.700000  87.915000 ;
        RECT 54.355000 87.915000 74.700000  88.065000 ;
        RECT 54.505000 88.065000 74.700000  88.215000 ;
        RECT 54.655000 88.215000 74.700000  88.365000 ;
        RECT 54.805000 88.365000 74.700000  88.515000 ;
        RECT 54.955000 88.515000 74.700000  88.665000 ;
        RECT 55.105000 88.665000 74.700000  88.815000 ;
        RECT 55.255000 88.815000 74.700000  88.965000 ;
        RECT 55.405000 88.965000 74.700000  89.115000 ;
        RECT 55.555000 89.115000 74.700000  89.265000 ;
        RECT 55.705000 89.265000 74.700000  89.415000 ;
        RECT 55.855000 89.415000 74.700000  89.565000 ;
        RECT 56.005000 89.565000 74.700000  89.715000 ;
        RECT 56.155000 89.715000 74.700000  89.865000 ;
        RECT 56.305000 89.865000 74.700000  90.015000 ;
        RECT 56.455000 90.015000 74.700000  90.165000 ;
        RECT 56.605000 90.165000 74.700000  90.315000 ;
        RECT 56.755000 90.315000 74.700000  90.465000 ;
        RECT 56.905000 90.465000 74.700000  90.615000 ;
        RECT 57.055000 90.615000 74.700000  90.765000 ;
        RECT 57.205000 90.765000 74.700000  90.915000 ;
        RECT 57.355000 90.915000 74.700000  91.065000 ;
        RECT 57.505000 91.065000 74.700000  91.215000 ;
        RECT 57.655000 91.215000 74.700000  91.365000 ;
        RECT 57.805000 91.365000 74.700000  91.515000 ;
        RECT 57.955000 91.515000 74.700000  91.665000 ;
        RECT 58.105000 91.665000 74.700000  91.815000 ;
        RECT 58.255000 91.815000 74.700000  91.965000 ;
        RECT 58.405000 91.965000 74.700000  92.115000 ;
        RECT 58.555000 92.115000 74.700000  92.265000 ;
        RECT 58.705000 92.265000 74.700000  92.415000 ;
        RECT 58.855000 92.415000 74.700000  92.565000 ;
        RECT 59.005000 92.565000 74.700000  92.715000 ;
        RECT 59.155000 92.715000 74.700000  92.865000 ;
        RECT 59.305000 92.865000 74.700000  93.015000 ;
        RECT 59.455000 93.015000 74.700000  93.165000 ;
        RECT 59.605000 93.165000 74.700000  93.315000 ;
        RECT 59.755000 93.315000 74.700000  93.465000 ;
        RECT 59.905000 93.465000 74.700000  93.615000 ;
        RECT 60.055000 93.615000 74.700000  93.765000 ;
        RECT 60.205000 93.765000 74.700000  93.915000 ;
        RECT 60.355000 93.915000 74.700000  94.065000 ;
        RECT 60.505000 94.065000 74.700000  94.215000 ;
        RECT 60.655000 94.215000 74.700000  94.365000 ;
        RECT 60.805000 94.365000 74.700000  94.515000 ;
        RECT 60.955000 94.515000 74.700000  94.665000 ;
        RECT 61.105000 94.665000 74.700000  94.815000 ;
        RECT 61.255000 94.815000 74.700000  94.965000 ;
        RECT 61.405000 94.965000 74.700000  95.115000 ;
        RECT 61.555000 95.115000 74.700000  95.265000 ;
        RECT 61.705000 95.265000 74.700000  95.415000 ;
        RECT 61.855000 95.415000 74.700000  95.565000 ;
        RECT 62.005000 95.565000 74.700000  95.715000 ;
        RECT 62.045000 95.715000 74.700000  95.755000 ;
        RECT 62.045000 95.755000 74.700000 172.235000 ;
    END
  END P_CORE
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT  0.500000   0.000000 20.495000   1.485000 ;
        RECT  0.500000   1.485000 20.425000   1.555000 ;
        RECT  0.500000   1.555000 20.355000   1.625000 ;
        RECT  0.500000   1.625000 20.285000   1.695000 ;
        RECT  0.500000   1.695000 20.215000   1.765000 ;
        RECT  0.500000   1.765000 20.145000   1.835000 ;
        RECT  0.500000   1.835000 20.075000   1.905000 ;
        RECT  0.500000   1.905000 20.005000   1.975000 ;
        RECT  0.500000   1.975000 19.935000   2.045000 ;
        RECT  0.500000   2.045000 19.865000   2.115000 ;
        RECT  0.500000   2.115000 19.795000   2.185000 ;
        RECT  0.500000   2.185000 19.725000   2.255000 ;
        RECT  0.500000   2.255000 19.655000   2.325000 ;
        RECT  0.500000   2.325000 19.585000   2.395000 ;
        RECT  0.500000   2.395000 19.515000   2.465000 ;
        RECT  0.500000   2.465000 19.445000   2.535000 ;
        RECT  0.500000   2.535000 19.375000   2.605000 ;
        RECT  0.500000   2.605000 19.305000   2.675000 ;
        RECT  0.500000   2.675000 19.235000   2.745000 ;
        RECT  0.500000   2.745000 19.165000   2.815000 ;
        RECT  0.500000   2.815000 19.095000   2.885000 ;
        RECT  0.500000   2.885000 19.025000   2.955000 ;
        RECT  0.500000   2.955000 18.955000   3.025000 ;
        RECT  0.500000   3.025000 18.885000   3.095000 ;
        RECT  0.500000   3.095000 18.815000   3.165000 ;
        RECT  0.500000   3.165000 18.745000   3.235000 ;
        RECT  0.500000   3.235000 18.675000   3.305000 ;
        RECT  0.500000   3.305000 18.605000   3.375000 ;
        RECT  0.500000   3.375000 18.535000   3.445000 ;
        RECT  0.500000   3.445000 18.465000   3.515000 ;
        RECT  0.500000   3.515000 18.395000   3.585000 ;
        RECT  0.500000   3.585000 18.325000   3.655000 ;
        RECT  0.500000   3.655000 18.255000   3.725000 ;
        RECT  0.500000   3.725000 18.185000   3.795000 ;
        RECT  0.500000   3.795000 18.115000   3.865000 ;
        RECT  0.500000   3.865000 18.045000   3.935000 ;
        RECT  0.500000   3.935000 17.975000   4.005000 ;
        RECT  0.500000   4.005000 17.905000   4.075000 ;
        RECT  0.500000   4.075000 17.835000   4.145000 ;
        RECT  0.500000   4.145000 17.765000   4.215000 ;
        RECT  0.500000   4.215000 17.695000   4.285000 ;
        RECT  0.500000   4.285000 17.625000   4.355000 ;
        RECT  0.500000   4.355000 17.555000   4.425000 ;
        RECT  0.500000   4.425000 17.485000   4.495000 ;
        RECT  0.500000   4.495000 17.415000   4.565000 ;
        RECT  0.500000   4.565000 17.345000   4.635000 ;
        RECT  0.500000   4.635000 17.275000   4.705000 ;
        RECT  0.500000   4.705000 17.205000   4.775000 ;
        RECT  0.500000   4.775000 17.135000   4.845000 ;
        RECT  0.500000   4.845000 17.065000   4.915000 ;
        RECT  0.500000   4.915000 16.995000   4.985000 ;
        RECT  0.500000   4.985000 16.925000   5.055000 ;
        RECT  0.500000   5.055000 16.860000   5.120000 ;
        RECT  0.500000   5.120000 16.860000   7.655000 ;
        RECT  0.500000   7.655000 10.745000   7.725000 ;
        RECT  0.500000   7.725000 10.675000   7.795000 ;
        RECT  0.500000   7.795000 10.605000   7.865000 ;
        RECT  0.500000   7.865000 10.535000   7.935000 ;
        RECT  0.500000   7.935000 10.465000   8.005000 ;
        RECT  0.500000   8.005000 10.420000   8.050000 ;
        RECT  0.500000   8.050000 10.420000   9.820000 ;
        RECT  0.500000   9.820000 10.420000   9.890000 ;
        RECT  0.500000   9.890000 10.490000   9.960000 ;
        RECT  0.500000   9.960000 10.560000  10.030000 ;
        RECT  0.500000  10.030000 10.630000  10.100000 ;
        RECT  0.500000  10.100000 10.700000  10.170000 ;
        RECT  0.500000  10.170000 10.770000  10.215000 ;
        RECT  0.500000  10.215000 55.595000  17.080000 ;
        RECT  0.500000  17.080000 21.785000  17.150000 ;
        RECT  0.500000  17.150000 21.715000  17.220000 ;
        RECT  0.500000  17.220000 21.645000  17.290000 ;
        RECT  0.500000  17.290000 21.575000  17.360000 ;
        RECT  0.500000  17.360000 21.505000  17.430000 ;
        RECT  0.500000  17.430000 21.435000  17.500000 ;
        RECT  0.500000  17.500000 21.365000  17.570000 ;
        RECT  0.500000  17.570000 21.295000  17.640000 ;
        RECT  0.500000  17.640000 21.225000  17.710000 ;
        RECT  0.500000  17.710000 21.155000  17.780000 ;
        RECT  0.500000  17.780000 21.085000  17.850000 ;
        RECT  0.500000  17.850000 21.015000  17.920000 ;
        RECT  0.500000  17.920000 20.945000  17.990000 ;
        RECT  0.500000  17.990000 20.875000  18.060000 ;
        RECT  0.500000  18.060000 20.805000  18.130000 ;
        RECT  0.500000  18.130000 20.735000  18.200000 ;
        RECT  0.500000  18.200000 20.665000  18.270000 ;
        RECT  0.500000  18.270000 20.595000  18.340000 ;
        RECT  0.500000  18.340000 20.525000  18.410000 ;
        RECT  0.500000  18.410000 20.455000  18.480000 ;
        RECT  0.500000  18.480000 20.385000  18.550000 ;
        RECT  0.500000  18.550000 20.315000  18.620000 ;
        RECT  0.500000  18.620000 20.245000  18.690000 ;
        RECT  0.500000  18.690000 20.175000  18.760000 ;
        RECT  0.500000  18.760000 20.105000  18.830000 ;
        RECT  0.500000  18.830000 20.035000  18.900000 ;
        RECT  0.500000  18.900000 19.965000  18.970000 ;
        RECT  0.500000  18.970000 19.895000  19.040000 ;
        RECT  0.500000  19.040000 19.825000  19.110000 ;
        RECT  0.500000  19.110000 19.755000  19.180000 ;
        RECT  0.500000  19.180000 19.685000  19.250000 ;
        RECT  0.500000  19.250000 19.615000  19.320000 ;
        RECT  0.500000  19.320000 19.545000  19.390000 ;
        RECT  0.500000  19.390000 19.475000  19.460000 ;
        RECT  0.500000  19.460000 19.405000  19.530000 ;
        RECT  0.500000  19.530000 19.335000  19.600000 ;
        RECT  0.500000  19.600000 19.265000  19.670000 ;
        RECT  0.500000  19.670000 19.195000  19.740000 ;
        RECT  0.500000  19.740000 19.125000  19.810000 ;
        RECT  0.500000  19.810000 19.055000  19.880000 ;
        RECT  0.500000  19.880000 18.985000  19.950000 ;
        RECT  0.500000  19.950000 18.915000  20.020000 ;
        RECT  0.500000  20.020000 18.845000  20.090000 ;
        RECT  0.500000  20.090000 18.775000  20.160000 ;
        RECT  0.500000  20.160000 18.705000  20.230000 ;
        RECT  0.500000  20.230000 18.635000  20.300000 ;
        RECT  0.500000  20.300000 18.565000  20.370000 ;
        RECT  0.500000  20.370000 18.495000  20.440000 ;
        RECT  0.500000  20.440000 18.425000  20.510000 ;
        RECT  0.500000  20.510000 18.355000  20.580000 ;
        RECT  0.500000  20.580000 18.285000  20.650000 ;
        RECT  0.500000  20.650000 18.215000  20.720000 ;
        RECT  0.500000  20.720000 18.145000  20.790000 ;
        RECT  0.500000  20.790000 18.075000  20.860000 ;
        RECT  0.500000  20.860000 18.005000  20.930000 ;
        RECT  0.500000  20.930000 17.935000  21.000000 ;
        RECT  0.500000  21.000000 17.865000  21.070000 ;
        RECT  0.500000  21.070000 17.795000  21.140000 ;
        RECT  0.500000  21.140000 17.725000  21.210000 ;
        RECT  0.500000  21.210000 17.655000  21.280000 ;
        RECT  0.500000  21.280000 17.585000  21.350000 ;
        RECT  0.500000  21.350000 17.515000  21.420000 ;
        RECT  0.500000  21.420000 17.445000  21.490000 ;
        RECT  0.500000  21.490000 17.375000  21.560000 ;
        RECT  0.500000  21.560000 17.305000  21.630000 ;
        RECT  0.500000  21.630000 17.235000  21.700000 ;
        RECT  0.500000  21.700000 17.165000  21.770000 ;
        RECT  0.500000  21.770000 17.095000  21.840000 ;
        RECT  0.500000  21.840000 17.025000  21.910000 ;
        RECT  0.500000  21.910000 16.955000  21.980000 ;
        RECT  0.500000  21.980000 16.885000  22.050000 ;
        RECT  0.500000  22.050000 16.815000  22.120000 ;
        RECT  0.500000  22.120000 16.745000  22.190000 ;
        RECT  0.500000  22.190000 16.675000  22.260000 ;
        RECT  0.500000  22.260000 16.605000  22.330000 ;
        RECT  0.500000  22.330000 16.535000  22.400000 ;
        RECT  0.500000  22.400000 16.465000  22.470000 ;
        RECT  0.500000  22.470000 16.395000  22.540000 ;
        RECT  0.500000  22.540000 16.325000  22.610000 ;
        RECT  0.500000  22.610000 16.255000  22.680000 ;
        RECT  0.500000  22.680000 16.185000  22.750000 ;
        RECT  0.500000  22.750000 16.115000  22.820000 ;
        RECT  0.500000  22.820000 16.045000  22.890000 ;
        RECT  0.500000  22.890000 15.975000  22.960000 ;
        RECT  0.500000  22.960000 15.905000  23.030000 ;
        RECT  0.500000  23.030000 15.835000  23.100000 ;
        RECT  0.500000  23.100000 15.765000  23.170000 ;
        RECT  0.500000  23.170000 15.695000  23.240000 ;
        RECT  0.500000  23.240000 15.625000  23.310000 ;
        RECT  0.500000  23.310000 15.555000  23.380000 ;
        RECT  0.500000  23.380000 15.485000  23.450000 ;
        RECT  0.500000  23.450000 15.415000  23.520000 ;
        RECT  0.500000  23.520000 15.345000  23.590000 ;
        RECT  0.500000  23.590000 15.275000  23.660000 ;
        RECT  0.500000  23.660000 15.205000  23.730000 ;
        RECT  0.500000  23.730000 15.135000  23.800000 ;
        RECT  0.500000  23.800000 15.065000  23.870000 ;
        RECT  0.500000  23.870000 14.995000  23.940000 ;
        RECT  0.500000  23.940000 14.925000  24.010000 ;
        RECT  0.500000  24.010000 14.855000  24.080000 ;
        RECT  0.500000  24.080000 14.785000  24.150000 ;
        RECT  0.500000  24.150000 14.715000  24.220000 ;
        RECT  0.500000  24.220000 14.645000  24.290000 ;
        RECT  0.500000  24.290000 14.575000  24.360000 ;
        RECT  0.500000  24.360000 14.505000  24.430000 ;
        RECT  0.500000  24.430000 14.435000  24.500000 ;
        RECT  0.500000  24.500000 14.365000  24.570000 ;
        RECT  0.500000  24.570000 14.295000  24.640000 ;
        RECT  0.500000  24.640000 14.225000  24.710000 ;
        RECT  0.500000  24.710000 14.155000  24.780000 ;
        RECT  0.500000  24.780000 14.085000  24.850000 ;
        RECT  0.500000  24.850000 14.015000  24.920000 ;
        RECT  0.500000  24.920000 13.945000  24.990000 ;
        RECT  0.500000  24.990000 13.875000  25.060000 ;
        RECT  0.500000  25.060000 13.805000  25.130000 ;
        RECT  0.500000  25.130000 13.750000  25.185000 ;
        RECT  0.500000  25.185000 13.750000  74.295000 ;
        RECT  0.500000  74.295000 13.750000  74.365000 ;
        RECT  0.500000  74.365000 13.820000  74.435000 ;
        RECT  0.500000  74.435000 13.890000  74.505000 ;
        RECT  0.500000  74.505000 13.960000 129.935000 ;
        RECT  0.500000 129.935000 13.960000 130.005000 ;
        RECT  0.500000 130.005000 14.030000 130.075000 ;
        RECT  0.500000 130.075000 14.100000 130.145000 ;
        RECT  0.500000 130.145000 14.170000 130.215000 ;
        RECT  0.500000 130.215000 14.240000 130.285000 ;
        RECT  0.500000 130.285000 14.310000 130.355000 ;
        RECT  0.500000 130.355000 14.380000 130.425000 ;
        RECT  0.500000 130.425000 14.450000 130.495000 ;
        RECT  0.500000 130.495000 14.520000 130.565000 ;
        RECT  0.500000 130.565000 14.590000 130.635000 ;
        RECT  0.500000 130.635000 14.660000 130.705000 ;
        RECT  0.500000 130.705000 14.730000 130.775000 ;
        RECT  0.500000 130.775000 14.800000 130.845000 ;
        RECT  0.500000 130.845000 14.870000 130.915000 ;
        RECT  0.500000 130.915000 14.940000 130.985000 ;
        RECT  0.500000 130.985000 68.010000 133.630000 ;
        RECT  0.500000 133.630000 14.940000 133.700000 ;
        RECT  0.500000 133.700000 14.870000 133.770000 ;
        RECT  0.500000 133.770000 14.800000 133.840000 ;
        RECT  0.500000 133.840000 14.730000 133.910000 ;
        RECT  0.500000 133.910000 14.660000 133.980000 ;
        RECT  0.500000 133.980000 14.590000 134.050000 ;
        RECT  0.500000 134.050000 14.520000 134.120000 ;
        RECT  0.500000 134.120000 14.450000 134.190000 ;
        RECT  0.500000 134.190000 14.380000 134.260000 ;
        RECT  0.500000 134.260000 14.310000 134.330000 ;
        RECT  0.500000 134.330000 14.240000 134.400000 ;
        RECT  0.500000 134.400000 14.170000 134.470000 ;
        RECT  0.500000 134.470000 14.100000 134.540000 ;
        RECT  0.500000 134.540000 14.030000 134.610000 ;
        RECT  0.500000 134.610000 13.960000 134.680000 ;
        RECT  0.500000 134.680000 13.960000 139.940000 ;
        RECT  0.500000 139.940000 13.960000 140.010000 ;
        RECT  0.500000 140.010000 14.030000 140.080000 ;
        RECT  0.500000 140.080000 14.100000 140.150000 ;
        RECT  0.500000 140.150000 14.170000 140.220000 ;
        RECT  0.500000 140.220000 14.240000 140.290000 ;
        RECT  0.500000 140.290000 14.310000 140.360000 ;
        RECT  0.500000 140.360000 14.380000 140.430000 ;
        RECT  0.500000 140.430000 14.450000 140.500000 ;
        RECT  0.500000 140.500000 14.520000 140.570000 ;
        RECT  0.500000 140.570000 14.590000 140.640000 ;
        RECT  0.500000 140.640000 14.660000 140.710000 ;
        RECT  0.500000 140.710000 14.730000 140.780000 ;
        RECT  0.500000 140.780000 14.800000 140.850000 ;
        RECT  0.500000 140.850000 14.870000 140.920000 ;
        RECT  0.500000 140.920000 14.940000 140.990000 ;
        RECT  0.500000 140.990000 68.010000 143.630000 ;
        RECT  0.500000 143.630000 14.940000 143.700000 ;
        RECT  0.500000 143.700000 14.870000 143.770000 ;
        RECT  0.500000 143.770000 14.800000 143.840000 ;
        RECT  0.500000 143.840000 14.730000 143.910000 ;
        RECT  0.500000 143.910000 14.660000 143.980000 ;
        RECT  0.500000 143.980000 14.590000 144.050000 ;
        RECT  0.500000 144.050000 14.520000 144.120000 ;
        RECT  0.500000 144.120000 14.450000 144.190000 ;
        RECT  0.500000 144.190000 14.380000 144.260000 ;
        RECT  0.500000 144.260000 14.310000 144.330000 ;
        RECT  0.500000 144.330000 14.240000 144.400000 ;
        RECT  0.500000 144.400000 14.170000 144.470000 ;
        RECT  0.500000 144.470000 14.100000 144.540000 ;
        RECT  0.500000 144.540000 14.030000 144.610000 ;
        RECT  0.500000 144.610000 13.960000 144.680000 ;
        RECT  0.500000 144.680000 13.960000 149.940000 ;
        RECT  0.500000 149.940000 13.960000 150.010000 ;
        RECT  0.500000 150.010000 14.030000 150.080000 ;
        RECT  0.500000 150.080000 14.100000 150.150000 ;
        RECT  0.500000 150.150000 14.170000 150.220000 ;
        RECT  0.500000 150.220000 14.240000 150.290000 ;
        RECT  0.500000 150.290000 14.310000 150.360000 ;
        RECT  0.500000 150.360000 14.380000 150.430000 ;
        RECT  0.500000 150.430000 14.450000 150.500000 ;
        RECT  0.500000 150.500000 14.520000 150.570000 ;
        RECT  0.500000 150.570000 14.590000 150.640000 ;
        RECT  0.500000 150.640000 14.660000 150.710000 ;
        RECT  0.500000 150.710000 14.730000 150.780000 ;
        RECT  0.500000 150.780000 14.800000 150.850000 ;
        RECT  0.500000 150.850000 14.870000 150.920000 ;
        RECT  0.500000 150.920000 14.940000 150.990000 ;
        RECT  0.500000 150.990000 68.010000 153.630000 ;
        RECT  0.500000 153.630000 14.940000 153.700000 ;
        RECT  0.500000 153.700000 14.870000 153.770000 ;
        RECT  0.500000 153.770000 14.800000 153.840000 ;
        RECT  0.500000 153.840000 14.730000 153.910000 ;
        RECT  0.500000 153.910000 14.660000 153.980000 ;
        RECT  0.500000 153.980000 14.590000 154.050000 ;
        RECT  0.500000 154.050000 14.520000 154.120000 ;
        RECT  0.500000 154.120000 14.450000 154.190000 ;
        RECT  0.500000 154.190000 14.380000 154.260000 ;
        RECT  0.500000 154.260000 14.310000 154.330000 ;
        RECT  0.500000 154.330000 14.240000 154.400000 ;
        RECT  0.500000 154.400000 14.170000 154.470000 ;
        RECT  0.500000 154.470000 14.100000 154.540000 ;
        RECT  0.500000 154.540000 14.030000 154.610000 ;
        RECT  0.500000 154.610000 13.960000 154.680000 ;
        RECT  0.500000 154.680000 13.960000 159.940000 ;
        RECT  0.500000 159.940000 13.960000 160.010000 ;
        RECT  0.500000 160.010000 14.030000 160.080000 ;
        RECT  0.500000 160.080000 14.100000 160.150000 ;
        RECT  0.500000 160.150000 14.170000 160.220000 ;
        RECT  0.500000 160.220000 14.240000 160.290000 ;
        RECT  0.500000 160.290000 14.310000 160.360000 ;
        RECT  0.500000 160.360000 14.380000 160.430000 ;
        RECT  0.500000 160.430000 14.450000 160.500000 ;
        RECT  0.500000 160.500000 14.520000 160.570000 ;
        RECT  0.500000 160.570000 14.590000 160.640000 ;
        RECT  0.500000 160.640000 14.660000 160.710000 ;
        RECT  0.500000 160.710000 14.730000 160.780000 ;
        RECT  0.500000 160.780000 14.800000 160.850000 ;
        RECT  0.500000 160.850000 14.870000 160.920000 ;
        RECT  0.500000 160.920000 14.940000 160.990000 ;
        RECT  0.500000 160.990000 68.010000 163.630000 ;
        RECT  0.500000 163.630000 14.940000 163.700000 ;
        RECT  0.500000 163.700000 14.870000 163.770000 ;
        RECT  0.500000 163.770000 14.800000 163.840000 ;
        RECT  0.500000 163.840000 14.730000 163.910000 ;
        RECT  0.500000 163.910000 14.660000 163.980000 ;
        RECT  0.500000 163.980000 14.590000 164.050000 ;
        RECT  0.500000 164.050000 14.520000 164.120000 ;
        RECT  0.500000 164.120000 14.450000 164.190000 ;
        RECT  0.500000 164.190000 14.380000 164.260000 ;
        RECT  0.500000 164.260000 14.310000 164.330000 ;
        RECT  0.500000 164.330000 14.240000 164.400000 ;
        RECT  0.500000 164.400000 14.170000 164.470000 ;
        RECT  0.500000 164.470000 14.100000 164.540000 ;
        RECT  0.500000 164.540000 14.030000 164.610000 ;
        RECT  0.500000 164.610000 13.960000 164.680000 ;
        RECT  0.500000 164.680000 13.960000 169.940000 ;
        RECT  0.500000 169.940000 13.960000 170.010000 ;
        RECT  0.500000 170.010000 14.030000 170.080000 ;
        RECT  0.500000 170.080000 14.100000 170.150000 ;
        RECT  0.500000 170.150000 14.170000 170.220000 ;
        RECT  0.500000 170.220000 14.240000 170.290000 ;
        RECT  0.500000 170.290000 14.310000 170.360000 ;
        RECT  0.500000 170.360000 14.380000 170.430000 ;
        RECT  0.500000 170.430000 14.450000 170.500000 ;
        RECT  0.500000 170.500000 14.520000 170.570000 ;
        RECT  0.500000 170.570000 14.590000 170.640000 ;
        RECT  0.500000 170.640000 14.660000 170.710000 ;
        RECT  0.500000 170.710000 14.730000 170.780000 ;
        RECT  0.500000 170.780000 14.800000 170.850000 ;
        RECT  0.500000 170.850000 14.870000 170.920000 ;
        RECT  0.500000 170.920000 14.940000 170.990000 ;
        RECT  0.500000 170.990000 68.010000 173.630000 ;
        RECT  0.500000 173.630000 14.940000 173.700000 ;
        RECT  0.500000 173.700000 14.870000 173.770000 ;
        RECT  0.500000 173.770000 14.800000 173.840000 ;
        RECT  0.500000 173.840000 14.730000 173.910000 ;
        RECT  0.500000 173.910000 14.660000 173.980000 ;
        RECT  0.500000 173.980000 14.590000 174.050000 ;
        RECT  0.500000 174.050000 14.520000 174.120000 ;
        RECT  0.500000 174.120000 14.450000 174.190000 ;
        RECT  0.500000 174.190000 14.380000 174.260000 ;
        RECT  0.500000 174.260000 14.310000 174.330000 ;
        RECT  0.500000 174.330000 14.240000 174.400000 ;
        RECT  0.500000 174.400000 14.170000 174.470000 ;
        RECT  0.500000 174.470000 14.100000 174.540000 ;
        RECT  0.500000 174.540000 14.030000 174.610000 ;
        RECT  0.500000 174.610000 13.960000 174.680000 ;
        RECT  0.500000 174.680000 13.960000 179.940000 ;
        RECT  0.500000 179.940000 13.960000 180.010000 ;
        RECT  0.500000 180.010000 14.030000 180.080000 ;
        RECT  0.500000 180.080000 14.100000 180.150000 ;
        RECT  0.500000 180.150000 14.170000 180.220000 ;
        RECT  0.500000 180.220000 14.240000 180.290000 ;
        RECT  0.500000 180.290000 14.310000 180.360000 ;
        RECT  0.500000 180.360000 14.380000 180.430000 ;
        RECT  0.500000 180.430000 14.450000 180.500000 ;
        RECT  0.500000 180.500000 14.520000 180.570000 ;
        RECT  0.500000 180.570000 14.590000 180.640000 ;
        RECT  0.500000 180.640000 14.660000 180.710000 ;
        RECT  0.500000 180.710000 14.730000 180.780000 ;
        RECT  0.500000 180.780000 14.800000 180.850000 ;
        RECT  0.500000 180.850000 14.870000 180.920000 ;
        RECT  0.500000 180.920000 14.940000 180.990000 ;
        RECT  0.500000 180.990000 68.010000 183.630000 ;
        RECT  0.500000 183.630000 14.940000 183.700000 ;
        RECT  0.500000 183.700000 14.870000 183.770000 ;
        RECT  0.500000 183.770000 14.800000 183.840000 ;
        RECT  0.500000 183.840000 14.730000 183.910000 ;
        RECT  0.500000 183.910000 14.660000 183.980000 ;
        RECT  0.500000 183.980000 14.590000 184.050000 ;
        RECT  0.500000 184.050000 14.520000 184.120000 ;
        RECT  0.500000 184.120000 14.450000 184.190000 ;
        RECT  0.500000 184.190000 14.380000 184.260000 ;
        RECT  0.500000 184.260000 14.310000 184.330000 ;
        RECT  0.500000 184.330000 14.240000 184.400000 ;
        RECT  0.500000 184.400000 14.170000 184.470000 ;
        RECT  0.500000 184.470000 14.100000 184.540000 ;
        RECT  0.500000 184.540000 14.030000 184.610000 ;
        RECT  0.500000 184.610000 13.960000 184.680000 ;
        RECT  0.500000 184.680000 13.960000 189.940000 ;
        RECT  0.500000 189.940000 13.960000 190.010000 ;
        RECT  0.500000 190.010000 14.030000 190.080000 ;
        RECT  0.500000 190.080000 14.100000 190.150000 ;
        RECT  0.500000 190.150000 14.170000 190.220000 ;
        RECT  0.500000 190.220000 14.240000 190.290000 ;
        RECT  0.500000 190.290000 14.310000 190.360000 ;
        RECT  0.500000 190.360000 14.380000 190.430000 ;
        RECT  0.500000 190.430000 14.450000 190.500000 ;
        RECT  0.500000 190.500000 14.520000 190.570000 ;
        RECT  0.500000 190.570000 14.590000 190.640000 ;
        RECT  0.500000 190.640000 14.660000 190.710000 ;
        RECT  0.500000 190.710000 14.730000 190.780000 ;
        RECT  0.500000 190.780000 14.800000 190.850000 ;
        RECT  0.500000 190.850000 14.870000 190.920000 ;
        RECT  0.500000 190.920000 14.940000 190.990000 ;
        RECT  0.500000 190.990000 68.010000 193.630000 ;
        RECT 11.635000  10.210000 55.595000  10.215000 ;
        RECT 11.695000   7.655000 16.860000   7.725000 ;
        RECT 11.700000  10.145000 55.595000  10.210000 ;
        RECT 11.765000   7.725000 16.860000   7.795000 ;
        RECT 11.765000  10.080000 55.595000  10.145000 ;
        RECT 11.805000  10.040000 17.535000  10.080000 ;
        RECT 11.835000   7.795000 16.860000   7.865000 ;
        RECT 11.875000   9.970000 17.465000  10.040000 ;
        RECT 11.905000   7.865000 16.860000   7.935000 ;
        RECT 11.945000   9.900000 17.395000   9.970000 ;
        RECT 11.975000   7.935000 16.860000   8.005000 ;
        RECT 12.015000   8.005000 16.860000   8.045000 ;
        RECT 12.015000   8.045000 16.860000   9.365000 ;
        RECT 12.015000   9.365000 16.860000   9.435000 ;
        RECT 12.015000   9.435000 16.930000   9.505000 ;
        RECT 12.015000   9.505000 17.000000   9.575000 ;
        RECT 12.015000   9.575000 17.070000   9.645000 ;
        RECT 12.015000   9.645000 17.140000   9.715000 ;
        RECT 12.015000   9.715000 17.210000   9.785000 ;
        RECT 12.015000   9.785000 17.280000   9.830000 ;
        RECT 12.015000   9.830000 17.325000   9.900000 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 16.135000 31.010000 74.700000 33.650000 ;
        RECT 16.135000 40.990000 74.700000 43.630000 ;
        RECT 16.135000 51.010000 74.700000 53.650000 ;
        RECT 16.135000 60.990000 74.700000 63.630000 ;
        RECT 16.135000 70.990000 74.700000 73.630000 ;
        RECT 54.095000  0.000000 74.700000  7.815000 ;
        RECT 54.095000 19.990000 74.700000 21.695000 ;
        RECT 54.150000 19.935000 74.700000 19.990000 ;
        RECT 54.165000  7.815000 74.700000  7.885000 ;
        RECT 54.220000 19.865000 74.700000 19.935000 ;
        RECT 54.235000  7.885000 74.700000  7.955000 ;
        RECT 54.290000 19.795000 74.700000 19.865000 ;
        RECT 54.305000  7.955000 74.700000  8.025000 ;
        RECT 54.360000 19.725000 74.700000 19.795000 ;
        RECT 54.375000  8.025000 74.700000  8.095000 ;
        RECT 54.430000 19.655000 74.700000 19.725000 ;
        RECT 54.445000  8.095000 74.700000  8.165000 ;
        RECT 54.500000 19.585000 74.700000 19.655000 ;
        RECT 54.515000  8.165000 74.700000  8.235000 ;
        RECT 54.570000 19.515000 74.700000 19.585000 ;
        RECT 54.585000  8.235000 74.700000  8.305000 ;
        RECT 54.640000 19.445000 74.700000 19.515000 ;
        RECT 54.655000  8.305000 74.700000  8.375000 ;
        RECT 54.710000 19.375000 74.700000 19.445000 ;
        RECT 54.725000  8.375000 74.700000  8.445000 ;
        RECT 54.780000 19.305000 74.700000 19.375000 ;
        RECT 54.795000  8.445000 74.700000  8.515000 ;
        RECT 54.850000 19.235000 74.700000 19.305000 ;
        RECT 54.865000  8.515000 74.700000  8.585000 ;
        RECT 54.920000 19.165000 74.700000 19.235000 ;
        RECT 54.935000  8.585000 74.700000  8.655000 ;
        RECT 54.990000 19.095000 74.700000 19.165000 ;
        RECT 55.005000  8.655000 74.700000  8.725000 ;
        RECT 55.060000 19.025000 74.700000 19.095000 ;
        RECT 55.075000  8.725000 74.700000  8.795000 ;
        RECT 55.130000 18.955000 74.700000 19.025000 ;
        RECT 55.145000  8.795000 74.700000  8.865000 ;
        RECT 55.200000 18.885000 74.700000 18.955000 ;
        RECT 55.215000  8.865000 74.700000  8.935000 ;
        RECT 55.270000 18.815000 74.700000 18.885000 ;
        RECT 55.285000  8.935000 74.700000  9.005000 ;
        RECT 55.340000 18.745000 74.700000 18.815000 ;
        RECT 55.355000  9.005000 74.700000  9.075000 ;
        RECT 55.410000 18.675000 74.700000 18.745000 ;
        RECT 55.425000  9.075000 74.700000  9.145000 ;
        RECT 55.480000 18.605000 74.700000 18.675000 ;
        RECT 55.495000  9.145000 74.700000  9.215000 ;
        RECT 55.550000 18.535000 74.700000 18.605000 ;
        RECT 55.565000  9.215000 74.700000  9.285000 ;
        RECT 55.620000 18.465000 74.700000 18.535000 ;
        RECT 55.635000  9.285000 74.700000  9.355000 ;
        RECT 55.690000 18.395000 74.700000 18.465000 ;
        RECT 55.705000  9.355000 74.700000  9.425000 ;
        RECT 55.760000 18.325000 74.700000 18.395000 ;
        RECT 55.775000  9.425000 74.700000  9.495000 ;
        RECT 55.830000 18.255000 74.700000 18.325000 ;
        RECT 55.845000  9.495000 74.700000  9.565000 ;
        RECT 55.900000 18.185000 74.700000 18.255000 ;
        RECT 55.915000  9.565000 74.700000  9.635000 ;
        RECT 55.970000 18.115000 74.700000 18.185000 ;
        RECT 55.985000  9.635000 74.700000  9.705000 ;
        RECT 56.040000 18.045000 74.700000 18.115000 ;
        RECT 56.055000  9.705000 74.700000  9.775000 ;
        RECT 56.110000 17.975000 74.700000 18.045000 ;
        RECT 56.125000  9.775000 74.700000  9.845000 ;
        RECT 56.180000 17.905000 74.700000 17.975000 ;
        RECT 56.195000  9.845000 74.700000  9.915000 ;
        RECT 56.250000  9.915000 74.700000  9.970000 ;
        RECT 56.250000  9.970000 74.700000 17.835000 ;
        RECT 56.250000 17.835000 74.700000 17.905000 ;
        RECT 62.325000 21.695000 74.700000 21.765000 ;
        RECT 62.395000 21.765000 74.700000 21.835000 ;
        RECT 62.465000 21.835000 74.700000 21.905000 ;
        RECT 62.535000 21.905000 74.700000 21.975000 ;
        RECT 62.605000 21.975000 74.700000 22.045000 ;
        RECT 62.675000 22.045000 74.700000 22.115000 ;
        RECT 62.745000 22.115000 74.700000 22.185000 ;
        RECT 62.815000 22.185000 74.700000 22.255000 ;
        RECT 62.885000 22.255000 74.700000 22.325000 ;
        RECT 62.955000 22.325000 74.700000 22.395000 ;
        RECT 63.025000 22.395000 74.700000 22.465000 ;
        RECT 63.095000 22.465000 74.700000 22.535000 ;
        RECT 63.165000 22.535000 74.700000 22.605000 ;
        RECT 63.235000 22.605000 74.700000 22.675000 ;
        RECT 63.305000 22.675000 74.700000 22.745000 ;
        RECT 63.375000 22.745000 74.700000 22.815000 ;
        RECT 63.445000 22.815000 74.700000 22.885000 ;
        RECT 63.515000 22.885000 74.700000 22.955000 ;
        RECT 63.585000 22.955000 74.700000 23.025000 ;
        RECT 63.655000 23.025000 74.700000 23.095000 ;
        RECT 63.725000 23.095000 74.700000 23.165000 ;
        RECT 63.795000 23.165000 74.700000 23.235000 ;
        RECT 63.865000 23.235000 74.700000 23.305000 ;
        RECT 63.935000 23.305000 74.700000 23.375000 ;
        RECT 64.005000 23.375000 74.700000 23.445000 ;
        RECT 64.075000 23.445000 74.700000 23.515000 ;
        RECT 64.145000 23.515000 74.700000 23.585000 ;
        RECT 64.215000 23.585000 74.700000 23.655000 ;
        RECT 64.285000 23.655000 74.700000 23.725000 ;
        RECT 64.355000 23.725000 74.700000 23.795000 ;
        RECT 64.425000 23.795000 74.700000 23.865000 ;
        RECT 64.495000 23.865000 74.700000 23.935000 ;
        RECT 64.565000 23.935000 74.700000 24.005000 ;
        RECT 64.635000 24.005000 74.700000 24.075000 ;
        RECT 64.705000 24.075000 74.700000 24.145000 ;
        RECT 64.775000 24.145000 74.700000 24.215000 ;
        RECT 64.845000 24.215000 74.700000 24.285000 ;
        RECT 64.880000 31.000000 74.700000 31.010000 ;
        RECT 64.915000 24.285000 74.700000 24.355000 ;
        RECT 64.950000 30.930000 74.700000 31.000000 ;
        RECT 64.950000 40.985000 74.700000 40.990000 ;
        RECT 64.950000 51.005000 74.700000 51.010000 ;
        RECT 64.985000 24.355000 74.700000 24.425000 ;
        RECT 65.015000 60.920000 74.700000 60.990000 ;
        RECT 65.015000 63.630000 74.700000 63.700000 ;
        RECT 65.015000 70.920000 74.700000 70.990000 ;
        RECT 65.020000 30.860000 74.700000 30.930000 ;
        RECT 65.020000 40.915000 74.700000 40.985000 ;
        RECT 65.020000 50.935000 74.700000 51.005000 ;
        RECT 65.030000 33.650000 74.700000 33.720000 ;
        RECT 65.030000 43.630000 74.700000 43.700000 ;
        RECT 65.030000 53.650000 74.700000 53.720000 ;
        RECT 65.055000 24.425000 74.700000 24.495000 ;
        RECT 65.085000 60.850000 74.700000 60.920000 ;
        RECT 65.085000 63.700000 74.700000 63.770000 ;
        RECT 65.085000 70.850000 74.700000 70.920000 ;
        RECT 65.090000 30.790000 74.700000 30.860000 ;
        RECT 65.090000 40.845000 74.700000 40.915000 ;
        RECT 65.090000 50.865000 74.700000 50.935000 ;
        RECT 65.100000 33.720000 74.700000 33.790000 ;
        RECT 65.100000 43.700000 74.700000 43.770000 ;
        RECT 65.100000 53.720000 74.700000 53.790000 ;
        RECT 65.125000 24.495000 74.700000 24.565000 ;
        RECT 65.155000 60.780000 74.700000 60.850000 ;
        RECT 65.155000 63.770000 74.700000 63.840000 ;
        RECT 65.155000 70.780000 74.700000 70.850000 ;
        RECT 65.160000 30.720000 74.700000 30.790000 ;
        RECT 65.160000 40.775000 74.700000 40.845000 ;
        RECT 65.160000 50.795000 74.700000 50.865000 ;
        RECT 65.170000 33.790000 74.700000 33.860000 ;
        RECT 65.170000 43.770000 74.700000 43.840000 ;
        RECT 65.170000 53.790000 74.700000 53.860000 ;
        RECT 65.195000 24.565000 74.700000 24.635000 ;
        RECT 65.225000 60.710000 74.700000 60.780000 ;
        RECT 65.225000 63.840000 74.700000 63.910000 ;
        RECT 65.225000 70.710000 74.700000 70.780000 ;
        RECT 65.230000 30.650000 74.700000 30.720000 ;
        RECT 65.230000 40.705000 74.700000 40.775000 ;
        RECT 65.230000 50.725000 74.700000 50.795000 ;
        RECT 65.240000 33.860000 74.700000 33.930000 ;
        RECT 65.240000 43.840000 74.700000 43.910000 ;
        RECT 65.240000 53.860000 74.700000 53.930000 ;
        RECT 65.265000 24.635000 74.700000 24.705000 ;
        RECT 65.270000 73.630000 68.740000 73.700000 ;
        RECT 65.295000 60.640000 74.700000 60.710000 ;
        RECT 65.295000 63.910000 74.700000 63.980000 ;
        RECT 65.295000 70.640000 74.700000 70.710000 ;
        RECT 65.300000 30.580000 74.700000 30.650000 ;
        RECT 65.300000 40.635000 74.700000 40.705000 ;
        RECT 65.300000 50.655000 74.700000 50.725000 ;
        RECT 65.310000 33.930000 74.700000 34.000000 ;
        RECT 65.310000 43.910000 74.700000 43.980000 ;
        RECT 65.310000 53.930000 74.700000 54.000000 ;
        RECT 65.335000 24.705000 74.700000 24.775000 ;
        RECT 65.340000 73.700000 68.670000 73.770000 ;
        RECT 65.365000 60.570000 74.700000 60.640000 ;
        RECT 65.365000 63.980000 74.700000 64.050000 ;
        RECT 65.365000 70.570000 74.700000 70.640000 ;
        RECT 65.370000 30.510000 74.700000 30.580000 ;
        RECT 65.370000 40.565000 74.700000 40.635000 ;
        RECT 65.370000 50.585000 74.700000 50.655000 ;
        RECT 65.380000 34.000000 74.700000 34.070000 ;
        RECT 65.380000 43.980000 74.700000 44.050000 ;
        RECT 65.380000 54.000000 74.700000 54.070000 ;
        RECT 65.405000 24.775000 74.700000 24.845000 ;
        RECT 65.410000 73.770000 68.600000 73.840000 ;
        RECT 65.435000 60.500000 74.700000 60.570000 ;
        RECT 65.435000 64.050000 74.700000 64.120000 ;
        RECT 65.435000 70.500000 74.700000 70.570000 ;
        RECT 65.440000 30.440000 74.700000 30.510000 ;
        RECT 65.440000 40.495000 74.700000 40.565000 ;
        RECT 65.440000 50.515000 74.700000 50.585000 ;
        RECT 65.450000 34.070000 74.700000 34.140000 ;
        RECT 65.450000 44.050000 74.700000 44.120000 ;
        RECT 65.450000 54.070000 74.700000 54.140000 ;
        RECT 65.475000 24.845000 74.700000 24.915000 ;
        RECT 65.480000 73.840000 68.530000 73.910000 ;
        RECT 65.505000 60.430000 74.700000 60.500000 ;
        RECT 65.505000 64.120000 74.700000 64.190000 ;
        RECT 65.505000 70.430000 74.700000 70.500000 ;
        RECT 65.510000 30.370000 74.700000 30.440000 ;
        RECT 65.510000 40.425000 74.700000 40.495000 ;
        RECT 65.510000 50.445000 74.700000 50.515000 ;
        RECT 65.520000 34.140000 74.700000 34.210000 ;
        RECT 65.520000 44.120000 74.700000 44.190000 ;
        RECT 65.520000 54.140000 74.700000 54.210000 ;
        RECT 65.545000 24.915000 74.700000 24.985000 ;
        RECT 65.550000 73.910000 68.460000 73.980000 ;
        RECT 65.575000 60.360000 74.700000 60.430000 ;
        RECT 65.575000 64.190000 74.700000 64.260000 ;
        RECT 65.575000 70.360000 74.700000 70.430000 ;
        RECT 65.580000 30.300000 74.700000 30.370000 ;
        RECT 65.580000 40.355000 74.700000 40.425000 ;
        RECT 65.580000 50.375000 74.700000 50.445000 ;
        RECT 65.590000 34.210000 74.700000 34.280000 ;
        RECT 65.590000 44.190000 74.700000 44.260000 ;
        RECT 65.590000 54.210000 74.700000 54.280000 ;
        RECT 65.615000 24.985000 74.700000 25.055000 ;
        RECT 65.620000 73.980000 68.390000 74.050000 ;
        RECT 65.645000 60.290000 74.700000 60.360000 ;
        RECT 65.645000 64.260000 74.700000 64.330000 ;
        RECT 65.645000 70.290000 74.700000 70.360000 ;
        RECT 65.650000 30.230000 74.700000 30.300000 ;
        RECT 65.650000 40.285000 74.700000 40.355000 ;
        RECT 65.650000 50.305000 74.700000 50.375000 ;
        RECT 65.660000 34.280000 74.700000 34.350000 ;
        RECT 65.660000 44.260000 74.700000 44.330000 ;
        RECT 65.660000 54.280000 74.700000 54.350000 ;
        RECT 65.685000 25.055000 74.700000 25.125000 ;
        RECT 65.690000 74.050000 68.320000 74.120000 ;
        RECT 65.715000 60.220000 74.700000 60.290000 ;
        RECT 65.715000 64.330000 74.700000 64.400000 ;
        RECT 65.715000 70.220000 74.700000 70.290000 ;
        RECT 65.720000 30.160000 74.700000 30.230000 ;
        RECT 65.720000 40.215000 74.700000 40.285000 ;
        RECT 65.720000 50.235000 74.700000 50.305000 ;
        RECT 65.730000 34.350000 74.700000 34.420000 ;
        RECT 65.730000 44.330000 74.700000 44.400000 ;
        RECT 65.730000 54.350000 74.700000 54.420000 ;
        RECT 65.755000 25.125000 74.700000 25.195000 ;
        RECT 65.760000 74.120000 68.250000 74.190000 ;
        RECT 65.785000 60.150000 74.700000 60.220000 ;
        RECT 65.785000 64.400000 74.700000 64.470000 ;
        RECT 65.785000 70.150000 74.700000 70.220000 ;
        RECT 65.790000 30.090000 74.700000 30.160000 ;
        RECT 65.790000 40.145000 74.700000 40.215000 ;
        RECT 65.790000 50.165000 74.700000 50.235000 ;
        RECT 65.800000 34.420000 74.700000 34.490000 ;
        RECT 65.800000 44.400000 74.700000 44.470000 ;
        RECT 65.800000 54.420000 74.700000 54.490000 ;
        RECT 65.825000 25.195000 74.700000 25.265000 ;
        RECT 65.830000 74.190000 68.180000 74.260000 ;
        RECT 65.855000 60.080000 74.700000 60.150000 ;
        RECT 65.855000 64.470000 74.700000 64.540000 ;
        RECT 65.855000 70.080000 74.700000 70.150000 ;
        RECT 65.860000 30.020000 74.700000 30.090000 ;
        RECT 65.860000 40.075000 74.700000 40.145000 ;
        RECT 65.860000 50.095000 74.700000 50.165000 ;
        RECT 65.870000 34.490000 74.700000 34.560000 ;
        RECT 65.870000 44.470000 74.700000 44.540000 ;
        RECT 65.870000 54.490000 74.700000 54.560000 ;
        RECT 65.895000 25.265000 74.700000 25.335000 ;
        RECT 65.900000 74.260000 68.110000 74.330000 ;
        RECT 65.925000 60.010000 74.700000 60.080000 ;
        RECT 65.925000 64.540000 74.700000 64.610000 ;
        RECT 65.925000 70.010000 74.700000 70.080000 ;
        RECT 65.930000 29.950000 74.700000 30.020000 ;
        RECT 65.930000 40.005000 74.700000 40.075000 ;
        RECT 65.930000 50.025000 74.700000 50.095000 ;
        RECT 65.940000 34.560000 74.700000 34.630000 ;
        RECT 65.940000 44.540000 74.700000 44.610000 ;
        RECT 65.940000 54.560000 74.700000 54.630000 ;
        RECT 65.965000 25.335000 74.700000 25.405000 ;
        RECT 65.970000 74.330000 68.040000 74.400000 ;
        RECT 65.995000 54.630000 74.700000 54.685000 ;
        RECT 65.995000 54.685000 74.700000 59.940000 ;
        RECT 65.995000 59.940000 74.700000 60.010000 ;
        RECT 65.995000 64.610000 74.700000 64.680000 ;
        RECT 65.995000 64.680000 74.700000 69.940000 ;
        RECT 65.995000 69.940000 74.700000 70.010000 ;
        RECT 66.000000 25.405000 74.700000 25.440000 ;
        RECT 66.000000 25.440000 74.700000 29.880000 ;
        RECT 66.000000 29.880000 74.700000 29.950000 ;
        RECT 66.000000 34.630000 74.700000 34.690000 ;
        RECT 66.000000 34.690000 74.700000 39.935000 ;
        RECT 66.000000 39.935000 74.700000 40.005000 ;
        RECT 66.000000 44.610000 74.700000 44.670000 ;
        RECT 66.000000 44.670000 74.700000 49.955000 ;
        RECT 66.000000 49.955000 74.700000 50.025000 ;
        RECT 66.000000 74.400000 68.010000 74.430000 ;
        RECT 66.000000 74.430000 68.010000 98.560000 ;
    END
  END SRC_BDY_LVC2
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  0.240000  17.210000  2.995000  19.200000 ;
      RECT  1.350000   1.020000  7.110000   1.190000 ;
      RECT  1.350000   1.190000  1.520000  17.040000 ;
      RECT  1.350000  17.040000  7.110000  17.210000 ;
      RECT  1.760000  19.630000  9.385000  20.140000 ;
      RECT  1.760000  20.140000  2.685000  23.060000 ;
      RECT  1.845000   3.220000  2.015000   8.960000 ;
      RECT  1.845000   9.710000  2.015000  16.610000 ;
      RECT  2.070000   1.610000  6.390000   1.780000 ;
      RECT  2.070000   9.260000  6.390000   9.430000 ;
      RECT  2.305000   2.490000  2.475000   8.960000 ;
      RECT  2.305000  10.140000  2.475000  15.440000 ;
      RECT  2.765000   3.220000  2.935000   8.960000 ;
      RECT  2.765000   9.710000  2.935000  16.610000 ;
      RECT  3.225000   2.490000  3.395000   8.960000 ;
      RECT  3.225000  10.140000  3.395000  15.440000 ;
      RECT  3.685000   3.220000  3.855000   8.960000 ;
      RECT  3.685000   9.710000  3.855000  16.610000 ;
      RECT  4.145000   2.490000  4.315000   8.960000 ;
      RECT  4.145000  10.140000  4.315000  15.440000 ;
      RECT  4.605000   3.220000  4.775000   8.960000 ;
      RECT  4.605000   9.710000  4.775000  16.610000 ;
      RECT  4.975000  22.290000 10.650000  23.010000 ;
      RECT  5.065000   2.490000  5.235000   8.960000 ;
      RECT  5.065000  10.140000  5.235000  15.440000 ;
      RECT  5.525000   3.220000  5.695000   8.960000 ;
      RECT  5.525000   9.710000  5.695000  16.610000 ;
      RECT  5.890000  23.010000 10.650000  23.015000 ;
      RECT  5.985000   2.490000  6.155000   8.960000 ;
      RECT  5.985000  10.140000  6.155000  15.440000 ;
      RECT  6.445000   2.060000  6.615000   8.960000 ;
      RECT  6.445000   9.710000  6.615000  16.610000 ;
      RECT  6.940000   1.190000  7.110000  17.040000 ;
      RECT  8.340000 196.360000  8.670000 196.420000 ;
      RECT  8.345000   1.410000 16.655000  18.350000 ;
      RECT  8.420000 195.890000  8.590000 196.360000 ;
      RECT  9.155000 106.965000 10.280000 196.850000 ;
      RECT  9.155000 196.850000 69.720000 197.380000 ;
      RECT  9.185000  23.825000 69.720000  24.355000 ;
      RECT  9.185000  24.355000 10.280000  82.980000 ;
      RECT  9.185000  82.980000 21.740000  83.150000 ;
      RECT  9.185000  83.150000 10.280000  99.490000 ;
      RECT  9.730000  99.490000 10.280000 106.965000 ;
      RECT 10.920000  83.820000 11.830000  84.585000 ;
      RECT 11.065000 168.280000 12.050000 194.935000 ;
      RECT 11.065000 194.935000 68.495000 195.885000 ;
      RECT 11.095000 144.465000 11.795000 144.635000 ;
      RECT 11.095000 144.635000 21.320000 145.145000 ;
      RECT 11.095000 145.145000 12.050000 168.280000 ;
      RECT 11.275000  25.065000 68.140000  26.075000 ;
      RECT 11.275000  26.075000 12.220000  34.040000 ;
      RECT 11.275000  36.745000 12.220000  43.620000 ;
      RECT 11.275000  46.905000 12.220000  81.705000 ;
      RECT 11.275000  81.705000 23.280000  82.180000 ;
      RECT 11.275000  82.180000 68.140000  82.215000 ;
      RECT 11.370000  34.040000 12.220000  36.745000 ;
      RECT 11.370000  43.620000 12.220000  46.905000 ;
      RECT 12.405000 184.140000 66.575000 186.620000 ;
      RECT 12.430000 184.100000 66.575000 184.140000 ;
      RECT 12.750000  75.785000 12.920000  80.300000 ;
      RECT 12.975000  81.045000 66.655000  81.215000 ;
      RECT 13.060000  44.100000 65.590000  46.620000 ;
      RECT 13.060000  64.100000 65.590000  66.620000 ;
      RECT 13.190000  34.100000 65.590000  36.620000 ;
      RECT 13.190000  54.100000 65.590000  56.620000 ;
      RECT 13.335000 174.100000 65.590000 176.620000 ;
      RECT 13.365000 145.615000 14.305000 145.620000 ;
      RECT 13.365000 145.620000 65.590000 146.620000 ;
      RECT 13.365000 154.100000 65.590000 156.620000 ;
      RECT 13.365000 164.100000 65.590000 166.620000 ;
      RECT 13.395000  26.900000 13.925000  33.570000 ;
      RECT 13.395000  36.900000 13.925000  43.570000 ;
      RECT 13.395000  46.900000 13.925000  53.570000 ;
      RECT 13.395000  56.900000 13.925000  63.570000 ;
      RECT 13.395000  66.900000 13.925000  71.725000 ;
      RECT 13.395000 186.900000 13.925000 193.570000 ;
      RECT 14.360000 194.100000 65.590000 194.270000 ;
      RECT 14.780000  26.900000 15.310000  33.570000 ;
      RECT 14.780000  36.900000 15.310000  43.570000 ;
      RECT 14.780000  46.900000 15.310000  53.570000 ;
      RECT 14.780000  56.900000 15.310000  63.570000 ;
      RECT 14.780000  66.900000 15.310000  71.725000 ;
      RECT 14.780000 186.900000 15.310000 193.570000 ;
      RECT 14.790000  26.840000 15.300000  26.900000 ;
      RECT 14.790000  33.570000 15.300000  33.630000 ;
      RECT 14.790000  36.840000 15.300000  36.900000 ;
      RECT 14.790000  43.570000 15.300000  43.630000 ;
      RECT 14.790000  46.840000 15.300000  46.900000 ;
      RECT 14.790000  53.570000 15.300000  53.630000 ;
      RECT 14.790000  56.840000 15.300000  56.900000 ;
      RECT 14.790000  63.570000 15.300000  63.630000 ;
      RECT 14.790000  66.840000 15.300000  66.900000 ;
      RECT 14.790000 186.840000 15.300000 186.900000 ;
      RECT 14.790000 193.570000 15.300000 193.630000 ;
      RECT 15.865000 146.900000 16.395000 153.570000 ;
      RECT 15.865000 156.900000 16.395000 163.570000 ;
      RECT 15.865000 166.900000 16.395000 173.570000 ;
      RECT 16.165000  26.900000 16.695000  33.570000 ;
      RECT 16.165000  36.900000 16.695000  43.570000 ;
      RECT 16.165000  46.900000 16.695000  53.570000 ;
      RECT 16.165000  56.900000 16.695000  63.570000 ;
      RECT 16.165000  66.900000 16.695000  71.725000 ;
      RECT 16.165000 176.900000 16.695000 183.570000 ;
      RECT 16.165000 186.900000 16.695000 193.570000 ;
      RECT 17.000000  17.580000 56.200000  18.350000 ;
      RECT 17.030000  75.785000 17.200000  80.300000 ;
      RECT 17.550000  26.900000 18.080000  33.570000 ;
      RECT 17.550000  36.900000 18.080000  43.570000 ;
      RECT 17.550000  46.900000 18.080000  53.570000 ;
      RECT 17.550000  56.900000 18.080000  63.570000 ;
      RECT 17.550000  66.900000 18.080000  71.725000 ;
      RECT 17.550000 176.900000 18.080000 183.570000 ;
      RECT 17.550000 186.900000 18.080000 193.570000 ;
      RECT 17.560000  26.840000 18.070000  26.900000 ;
      RECT 17.560000  33.570000 18.070000  33.630000 ;
      RECT 17.560000  36.840000 18.070000  36.900000 ;
      RECT 17.560000  43.570000 18.070000  43.630000 ;
      RECT 17.560000  46.840000 18.070000  46.900000 ;
      RECT 17.560000  53.570000 18.070000  53.630000 ;
      RECT 17.560000  56.840000 18.070000  56.900000 ;
      RECT 17.560000  63.570000 18.070000  63.630000 ;
      RECT 17.560000  66.840000 18.070000  66.900000 ;
      RECT 17.560000 176.840000 18.070000 176.900000 ;
      RECT 17.560000 183.570000 18.070000 183.630000 ;
      RECT 17.560000 186.840000 18.070000 186.900000 ;
      RECT 17.560000 193.570000 18.070000 193.630000 ;
      RECT 17.955000 146.900000 18.485000 153.570000 ;
      RECT 17.955000 156.900000 18.485000 163.570000 ;
      RECT 17.955000 166.900000 18.485000 173.570000 ;
      RECT 17.965000 146.840000 18.475000 146.900000 ;
      RECT 17.965000 153.570000 18.475000 153.630000 ;
      RECT 17.965000 156.840000 18.475000 156.900000 ;
      RECT 17.965000 163.570000 18.475000 163.630000 ;
      RECT 17.965000 166.840000 18.475000 166.900000 ;
      RECT 17.965000 173.570000 18.475000 173.630000 ;
      RECT 18.935000  26.900000 19.465000  33.570000 ;
      RECT 18.935000  36.900000 19.465000  43.570000 ;
      RECT 18.935000  46.900000 19.465000  53.570000 ;
      RECT 18.935000  56.900000 19.465000  63.570000 ;
      RECT 18.935000  66.900000 19.465000  71.725000 ;
      RECT 18.935000 176.900000 19.465000 183.570000 ;
      RECT 18.935000 186.900000 19.465000 193.570000 ;
      RECT 19.495000  83.820000 20.405000  84.585000 ;
      RECT 20.045000 146.900000 20.575000 153.570000 ;
      RECT 20.045000 156.900000 20.575000 163.570000 ;
      RECT 20.045000 166.900000 20.575000 173.570000 ;
      RECT 20.320000  26.900000 20.850000  33.570000 ;
      RECT 20.320000  36.900000 20.850000  43.570000 ;
      RECT 20.320000  46.900000 20.850000  53.570000 ;
      RECT 20.320000  56.900000 20.850000  63.570000 ;
      RECT 20.320000  66.900000 20.850000  71.725000 ;
      RECT 20.320000 176.900000 20.850000 183.570000 ;
      RECT 20.320000 186.900000 20.850000 193.570000 ;
      RECT 20.330000  26.840000 20.840000  26.900000 ;
      RECT 20.330000  33.570000 20.840000  33.630000 ;
      RECT 20.330000  36.840000 20.840000  36.900000 ;
      RECT 20.330000  43.570000 20.840000  43.630000 ;
      RECT 20.330000  46.840000 20.840000  46.900000 ;
      RECT 20.330000  53.570000 20.840000  53.630000 ;
      RECT 20.330000  56.840000 20.840000  56.900000 ;
      RECT 20.330000  63.570000 20.840000  63.630000 ;
      RECT 20.330000  66.840000 20.840000  66.900000 ;
      RECT 20.330000 176.840000 20.840000 176.900000 ;
      RECT 20.330000 183.570000 20.840000 183.630000 ;
      RECT 20.330000 186.840000 20.840000 186.900000 ;
      RECT 20.330000 193.570000 20.840000 193.630000 ;
      RECT 20.810000 100.865000 68.495000 101.035000 ;
      RECT 20.810000 101.035000 21.320000 109.275000 ;
      RECT 20.810000 109.275000 68.495000 109.445000 ;
      RECT 20.810000 109.445000 21.320000 117.770000 ;
      RECT 20.810000 117.770000 68.495000 117.940000 ;
      RECT 20.810000 117.940000 21.320000 144.635000 ;
      RECT 21.570000  83.150000 21.740000  99.925000 ;
      RECT 21.570000  99.925000 69.720000 100.095000 ;
      RECT 21.660000 128.010000 65.590000 128.515000 ;
      RECT 21.690000 134.100000 65.590000 136.620000 ;
      RECT 21.705000  26.900000 22.235000  33.570000 ;
      RECT 21.705000  36.900000 22.235000  43.570000 ;
      RECT 21.705000  46.900000 22.235000  53.570000 ;
      RECT 21.705000  56.900000 22.235000  63.570000 ;
      RECT 21.705000  66.900000 22.235000  71.725000 ;
      RECT 21.705000 176.900000 22.235000 183.570000 ;
      RECT 21.705000 186.900000 22.235000 193.570000 ;
      RECT 22.135000 146.900000 22.665000 153.570000 ;
      RECT 22.135000 156.900000 22.665000 163.570000 ;
      RECT 22.135000 166.900000 22.665000 173.570000 ;
      RECT 22.145000 146.840000 22.655000 146.900000 ;
      RECT 22.145000 153.570000 22.655000 153.630000 ;
      RECT 22.145000 156.840000 22.655000 156.900000 ;
      RECT 22.145000 163.570000 22.655000 163.630000 ;
      RECT 22.145000 166.840000 22.655000 166.900000 ;
      RECT 22.145000 173.570000 22.655000 173.630000 ;
      RECT 22.430000  82.215000 68.140000  82.350000 ;
      RECT 22.430000  82.350000 23.280000  90.675000 ;
      RECT 22.430000  90.675000 68.140000  90.845000 ;
      RECT 22.430000  90.845000 23.280000  97.890000 ;
      RECT 22.600000  97.890000 23.110000  98.990000 ;
      RECT 22.600000  98.990000 68.140000  99.160000 ;
      RECT 23.090000  26.900000 23.620000  33.570000 ;
      RECT 23.090000  36.900000 23.620000  43.570000 ;
      RECT 23.090000  46.900000 23.620000  53.570000 ;
      RECT 23.090000  56.900000 23.620000  63.570000 ;
      RECT 23.090000  66.900000 23.620000  71.725000 ;
      RECT 23.090000 176.900000 23.620000 183.570000 ;
      RECT 23.090000 186.900000 23.620000 193.570000 ;
      RECT 23.100000  26.840000 23.610000  26.900000 ;
      RECT 23.100000  33.570000 23.610000  33.630000 ;
      RECT 23.100000  36.840000 23.610000  36.900000 ;
      RECT 23.100000  43.570000 23.610000  43.630000 ;
      RECT 23.100000  46.840000 23.610000  46.900000 ;
      RECT 23.100000  53.570000 23.610000  53.630000 ;
      RECT 23.100000  56.840000 23.610000  56.900000 ;
      RECT 23.100000  63.570000 23.610000  63.630000 ;
      RECT 23.100000  66.840000 23.610000  66.900000 ;
      RECT 23.100000 176.840000 23.610000 176.900000 ;
      RECT 23.100000 183.570000 23.610000 183.630000 ;
      RECT 23.100000 186.840000 23.610000 186.900000 ;
      RECT 23.100000 193.570000 23.610000 193.630000 ;
      RECT 23.405000 144.100000 65.590000 145.620000 ;
      RECT 23.635000 101.385000 24.045000 108.175000 ;
      RECT 23.635000 109.880000 24.045000 115.550000 ;
      RECT 23.635000 120.080000 24.045000 125.295000 ;
      RECT 23.685000  82.785000 24.215000  89.575000 ;
      RECT 23.685000  91.280000 24.215000  98.070000 ;
      RECT 23.805000 115.550000 24.045000 116.670000 ;
      RECT 23.805000 118.955000 24.045000 120.080000 ;
      RECT 23.805000 125.295000 24.045000 125.745000 ;
      RECT 24.225000 128.730000 24.755000 133.760000 ;
      RECT 24.225000 136.900000 24.755000 143.570000 ;
      RECT 24.225000 146.900000 24.755000 153.570000 ;
      RECT 24.225000 156.900000 24.755000 163.570000 ;
      RECT 24.225000 166.900000 24.755000 173.570000 ;
      RECT 24.475000  26.900000 25.005000  33.570000 ;
      RECT 24.475000  36.900000 25.005000  43.570000 ;
      RECT 24.475000  46.900000 25.005000  53.570000 ;
      RECT 24.475000  56.900000 25.005000  63.570000 ;
      RECT 24.475000  66.900000 25.005000  71.725000 ;
      RECT 24.475000 176.900000 25.005000 183.570000 ;
      RECT 24.475000 186.900000 25.005000 193.570000 ;
      RECT 24.615000  90.045000 66.655000  90.215000 ;
      RECT 24.615000  98.540000 66.655000  98.710000 ;
      RECT 24.670000 108.645000 66.655000 108.815000 ;
      RECT 24.670000 117.140000 66.655000 117.310000 ;
      RECT 24.670000 118.315000 66.655000 118.485000 ;
      RECT 25.310000  75.785000 25.480000  80.300000 ;
      RECT 25.310000  82.915000 25.480000  89.020000 ;
      RECT 25.310000  91.930000 25.480000  96.925000 ;
      RECT 25.365000 101.385000 25.535000 106.255000 ;
      RECT 25.365000 110.450000 25.535000 115.330000 ;
      RECT 25.365000 120.080000 25.535000 124.860000 ;
      RECT 25.860000  26.900000 26.390000  33.570000 ;
      RECT 25.860000  36.900000 26.390000  43.570000 ;
      RECT 25.860000  46.900000 26.390000  53.570000 ;
      RECT 25.860000  56.900000 26.390000  63.570000 ;
      RECT 25.860000  66.900000 26.390000  71.725000 ;
      RECT 25.860000 176.900000 26.390000 183.570000 ;
      RECT 25.860000 186.900000 26.390000 193.570000 ;
      RECT 25.870000  26.840000 26.380000  26.900000 ;
      RECT 25.870000  33.570000 26.380000  33.630000 ;
      RECT 25.870000  36.840000 26.380000  36.900000 ;
      RECT 25.870000  43.570000 26.380000  43.630000 ;
      RECT 25.870000  46.840000 26.380000  46.900000 ;
      RECT 25.870000  53.570000 26.380000  53.630000 ;
      RECT 25.870000  56.840000 26.380000  56.900000 ;
      RECT 25.870000  63.570000 26.380000  63.630000 ;
      RECT 25.870000  66.840000 26.380000  66.900000 ;
      RECT 25.870000 176.840000 26.380000 176.900000 ;
      RECT 25.870000 183.570000 26.380000 183.630000 ;
      RECT 25.870000 186.840000 26.380000 186.900000 ;
      RECT 25.870000 193.570000 26.380000 193.630000 ;
      RECT 26.315000 128.730000 26.845000 133.715000 ;
      RECT 26.315000 136.900000 26.845000 143.570000 ;
      RECT 26.315000 146.900000 26.845000 153.570000 ;
      RECT 26.315000 156.900000 26.845000 163.570000 ;
      RECT 26.315000 166.900000 26.845000 173.570000 ;
      RECT 26.325000 136.840000 26.835000 136.900000 ;
      RECT 26.325000 143.570000 26.835000 143.630000 ;
      RECT 26.325000 146.840000 26.835000 146.900000 ;
      RECT 26.325000 153.570000 26.835000 153.630000 ;
      RECT 26.325000 156.840000 26.835000 156.900000 ;
      RECT 26.325000 163.570000 26.835000 163.630000 ;
      RECT 26.325000 166.840000 26.835000 166.900000 ;
      RECT 26.325000 173.570000 26.835000 173.630000 ;
      RECT 27.245000  26.900000 27.775000  33.570000 ;
      RECT 27.245000  36.900000 27.775000  43.570000 ;
      RECT 27.245000  46.900000 27.775000  53.570000 ;
      RECT 27.245000  56.900000 27.775000  63.570000 ;
      RECT 27.245000  66.900000 27.775000  71.725000 ;
      RECT 27.245000 176.900000 27.775000 183.570000 ;
      RECT 27.245000 186.900000 27.775000 193.570000 ;
      RECT 28.405000 128.860000 28.935000 133.760000 ;
      RECT 28.405000 136.900000 28.935000 143.570000 ;
      RECT 28.405000 146.900000 28.935000 153.570000 ;
      RECT 28.405000 156.900000 28.935000 163.570000 ;
      RECT 28.405000 166.900000 28.935000 173.570000 ;
      RECT 28.630000  26.900000 29.160000  33.570000 ;
      RECT 28.630000  36.900000 29.160000  43.570000 ;
      RECT 28.630000  46.900000 29.160000  53.570000 ;
      RECT 28.630000  56.900000 29.160000  63.570000 ;
      RECT 28.630000  66.900000 29.160000  71.725000 ;
      RECT 28.630000 176.900000 29.160000 183.570000 ;
      RECT 28.630000 186.900000 29.160000 193.570000 ;
      RECT 28.640000  26.840000 29.150000  26.900000 ;
      RECT 28.640000  33.570000 29.150000  33.630000 ;
      RECT 28.640000  36.840000 29.150000  36.900000 ;
      RECT 28.640000  43.570000 29.150000  43.630000 ;
      RECT 28.640000  46.840000 29.150000  46.900000 ;
      RECT 28.640000  53.570000 29.150000  53.630000 ;
      RECT 28.640000  56.840000 29.150000  56.900000 ;
      RECT 28.640000  63.570000 29.150000  63.630000 ;
      RECT 28.640000  66.840000 29.150000  66.900000 ;
      RECT 28.640000 176.840000 29.150000 176.900000 ;
      RECT 28.640000 183.570000 29.150000 183.630000 ;
      RECT 28.640000 186.840000 29.150000 186.900000 ;
      RECT 28.640000 193.570000 29.150000 193.630000 ;
      RECT 30.015000  26.900000 30.545000  33.570000 ;
      RECT 30.015000  36.900000 30.545000  43.570000 ;
      RECT 30.015000  46.900000 30.545000  53.570000 ;
      RECT 30.015000  56.900000 30.545000  63.570000 ;
      RECT 30.015000  66.900000 30.545000  71.725000 ;
      RECT 30.015000 176.900000 30.545000 183.570000 ;
      RECT 30.015000 186.900000 30.545000 193.570000 ;
      RECT 30.495000 128.730000 31.025000 133.715000 ;
      RECT 30.495000 136.900000 31.025000 143.570000 ;
      RECT 30.495000 146.900000 31.025000 153.570000 ;
      RECT 30.495000 156.900000 31.025000 163.570000 ;
      RECT 30.495000 166.900000 31.025000 173.570000 ;
      RECT 30.505000 136.840000 31.015000 136.900000 ;
      RECT 30.505000 143.570000 31.015000 143.630000 ;
      RECT 30.505000 146.840000 31.015000 146.900000 ;
      RECT 30.505000 153.570000 31.015000 153.630000 ;
      RECT 30.505000 156.840000 31.015000 156.900000 ;
      RECT 30.505000 163.570000 31.015000 163.630000 ;
      RECT 30.505000 166.840000 31.015000 166.900000 ;
      RECT 30.505000 173.570000 31.015000 173.630000 ;
      RECT 31.400000  26.900000 31.930000  33.570000 ;
      RECT 31.400000  36.900000 31.930000  43.570000 ;
      RECT 31.400000  46.900000 31.930000  53.570000 ;
      RECT 31.400000  56.900000 31.930000  63.570000 ;
      RECT 31.400000  66.900000 31.930000  71.725000 ;
      RECT 31.400000 176.900000 31.930000 183.570000 ;
      RECT 31.400000 186.900000 31.930000 193.570000 ;
      RECT 31.410000  26.840000 31.920000  26.900000 ;
      RECT 31.410000  33.570000 31.920000  33.630000 ;
      RECT 31.410000  36.840000 31.920000  36.900000 ;
      RECT 31.410000  43.570000 31.920000  43.630000 ;
      RECT 31.410000  46.840000 31.920000  46.900000 ;
      RECT 31.410000  53.570000 31.920000  53.630000 ;
      RECT 31.410000  56.840000 31.920000  56.900000 ;
      RECT 31.410000  63.570000 31.920000  63.630000 ;
      RECT 31.410000  66.840000 31.920000  66.900000 ;
      RECT 31.410000 176.840000 31.920000 176.900000 ;
      RECT 31.410000 183.570000 31.920000 183.630000 ;
      RECT 31.410000 186.840000 31.920000 186.900000 ;
      RECT 31.410000 193.570000 31.920000 193.630000 ;
      RECT 32.585000 128.730000 33.115000 133.755000 ;
      RECT 32.585000 136.900000 33.115000 143.570000 ;
      RECT 32.585000 146.900000 33.115000 153.570000 ;
      RECT 32.585000 156.900000 33.115000 163.570000 ;
      RECT 32.585000 166.900000 33.115000 173.570000 ;
      RECT 32.785000  26.900000 33.315000  33.570000 ;
      RECT 32.785000  36.900000 33.315000  43.570000 ;
      RECT 32.785000  46.900000 33.315000  53.570000 ;
      RECT 32.785000  56.900000 33.315000  63.570000 ;
      RECT 32.785000  66.900000 33.315000  71.725000 ;
      RECT 32.785000 176.900000 33.315000 183.570000 ;
      RECT 32.785000 186.900000 33.315000 193.570000 ;
      RECT 33.590000  75.785000 33.760000  80.300000 ;
      RECT 33.590000  82.915000 33.760000  89.020000 ;
      RECT 33.590000  91.930000 33.760000  96.925000 ;
      RECT 33.590000 101.385000 33.760000 106.255000 ;
      RECT 33.590000 110.450000 33.760000 115.270000 ;
      RECT 33.595000 120.080000 33.765000 124.860000 ;
      RECT 34.170000  26.900000 34.700000  33.570000 ;
      RECT 34.170000  36.900000 34.700000  43.570000 ;
      RECT 34.170000  46.900000 34.700000  53.570000 ;
      RECT 34.170000  56.900000 34.700000  63.570000 ;
      RECT 34.170000  66.900000 34.700000  71.725000 ;
      RECT 34.170000 176.900000 34.700000 183.570000 ;
      RECT 34.170000 186.900000 34.700000 193.570000 ;
      RECT 34.180000  26.840000 34.690000  26.900000 ;
      RECT 34.180000  33.570000 34.690000  33.630000 ;
      RECT 34.180000  36.840000 34.690000  36.900000 ;
      RECT 34.180000  43.570000 34.690000  43.630000 ;
      RECT 34.180000  46.840000 34.690000  46.900000 ;
      RECT 34.180000  53.570000 34.690000  53.630000 ;
      RECT 34.180000  56.840000 34.690000  56.900000 ;
      RECT 34.180000  63.570000 34.690000  63.630000 ;
      RECT 34.180000  66.840000 34.690000  66.900000 ;
      RECT 34.180000 176.840000 34.690000 176.900000 ;
      RECT 34.180000 183.570000 34.690000 183.630000 ;
      RECT 34.180000 186.840000 34.690000 186.900000 ;
      RECT 34.180000 193.570000 34.690000 193.630000 ;
      RECT 34.675000 128.730000 35.205000 133.840000 ;
      RECT 34.675000 136.900000 35.205000 143.570000 ;
      RECT 34.675000 146.900000 35.205000 153.570000 ;
      RECT 34.675000 156.900000 35.205000 163.570000 ;
      RECT 34.675000 166.900000 35.205000 173.570000 ;
      RECT 34.685000 136.840000 35.195000 136.900000 ;
      RECT 34.685000 143.570000 35.195000 143.630000 ;
      RECT 34.685000 146.840000 35.195000 146.900000 ;
      RECT 34.685000 153.570000 35.195000 153.630000 ;
      RECT 34.685000 156.840000 35.195000 156.900000 ;
      RECT 34.685000 163.570000 35.195000 163.630000 ;
      RECT 34.685000 166.840000 35.195000 166.900000 ;
      RECT 34.685000 173.570000 35.195000 173.630000 ;
      RECT 35.555000  26.900000 36.085000  33.570000 ;
      RECT 35.555000  36.900000 36.085000  43.570000 ;
      RECT 35.555000  46.900000 36.085000  53.570000 ;
      RECT 35.555000  56.900000 36.085000  63.570000 ;
      RECT 35.555000  66.900000 36.085000  71.725000 ;
      RECT 35.555000 176.900000 36.085000 183.570000 ;
      RECT 35.555000 186.900000 36.085000 193.570000 ;
      RECT 36.765000 128.730000 37.295000 133.755000 ;
      RECT 36.765000 136.900000 37.295000 143.570000 ;
      RECT 36.765000 146.900000 37.295000 153.570000 ;
      RECT 36.765000 156.900000 37.295000 163.570000 ;
      RECT 36.765000 166.900000 37.295000 173.570000 ;
      RECT 36.940000  26.900000 37.470000  33.570000 ;
      RECT 36.940000  36.900000 37.470000  43.570000 ;
      RECT 36.940000  46.900000 37.470000  53.570000 ;
      RECT 36.940000  56.900000 37.470000  63.570000 ;
      RECT 36.940000  66.900000 37.470000  71.725000 ;
      RECT 36.940000 176.900000 37.470000 183.570000 ;
      RECT 36.940000 186.900000 37.470000 193.570000 ;
      RECT 36.950000  26.840000 37.460000  26.900000 ;
      RECT 36.950000  33.570000 37.460000  33.630000 ;
      RECT 36.950000  36.840000 37.460000  36.900000 ;
      RECT 36.950000  43.570000 37.460000  43.630000 ;
      RECT 36.950000  46.840000 37.460000  46.900000 ;
      RECT 36.950000  53.570000 37.460000  53.630000 ;
      RECT 36.950000  56.840000 37.460000  56.900000 ;
      RECT 36.950000  63.570000 37.460000  63.630000 ;
      RECT 36.950000  66.840000 37.460000  66.900000 ;
      RECT 36.950000 176.840000 37.460000 176.900000 ;
      RECT 36.950000 183.570000 37.460000 183.630000 ;
      RECT 36.950000 186.840000 37.460000 186.900000 ;
      RECT 36.950000 193.570000 37.460000 193.630000 ;
      RECT 38.325000  26.900000 38.855000  33.570000 ;
      RECT 38.325000  36.900000 38.855000  43.570000 ;
      RECT 38.325000  46.900000 38.855000  53.570000 ;
      RECT 38.325000  56.900000 38.855000  63.570000 ;
      RECT 38.325000  66.900000 38.855000  71.725000 ;
      RECT 38.325000 176.900000 38.855000 183.570000 ;
      RECT 38.325000 186.900000 38.855000 193.570000 ;
      RECT 38.855000 128.730000 39.385000 133.925000 ;
      RECT 38.855000 136.900000 39.385000 143.570000 ;
      RECT 38.855000 146.900000 39.385000 153.570000 ;
      RECT 38.855000 156.900000 39.385000 163.570000 ;
      RECT 38.855000 166.900000 39.385000 173.570000 ;
      RECT 38.865000 136.840000 39.375000 136.900000 ;
      RECT 38.865000 143.570000 39.375000 143.630000 ;
      RECT 38.865000 146.840000 39.375000 146.900000 ;
      RECT 38.865000 153.570000 39.375000 153.630000 ;
      RECT 38.865000 156.840000 39.375000 156.900000 ;
      RECT 38.865000 163.570000 39.375000 163.630000 ;
      RECT 38.865000 166.840000 39.375000 166.900000 ;
      RECT 38.865000 173.570000 39.375000 173.630000 ;
      RECT 39.710000  26.900000 40.240000  33.570000 ;
      RECT 39.710000  36.900000 40.240000  43.570000 ;
      RECT 39.710000  46.900000 40.240000  53.570000 ;
      RECT 39.710000  56.900000 40.240000  63.570000 ;
      RECT 39.710000  66.900000 40.240000  71.725000 ;
      RECT 39.710000 176.900000 40.240000 183.570000 ;
      RECT 39.710000 186.900000 40.240000 193.570000 ;
      RECT 39.720000  26.840000 40.230000  26.900000 ;
      RECT 39.720000  33.570000 40.230000  33.630000 ;
      RECT 39.720000  36.840000 40.230000  36.900000 ;
      RECT 39.720000  43.570000 40.230000  43.630000 ;
      RECT 39.720000  46.840000 40.230000  46.900000 ;
      RECT 39.720000  53.570000 40.230000  53.630000 ;
      RECT 39.720000  56.840000 40.230000  56.900000 ;
      RECT 39.720000  63.570000 40.230000  63.630000 ;
      RECT 39.720000  66.840000 40.230000  66.900000 ;
      RECT 39.720000 176.840000 40.230000 176.900000 ;
      RECT 39.720000 183.570000 40.230000 183.630000 ;
      RECT 39.720000 186.840000 40.230000 186.900000 ;
      RECT 39.720000 193.570000 40.230000 193.630000 ;
      RECT 40.945000 128.730000 41.475000 133.755000 ;
      RECT 40.945000 136.900000 41.475000 143.570000 ;
      RECT 40.945000 146.900000 41.475000 153.570000 ;
      RECT 40.945000 156.900000 41.475000 163.570000 ;
      RECT 40.945000 166.900000 41.475000 173.570000 ;
      RECT 41.095000  26.900000 41.625000  33.570000 ;
      RECT 41.095000  36.900000 41.625000  43.570000 ;
      RECT 41.095000  46.900000 41.625000  53.570000 ;
      RECT 41.095000  56.900000 41.625000  63.570000 ;
      RECT 41.095000  66.900000 41.625000  71.725000 ;
      RECT 41.095000 176.900000 41.625000 183.570000 ;
      RECT 41.095000 186.900000 41.625000 193.570000 ;
      RECT 41.870000  75.785000 42.040000  80.300000 ;
      RECT 41.870000  82.915000 42.040000  89.020000 ;
      RECT 41.870000  91.930000 42.040000  96.925000 ;
      RECT 41.870000 101.385000 42.040000 106.255000 ;
      RECT 41.870000 110.450000 42.040000 115.270000 ;
      RECT 41.870000 120.080000 42.040000 124.860000 ;
      RECT 42.480000  26.900000 43.010000  33.570000 ;
      RECT 42.480000  36.900000 43.010000  43.570000 ;
      RECT 42.480000  46.900000 43.010000  53.570000 ;
      RECT 42.480000  56.900000 43.010000  63.570000 ;
      RECT 42.480000  66.900000 43.010000  71.725000 ;
      RECT 42.480000 176.900000 43.010000 183.570000 ;
      RECT 42.480000 186.900000 43.010000 193.570000 ;
      RECT 42.490000  26.840000 43.000000  26.900000 ;
      RECT 42.490000  33.570000 43.000000  33.630000 ;
      RECT 42.490000  36.840000 43.000000  36.900000 ;
      RECT 42.490000  43.570000 43.000000  43.630000 ;
      RECT 42.490000  46.840000 43.000000  46.900000 ;
      RECT 42.490000  53.570000 43.000000  53.630000 ;
      RECT 42.490000  56.840000 43.000000  56.900000 ;
      RECT 42.490000  63.570000 43.000000  63.630000 ;
      RECT 42.490000  66.840000 43.000000  66.900000 ;
      RECT 42.490000 176.840000 43.000000 176.900000 ;
      RECT 42.490000 183.570000 43.000000 183.630000 ;
      RECT 42.490000 186.840000 43.000000 186.900000 ;
      RECT 42.490000 193.570000 43.000000 193.630000 ;
      RECT 43.035000 128.730000 43.565000 133.925000 ;
      RECT 43.035000 136.900000 43.565000 143.570000 ;
      RECT 43.035000 146.900000 43.565000 153.570000 ;
      RECT 43.035000 156.900000 43.565000 163.570000 ;
      RECT 43.035000 166.900000 43.565000 173.570000 ;
      RECT 43.045000 136.840000 43.555000 136.900000 ;
      RECT 43.045000 143.570000 43.555000 143.630000 ;
      RECT 43.045000 146.840000 43.555000 146.900000 ;
      RECT 43.045000 153.570000 43.555000 153.630000 ;
      RECT 43.045000 156.840000 43.555000 156.900000 ;
      RECT 43.045000 163.570000 43.555000 163.630000 ;
      RECT 43.045000 166.840000 43.555000 166.900000 ;
      RECT 43.045000 173.570000 43.555000 173.630000 ;
      RECT 43.865000  26.900000 44.395000  33.570000 ;
      RECT 43.865000  36.900000 44.395000  43.570000 ;
      RECT 43.865000  46.900000 44.395000  53.570000 ;
      RECT 43.865000  56.900000 44.395000  63.570000 ;
      RECT 43.865000  66.900000 44.395000  71.725000 ;
      RECT 43.865000 176.900000 44.395000 183.570000 ;
      RECT 43.865000 186.900000 44.395000 193.570000 ;
      RECT 45.125000 128.730000 45.655000 133.755000 ;
      RECT 45.125000 136.900000 45.655000 143.570000 ;
      RECT 45.125000 146.900000 45.655000 153.570000 ;
      RECT 45.125000 156.900000 45.655000 163.570000 ;
      RECT 45.125000 166.900000 45.655000 173.570000 ;
      RECT 45.250000  26.900000 45.780000  33.570000 ;
      RECT 45.250000  36.900000 45.780000  43.570000 ;
      RECT 45.250000  46.900000 45.780000  53.570000 ;
      RECT 45.250000  56.900000 45.780000  63.570000 ;
      RECT 45.250000  66.900000 45.780000  71.725000 ;
      RECT 45.250000 176.900000 45.780000 183.570000 ;
      RECT 45.250000 186.900000 45.780000 193.570000 ;
      RECT 45.260000  26.840000 45.770000  26.900000 ;
      RECT 45.260000  33.570000 45.770000  33.630000 ;
      RECT 45.260000  36.840000 45.770000  36.900000 ;
      RECT 45.260000  43.570000 45.770000  43.630000 ;
      RECT 45.260000  46.840000 45.770000  46.900000 ;
      RECT 45.260000  53.570000 45.770000  53.630000 ;
      RECT 45.260000  56.840000 45.770000  56.900000 ;
      RECT 45.260000  63.570000 45.770000  63.630000 ;
      RECT 45.260000  66.840000 45.770000  66.900000 ;
      RECT 45.260000 176.840000 45.770000 176.900000 ;
      RECT 45.260000 183.570000 45.770000 183.630000 ;
      RECT 45.260000 186.840000 45.770000 186.900000 ;
      RECT 45.260000 193.570000 45.770000 193.630000 ;
      RECT 46.635000  26.900000 47.165000  33.570000 ;
      RECT 46.635000  36.900000 47.165000  43.570000 ;
      RECT 46.635000  46.900000 47.165000  53.570000 ;
      RECT 46.635000  56.900000 47.165000  63.570000 ;
      RECT 46.635000  66.900000 47.165000  71.725000 ;
      RECT 46.635000 176.900000 47.165000 183.570000 ;
      RECT 46.635000 186.900000 47.165000 193.570000 ;
      RECT 47.215000 128.730000 47.745000 133.925000 ;
      RECT 47.215000 136.900000 47.745000 143.570000 ;
      RECT 47.215000 146.900000 47.745000 153.570000 ;
      RECT 47.215000 156.900000 47.745000 163.570000 ;
      RECT 47.215000 166.900000 47.745000 173.570000 ;
      RECT 47.225000 136.840000 47.735000 136.900000 ;
      RECT 47.225000 143.570000 47.735000 143.630000 ;
      RECT 47.225000 146.840000 47.735000 146.900000 ;
      RECT 47.225000 153.570000 47.735000 153.630000 ;
      RECT 47.225000 156.840000 47.735000 156.900000 ;
      RECT 47.225000 163.570000 47.735000 163.630000 ;
      RECT 47.225000 166.840000 47.735000 166.900000 ;
      RECT 47.225000 173.570000 47.735000 173.630000 ;
      RECT 48.020000  26.900000 48.550000  33.570000 ;
      RECT 48.020000  36.900000 48.550000  43.570000 ;
      RECT 48.020000  46.900000 48.550000  53.570000 ;
      RECT 48.020000  56.900000 48.550000  63.570000 ;
      RECT 48.020000  66.900000 48.550000  71.725000 ;
      RECT 48.020000 176.900000 48.550000 183.570000 ;
      RECT 48.020000 186.900000 48.550000 193.570000 ;
      RECT 48.030000  26.840000 48.540000  26.900000 ;
      RECT 48.030000  33.570000 48.540000  33.630000 ;
      RECT 48.030000  36.840000 48.540000  36.900000 ;
      RECT 48.030000  43.570000 48.540000  43.630000 ;
      RECT 48.030000  46.840000 48.540000  46.900000 ;
      RECT 48.030000  53.570000 48.540000  53.630000 ;
      RECT 48.030000  56.840000 48.540000  56.900000 ;
      RECT 48.030000  63.570000 48.540000  63.630000 ;
      RECT 48.030000  66.840000 48.540000  66.900000 ;
      RECT 48.030000 176.840000 48.540000 176.900000 ;
      RECT 48.030000 183.570000 48.540000 183.630000 ;
      RECT 48.030000 186.840000 48.540000 186.900000 ;
      RECT 48.030000 193.570000 48.540000 193.630000 ;
      RECT 49.305000 128.730000 49.835000 133.755000 ;
      RECT 49.305000 136.900000 49.835000 143.570000 ;
      RECT 49.305000 146.900000 49.835000 153.570000 ;
      RECT 49.305000 156.900000 49.835000 163.570000 ;
      RECT 49.305000 166.900000 49.835000 173.570000 ;
      RECT 49.405000  26.900000 49.935000  33.570000 ;
      RECT 49.405000  36.900000 49.935000  43.570000 ;
      RECT 49.405000  46.900000 49.935000  53.570000 ;
      RECT 49.405000  56.900000 49.935000  63.570000 ;
      RECT 49.405000  66.900000 49.935000  71.725000 ;
      RECT 49.405000 176.900000 49.935000 183.570000 ;
      RECT 49.405000 186.900000 49.935000 193.570000 ;
      RECT 50.150000  75.785000 50.320000  80.300000 ;
      RECT 50.150000  82.915000 50.320000  89.020000 ;
      RECT 50.150000  91.930000 50.320000  96.925000 ;
      RECT 50.150000 101.385000 50.320000 106.255000 ;
      RECT 50.150000 110.450000 50.320000 115.270000 ;
      RECT 50.150000 120.080000 50.320000 124.860000 ;
      RECT 50.790000  26.900000 51.320000  33.570000 ;
      RECT 50.790000  36.900000 51.320000  43.570000 ;
      RECT 50.790000  46.900000 51.320000  53.570000 ;
      RECT 50.790000  56.900000 51.320000  63.570000 ;
      RECT 50.790000  66.900000 51.320000  71.725000 ;
      RECT 50.790000 176.900000 51.320000 183.570000 ;
      RECT 50.790000 186.900000 51.320000 193.570000 ;
      RECT 50.800000  26.840000 51.310000  26.900000 ;
      RECT 50.800000  33.570000 51.310000  33.630000 ;
      RECT 50.800000  36.840000 51.310000  36.900000 ;
      RECT 50.800000  43.570000 51.310000  43.630000 ;
      RECT 50.800000  46.840000 51.310000  46.900000 ;
      RECT 50.800000  53.570000 51.310000  53.630000 ;
      RECT 50.800000  56.840000 51.310000  56.900000 ;
      RECT 50.800000  63.570000 51.310000  63.630000 ;
      RECT 50.800000  66.840000 51.310000  66.900000 ;
      RECT 50.800000 176.840000 51.310000 176.900000 ;
      RECT 50.800000 183.570000 51.310000 183.630000 ;
      RECT 50.800000 186.840000 51.310000 186.900000 ;
      RECT 50.800000 193.570000 51.310000 193.630000 ;
      RECT 51.395000 128.730000 51.925000 133.925000 ;
      RECT 51.395000 136.900000 51.925000 143.570000 ;
      RECT 51.395000 146.900000 51.925000 153.570000 ;
      RECT 51.395000 156.900000 51.925000 163.570000 ;
      RECT 51.395000 166.900000 51.925000 173.570000 ;
      RECT 51.405000 136.840000 51.915000 136.900000 ;
      RECT 51.405000 143.570000 51.915000 143.630000 ;
      RECT 51.405000 146.840000 51.915000 146.900000 ;
      RECT 51.405000 153.570000 51.915000 153.630000 ;
      RECT 51.405000 156.840000 51.915000 156.900000 ;
      RECT 51.405000 163.570000 51.915000 163.630000 ;
      RECT 51.405000 166.840000 51.915000 166.900000 ;
      RECT 51.405000 173.570000 51.915000 173.630000 ;
      RECT 52.175000  26.900000 52.705000  33.570000 ;
      RECT 52.175000  36.900000 52.705000  43.570000 ;
      RECT 52.175000  46.900000 52.705000  53.570000 ;
      RECT 52.175000  56.900000 52.705000  63.570000 ;
      RECT 52.175000  66.900000 52.705000  71.725000 ;
      RECT 52.175000 176.900000 52.705000 183.570000 ;
      RECT 52.175000 186.900000 52.705000 193.570000 ;
      RECT 53.485000 128.730000 54.015000 133.755000 ;
      RECT 53.485000 136.900000 54.015000 143.570000 ;
      RECT 53.485000 146.900000 54.015000 153.570000 ;
      RECT 53.485000 156.900000 54.015000 163.570000 ;
      RECT 53.485000 166.900000 54.015000 173.570000 ;
      RECT 53.560000  26.900000 54.090000  33.570000 ;
      RECT 53.560000  36.900000 54.090000  43.570000 ;
      RECT 53.560000  46.900000 54.090000  53.570000 ;
      RECT 53.560000  56.900000 54.090000  63.570000 ;
      RECT 53.560000  66.900000 54.090000  71.725000 ;
      RECT 53.560000 176.900000 54.090000 183.570000 ;
      RECT 53.560000 186.900000 54.090000 193.570000 ;
      RECT 53.570000  26.840000 54.080000  26.900000 ;
      RECT 53.570000  33.570000 54.080000  33.630000 ;
      RECT 53.570000  36.840000 54.080000  36.900000 ;
      RECT 53.570000  43.570000 54.080000  43.630000 ;
      RECT 53.570000  46.840000 54.080000  46.900000 ;
      RECT 53.570000  53.570000 54.080000  53.630000 ;
      RECT 53.570000  56.840000 54.080000  56.900000 ;
      RECT 53.570000  63.570000 54.080000  63.630000 ;
      RECT 53.570000  66.840000 54.080000  66.900000 ;
      RECT 53.570000 176.840000 54.080000 176.900000 ;
      RECT 53.570000 183.570000 54.080000 183.630000 ;
      RECT 53.570000 186.840000 54.080000 186.900000 ;
      RECT 53.570000 193.570000 54.080000 193.630000 ;
      RECT 54.945000  26.900000 55.475000  33.570000 ;
      RECT 54.945000  36.900000 55.475000  43.570000 ;
      RECT 54.945000  46.900000 55.475000  53.570000 ;
      RECT 54.945000  56.900000 55.475000  63.570000 ;
      RECT 54.945000  66.900000 55.475000  71.725000 ;
      RECT 54.945000 176.900000 55.475000 183.570000 ;
      RECT 54.945000 186.900000 55.475000 193.570000 ;
      RECT 55.575000 128.730000 56.105000 133.925000 ;
      RECT 55.575000 136.900000 56.105000 143.570000 ;
      RECT 55.575000 146.900000 56.105000 153.570000 ;
      RECT 55.575000 156.900000 56.105000 163.570000 ;
      RECT 55.575000 166.900000 56.105000 173.570000 ;
      RECT 55.585000 136.840000 56.095000 136.900000 ;
      RECT 55.585000 143.570000 56.095000 143.630000 ;
      RECT 55.585000 146.840000 56.095000 146.900000 ;
      RECT 55.585000 153.570000 56.095000 153.630000 ;
      RECT 55.585000 156.840000 56.095000 156.900000 ;
      RECT 55.585000 163.570000 56.095000 163.630000 ;
      RECT 55.585000 166.840000 56.095000 166.900000 ;
      RECT 55.585000 173.570000 56.095000 173.630000 ;
      RECT 56.330000  26.900000 56.860000  33.570000 ;
      RECT 56.330000  36.900000 56.860000  43.570000 ;
      RECT 56.330000  46.900000 56.860000  53.570000 ;
      RECT 56.330000  56.900000 56.860000  63.570000 ;
      RECT 56.330000  66.900000 56.860000  71.725000 ;
      RECT 56.330000 176.900000 56.860000 183.570000 ;
      RECT 56.330000 186.900000 56.860000 193.570000 ;
      RECT 56.340000  26.840000 56.850000  26.900000 ;
      RECT 56.340000  33.570000 56.850000  33.630000 ;
      RECT 56.340000  36.840000 56.850000  36.900000 ;
      RECT 56.340000  43.570000 56.850000  43.630000 ;
      RECT 56.340000  46.840000 56.850000  46.900000 ;
      RECT 56.340000  53.570000 56.850000  53.630000 ;
      RECT 56.340000  56.840000 56.850000  56.900000 ;
      RECT 56.340000  63.570000 56.850000  63.630000 ;
      RECT 56.340000  66.840000 56.850000  66.900000 ;
      RECT 56.340000 176.840000 56.850000 176.900000 ;
      RECT 56.340000 183.570000 56.850000 183.630000 ;
      RECT 56.340000 186.840000 56.850000 186.900000 ;
      RECT 56.340000 193.570000 56.850000 193.630000 ;
      RECT 56.980000  16.365000 57.510000  16.895000 ;
      RECT 57.665000 128.730000 58.195000 133.755000 ;
      RECT 57.665000 136.900000 58.195000 143.570000 ;
      RECT 57.665000 146.900000 58.195000 153.570000 ;
      RECT 57.665000 156.900000 58.195000 163.570000 ;
      RECT 57.665000 166.900000 58.195000 173.570000 ;
      RECT 57.715000  26.900000 58.245000  33.570000 ;
      RECT 57.715000  36.900000 58.245000  43.570000 ;
      RECT 57.715000  46.900000 58.245000  53.570000 ;
      RECT 57.715000  56.900000 58.245000  63.570000 ;
      RECT 57.715000  66.900000 58.245000  71.725000 ;
      RECT 57.715000 176.900000 58.245000 183.570000 ;
      RECT 57.715000 186.900000 58.245000 193.570000 ;
      RECT 58.430000  75.785000 58.600000  80.300000 ;
      RECT 58.430000  82.915000 58.600000  89.020000 ;
      RECT 58.430000  91.930000 58.600000  96.925000 ;
      RECT 58.430000 101.385000 58.600000 106.255000 ;
      RECT 58.430000 110.450000 58.600000 115.270000 ;
      RECT 58.430000 120.080000 58.600000 124.860000 ;
      RECT 59.100000  26.900000 59.630000  33.570000 ;
      RECT 59.100000  36.900000 59.630000  43.570000 ;
      RECT 59.100000  46.900000 59.630000  53.570000 ;
      RECT 59.100000  56.900000 59.630000  63.570000 ;
      RECT 59.100000  66.900000 59.630000  71.725000 ;
      RECT 59.100000 176.900000 59.630000 183.570000 ;
      RECT 59.100000 186.900000 59.630000 193.570000 ;
      RECT 59.110000  26.840000 59.620000  26.900000 ;
      RECT 59.110000  33.570000 59.620000  33.630000 ;
      RECT 59.110000  36.840000 59.620000  36.900000 ;
      RECT 59.110000  43.570000 59.620000  43.630000 ;
      RECT 59.110000  46.840000 59.620000  46.900000 ;
      RECT 59.110000  53.570000 59.620000  53.630000 ;
      RECT 59.110000  56.840000 59.620000  56.900000 ;
      RECT 59.110000  63.570000 59.620000  63.630000 ;
      RECT 59.110000  66.840000 59.620000  66.900000 ;
      RECT 59.110000 176.840000 59.620000 176.900000 ;
      RECT 59.110000 183.570000 59.620000 183.630000 ;
      RECT 59.110000 186.840000 59.620000 186.900000 ;
      RECT 59.110000 193.570000 59.620000 193.630000 ;
      RECT 59.755000 128.730000 60.285000 133.925000 ;
      RECT 59.755000 136.900000 60.285000 143.570000 ;
      RECT 59.755000 146.900000 60.285000 153.570000 ;
      RECT 59.755000 156.900000 60.285000 163.570000 ;
      RECT 59.755000 166.900000 60.285000 173.570000 ;
      RECT 59.765000 136.840000 60.275000 136.900000 ;
      RECT 59.765000 143.570000 60.275000 143.630000 ;
      RECT 59.765000 146.840000 60.275000 146.900000 ;
      RECT 59.765000 153.570000 60.275000 153.630000 ;
      RECT 59.765000 156.840000 60.275000 156.900000 ;
      RECT 59.765000 163.570000 60.275000 163.630000 ;
      RECT 59.765000 166.840000 60.275000 166.900000 ;
      RECT 59.765000 173.570000 60.275000 173.630000 ;
      RECT 60.485000  26.900000 61.015000  33.570000 ;
      RECT 60.485000  36.900000 61.015000  43.570000 ;
      RECT 60.485000  46.900000 61.015000  53.570000 ;
      RECT 60.485000  56.900000 61.015000  63.570000 ;
      RECT 60.485000  66.900000 61.015000  71.725000 ;
      RECT 60.485000 176.900000 61.015000 183.570000 ;
      RECT 60.485000 186.900000 61.015000 193.570000 ;
      RECT 61.845000 128.730000 62.375000 133.755000 ;
      RECT 61.845000 136.900000 62.375000 143.570000 ;
      RECT 61.845000 146.900000 62.375000 153.570000 ;
      RECT 61.845000 156.900000 62.375000 163.570000 ;
      RECT 61.845000 166.900000 62.375000 173.570000 ;
      RECT 61.870000  26.900000 62.400000  33.570000 ;
      RECT 61.870000  36.900000 62.400000  43.570000 ;
      RECT 61.870000  46.900000 62.400000  53.570000 ;
      RECT 61.870000  56.900000 62.400000  63.570000 ;
      RECT 61.870000  66.900000 62.400000  71.725000 ;
      RECT 61.870000 176.900000 62.400000 183.570000 ;
      RECT 61.870000 186.900000 62.400000 193.570000 ;
      RECT 61.880000  26.840000 62.390000  26.900000 ;
      RECT 61.880000  33.570000 62.390000  33.630000 ;
      RECT 61.880000  36.840000 62.390000  36.900000 ;
      RECT 61.880000  43.570000 62.390000  43.630000 ;
      RECT 61.880000  46.840000 62.390000  46.900000 ;
      RECT 61.880000  53.570000 62.390000  53.630000 ;
      RECT 61.880000  56.840000 62.390000  56.900000 ;
      RECT 61.880000  63.570000 62.390000  63.630000 ;
      RECT 61.880000  66.840000 62.390000  66.900000 ;
      RECT 61.880000 176.840000 62.390000 176.900000 ;
      RECT 61.880000 183.570000 62.390000 183.630000 ;
      RECT 61.880000 186.840000 62.390000 186.900000 ;
      RECT 61.880000 193.570000 62.390000 193.630000 ;
      RECT 63.255000  26.900000 63.785000  33.570000 ;
      RECT 63.255000  36.900000 63.785000  43.570000 ;
      RECT 63.255000  46.900000 63.785000  53.570000 ;
      RECT 63.255000  56.900000 63.785000  63.570000 ;
      RECT 63.255000  66.900000 63.785000  71.725000 ;
      RECT 63.255000 176.900000 63.785000 183.570000 ;
      RECT 63.255000 186.900000 63.785000 193.570000 ;
      RECT 63.935000 128.730000 64.465000 133.925000 ;
      RECT 63.935000 136.900000 64.465000 143.570000 ;
      RECT 63.935000 146.900000 64.465000 153.570000 ;
      RECT 63.935000 156.900000 64.465000 163.570000 ;
      RECT 63.935000 166.900000 64.465000 173.570000 ;
      RECT 63.945000 136.840000 64.455000 136.900000 ;
      RECT 63.945000 143.570000 64.455000 143.630000 ;
      RECT 63.945000 146.840000 64.455000 146.900000 ;
      RECT 63.945000 153.570000 64.455000 153.630000 ;
      RECT 63.945000 156.840000 64.455000 156.900000 ;
      RECT 63.945000 163.570000 64.455000 163.630000 ;
      RECT 63.945000 166.840000 64.455000 166.900000 ;
      RECT 63.945000 173.570000 64.455000 173.630000 ;
      RECT 64.640000  26.900000 65.170000  33.570000 ;
      RECT 64.640000  36.900000 65.170000  43.570000 ;
      RECT 64.640000  46.900000 65.170000  53.570000 ;
      RECT 64.640000  56.900000 65.170000  63.570000 ;
      RECT 64.640000  66.900000 65.170000  71.725000 ;
      RECT 64.640000 176.900000 65.170000 183.570000 ;
      RECT 64.640000 186.900000 65.170000 193.570000 ;
      RECT 64.650000  26.840000 65.160000  26.900000 ;
      RECT 64.650000  33.570000 65.160000  33.630000 ;
      RECT 64.650000  36.840000 65.160000  36.900000 ;
      RECT 64.650000  43.570000 65.160000  43.630000 ;
      RECT 64.650000  46.840000 65.160000  46.900000 ;
      RECT 64.650000  53.570000 65.160000  53.630000 ;
      RECT 64.650000  56.840000 65.160000  56.900000 ;
      RECT 64.650000  63.570000 65.160000  63.630000 ;
      RECT 64.650000  66.840000 65.160000  66.900000 ;
      RECT 64.650000 176.840000 65.160000 176.900000 ;
      RECT 64.650000 183.570000 65.160000 183.630000 ;
      RECT 64.650000 186.840000 65.160000 186.900000 ;
      RECT 64.650000 193.570000 65.160000 193.630000 ;
      RECT 66.025000  26.900000 66.555000  33.570000 ;
      RECT 66.025000  36.900000 66.555000  43.570000 ;
      RECT 66.025000  46.900000 66.555000  53.570000 ;
      RECT 66.025000  56.900000 66.555000  63.570000 ;
      RECT 66.025000  66.900000 66.555000  71.725000 ;
      RECT 66.025000 128.730000 66.555000 133.755000 ;
      RECT 66.025000 136.900000 66.555000 143.570000 ;
      RECT 66.025000 146.900000 66.555000 153.570000 ;
      RECT 66.025000 156.900000 66.555000 163.570000 ;
      RECT 66.025000 166.900000 66.555000 173.570000 ;
      RECT 66.025000 176.900000 66.555000 183.570000 ;
      RECT 66.025000 186.900000 66.555000 193.570000 ;
      RECT 66.700000   1.205000 67.230000   1.735000 ;
      RECT 66.710000  75.785000 66.880000  80.535000 ;
      RECT 66.710000  82.785000 66.880000  89.375000 ;
      RECT 66.710000  91.280000 66.880000  97.870000 ;
      RECT 66.710000 101.385000 66.880000 106.255000 ;
      RECT 66.710000 110.450000 66.880000 115.270000 ;
      RECT 66.710000 120.080000 66.880000 124.860000 ;
      RECT 67.290000  26.075000 68.140000  82.180000 ;
      RECT 67.290000  82.350000 68.140000  90.675000 ;
      RECT 67.290000  90.845000 68.140000  98.990000 ;
      RECT 67.575000 101.035000 68.495000 109.275000 ;
      RECT 67.575000 109.445000 68.495000 117.770000 ;
      RECT 67.575000 117.940000 68.495000 194.935000 ;
      RECT 67.605000 100.840000 68.495000 100.865000 ;
      RECT 67.610000   1.080000 73.375000   1.250000 ;
      RECT 67.615000   1.250000 67.785000  17.100000 ;
      RECT 67.615000  17.100000 73.375000  17.270000 ;
      RECT 68.110000   3.280000 68.280000   9.020000 ;
      RECT 68.110000   9.770000 68.280000  16.670000 ;
      RECT 68.335000   1.670000 72.655000   1.840000 ;
      RECT 68.335000   9.320000 72.655000   9.490000 ;
      RECT 68.570000   2.550000 68.740000   9.020000 ;
      RECT 68.570000  10.200000 68.740000  15.660000 ;
      RECT 69.030000   3.280000 69.200000   9.020000 ;
      RECT 69.030000   9.770000 69.200000  16.670000 ;
      RECT 69.190000  24.355000 69.720000  99.925000 ;
      RECT 69.190000 100.095000 69.720000 196.850000 ;
      RECT 69.490000   2.550000 69.660000   9.020000 ;
      RECT 69.490000  10.200000 69.660000  15.660000 ;
      RECT 69.530000  19.010000 70.265000  19.610000 ;
      RECT 69.950000   3.280000 70.120000   9.020000 ;
      RECT 69.950000   9.770000 70.120000  16.670000 ;
      RECT 70.410000   2.550000 70.580000   9.020000 ;
      RECT 70.410000  10.200000 70.580000  15.660000 ;
      RECT 70.495000  17.960000 71.095000  18.695000 ;
      RECT 70.870000   3.280000 71.040000   9.020000 ;
      RECT 70.870000   9.770000 71.040000  16.670000 ;
      RECT 71.330000   2.550000 71.500000   9.020000 ;
      RECT 71.330000  10.200000 71.500000  15.660000 ;
      RECT 71.790000   3.280000 71.960000   9.020000 ;
      RECT 71.790000   9.770000 71.960000  16.670000 ;
      RECT 72.250000   2.550000 72.420000   9.020000 ;
      RECT 72.250000  10.200000 72.420000  15.660000 ;
      RECT 72.710000   2.120000 72.880000   9.020000 ;
      RECT 72.710000   9.770000 72.880000  16.670000 ;
      RECT 73.205000   1.250000 73.375000  17.100000 ;
      RECT 73.875000 196.920000 74.755000 197.780000 ;
    LAYER met1 ;
      RECT  0.000000   0.000000 25.930000   0.295000 ;
      RECT  0.000000   0.000000 26.070000   0.310000 ;
      RECT  0.000000   0.295000 25.930000   0.310000 ;
      RECT  0.000000   0.310000 25.945000   0.325000 ;
      RECT  0.000000   0.310000 75.000000 198.000000 ;
      RECT  0.000000   0.325000 75.000000   3.330000 ;
      RECT  0.000000   3.330000  3.005000 194.995000 ;
      RECT  0.000000 194.995000 75.000000 198.000000 ;
      RECT  3.000000   3.002000 24.390000   3.070000 ;
      RECT  3.000000   3.002000 24.390000   3.070000 ;
      RECT  3.000000   3.070000 24.460000   3.140000 ;
      RECT  3.000000   3.070000 24.460000   3.140000 ;
      RECT  3.000000   3.140000 24.530000   3.210000 ;
      RECT  3.000000   3.140000 24.530000   3.210000 ;
      RECT  3.000000   3.210000 24.600000   3.280000 ;
      RECT  3.000000   3.210000 24.600000   3.280000 ;
      RECT  3.000000   3.280000 24.670000   3.325000 ;
      RECT  3.000000   3.280000 24.670000   3.325000 ;
      RECT  3.000000   3.325000 72.000000 195.000000 ;
      RECT 27.840000   0.000000 75.000000   0.310000 ;
      RECT 27.950000   0.320000 75.000000   0.325000 ;
      RECT 27.965000   0.305000 75.000000   0.320000 ;
      RECT 27.980000   0.000000 75.000000   0.290000 ;
      RECT 27.980000   0.290000 75.000000   0.305000 ;
      RECT 30.950000   3.000000 72.000000   6.330000 ;
      RECT 71.995000   3.330000 75.000000 194.995000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  0.220000 193.910000 ;
      RECT  0.000000   0.000000  0.220000 193.910000 ;
      RECT  0.000000 193.910000 75.000000 198.000000 ;
      RECT  0.000000 193.910000 75.000000 198.000000 ;
      RECT 10.700000   8.165000 11.735000   9.705000 ;
      RECT 10.700000   8.165000 11.735000   9.705000 ;
      RECT 10.700000   9.705000 11.735000   9.715000 ;
      RECT 10.705000   8.160000 11.735000   8.165000 ;
      RECT 10.705000   8.160000 11.735000   8.165000 ;
      RECT 10.705000   9.705000 11.735000   9.710000 ;
      RECT 10.710000   9.710000 11.735000   9.715000 ;
      RECT 10.710000   9.715000 11.515000   9.935000 ;
      RECT 10.720000   8.145000 11.720000   8.160000 ;
      RECT 10.780000   9.715000 11.665000   9.785000 ;
      RECT 10.790000   8.075000 11.650000   8.145000 ;
      RECT 10.850000   9.785000 11.595000   9.855000 ;
      RECT 10.860000   8.005000 11.580000   8.075000 ;
      RECT 10.920000   9.855000 11.525000   9.925000 ;
      RECT 10.930000   7.935000 11.510000   8.005000 ;
      RECT 10.930000   7.935000 11.735000   8.160000 ;
      RECT 10.930000   9.925000 11.515000   9.935000 ;
      RECT 14.030000  25.300000 65.465000  25.370000 ;
      RECT 14.030000  25.300000 65.465000  25.370000 ;
      RECT 14.030000  25.300000 65.860000  25.500000 ;
      RECT 14.030000  25.370000 65.535000  25.440000 ;
      RECT 14.030000  25.370000 65.535000  25.440000 ;
      RECT 14.030000  25.440000 65.605000  25.510000 ;
      RECT 14.030000  25.440000 65.605000  25.510000 ;
      RECT 14.030000  25.500000 65.860000  29.820000 ;
      RECT 14.030000  25.510000 65.675000  25.555000 ;
      RECT 14.030000  25.510000 65.675000  25.555000 ;
      RECT 14.030000  25.555000 65.720000  29.765000 ;
      RECT 14.030000  29.765000 65.650000  29.835000 ;
      RECT 14.030000  29.765000 65.650000  29.835000 ;
      RECT 14.030000  29.820000 64.810000  30.870000 ;
      RECT 14.030000  29.835000 65.580000  29.905000 ;
      RECT 14.030000  29.835000 65.580000  29.905000 ;
      RECT 14.030000  29.905000 65.510000  29.975000 ;
      RECT 14.030000  29.905000 65.510000  29.975000 ;
      RECT 14.030000  29.975000 65.440000  30.045000 ;
      RECT 14.030000  29.975000 65.440000  30.045000 ;
      RECT 14.030000  30.045000 65.370000  30.115000 ;
      RECT 14.030000  30.045000 65.370000  30.115000 ;
      RECT 14.030000  30.115000 65.300000  30.185000 ;
      RECT 14.030000  30.115000 65.300000  30.185000 ;
      RECT 14.030000  30.185000 65.230000  30.255000 ;
      RECT 14.030000  30.185000 65.230000  30.255000 ;
      RECT 14.030000  30.255000 65.160000  30.325000 ;
      RECT 14.030000  30.255000 65.160000  30.325000 ;
      RECT 14.030000  30.325000 65.090000  30.395000 ;
      RECT 14.030000  30.325000 65.090000  30.395000 ;
      RECT 14.030000  30.395000 65.020000  30.465000 ;
      RECT 14.030000  30.395000 65.020000  30.465000 ;
      RECT 14.030000  30.465000 64.950000  30.535000 ;
      RECT 14.030000  30.465000 64.950000  30.535000 ;
      RECT 14.030000  30.535000 64.880000  30.605000 ;
      RECT 14.030000  30.535000 64.880000  30.605000 ;
      RECT 14.030000  30.605000 64.810000  30.675000 ;
      RECT 14.030000  30.605000 64.810000  30.675000 ;
      RECT 14.030000  30.675000 64.755000  30.730000 ;
      RECT 14.030000  30.675000 64.755000  30.730000 ;
      RECT 14.030000  30.730000 15.855000  33.930000 ;
      RECT 14.030000  30.870000 15.995000  33.790000 ;
      RECT 14.030000  33.790000 65.860000  34.750000 ;
      RECT 14.030000  33.930000 64.845000  34.000000 ;
      RECT 14.030000  33.930000 64.845000  34.000000 ;
      RECT 14.030000  34.000000 64.915000  34.070000 ;
      RECT 14.030000  34.000000 64.915000  34.070000 ;
      RECT 14.030000  34.070000 64.985000  34.140000 ;
      RECT 14.030000  34.070000 64.985000  34.140000 ;
      RECT 14.030000  34.140000 65.055000  34.210000 ;
      RECT 14.030000  34.140000 65.055000  34.210000 ;
      RECT 14.030000  34.210000 65.125000  34.280000 ;
      RECT 14.030000  34.210000 65.125000  34.280000 ;
      RECT 14.030000  34.280000 65.195000  34.350000 ;
      RECT 14.030000  34.280000 65.195000  34.350000 ;
      RECT 14.030000  34.350000 65.265000  34.420000 ;
      RECT 14.030000  34.350000 65.265000  34.420000 ;
      RECT 14.030000  34.420000 65.335000  34.490000 ;
      RECT 14.030000  34.420000 65.335000  34.490000 ;
      RECT 14.030000  34.490000 65.405000  34.560000 ;
      RECT 14.030000  34.490000 65.405000  34.560000 ;
      RECT 14.030000  34.560000 65.475000  34.630000 ;
      RECT 14.030000  34.560000 65.475000  34.630000 ;
      RECT 14.030000  34.630000 65.545000  34.700000 ;
      RECT 14.030000  34.630000 65.545000  34.700000 ;
      RECT 14.030000  34.700000 65.615000  34.770000 ;
      RECT 14.030000  34.700000 65.615000  34.770000 ;
      RECT 14.030000  34.750000 65.860000  39.875000 ;
      RECT 14.030000  34.770000 65.685000  34.805000 ;
      RECT 14.030000  34.770000 65.685000  34.805000 ;
      RECT 14.030000  34.805000 65.720000  39.820000 ;
      RECT 14.030000  39.820000 65.650000  39.890000 ;
      RECT 14.030000  39.820000 65.650000  39.890000 ;
      RECT 14.030000  39.875000 64.885000  40.850000 ;
      RECT 14.030000  39.890000 65.580000  39.960000 ;
      RECT 14.030000  39.890000 65.580000  39.960000 ;
      RECT 14.030000  39.960000 65.510000  40.030000 ;
      RECT 14.030000  39.960000 65.510000  40.030000 ;
      RECT 14.030000  40.030000 65.440000  40.100000 ;
      RECT 14.030000  40.030000 65.440000  40.100000 ;
      RECT 14.030000  40.100000 65.370000  40.170000 ;
      RECT 14.030000  40.100000 65.370000  40.170000 ;
      RECT 14.030000  40.170000 65.300000  40.240000 ;
      RECT 14.030000  40.170000 65.300000  40.240000 ;
      RECT 14.030000  40.240000 65.230000  40.310000 ;
      RECT 14.030000  40.240000 65.230000  40.310000 ;
      RECT 14.030000  40.310000 65.160000  40.380000 ;
      RECT 14.030000  40.310000 65.160000  40.380000 ;
      RECT 14.030000  40.380000 65.090000  40.450000 ;
      RECT 14.030000  40.380000 65.090000  40.450000 ;
      RECT 14.030000  40.450000 65.020000  40.520000 ;
      RECT 14.030000  40.450000 65.020000  40.520000 ;
      RECT 14.030000  40.520000 64.950000  40.590000 ;
      RECT 14.030000  40.520000 64.950000  40.590000 ;
      RECT 14.030000  40.590000 64.880000  40.660000 ;
      RECT 14.030000  40.590000 64.880000  40.660000 ;
      RECT 14.030000  40.660000 64.830000  40.710000 ;
      RECT 14.030000  40.660000 64.830000  40.710000 ;
      RECT 14.030000  40.710000 15.855000  43.910000 ;
      RECT 14.030000  40.850000 15.995000  43.770000 ;
      RECT 14.030000  43.770000 65.860000  44.730000 ;
      RECT 14.030000  43.910000 64.845000  43.980000 ;
      RECT 14.030000  43.910000 64.845000  43.980000 ;
      RECT 14.030000  43.980000 64.915000  44.050000 ;
      RECT 14.030000  43.980000 64.915000  44.050000 ;
      RECT 14.030000  44.050000 64.985000  44.120000 ;
      RECT 14.030000  44.050000 64.985000  44.120000 ;
      RECT 14.030000  44.120000 65.055000  44.190000 ;
      RECT 14.030000  44.120000 65.055000  44.190000 ;
      RECT 14.030000  44.190000 65.125000  44.260000 ;
      RECT 14.030000  44.190000 65.125000  44.260000 ;
      RECT 14.030000  44.260000 65.195000  44.330000 ;
      RECT 14.030000  44.260000 65.195000  44.330000 ;
      RECT 14.030000  44.330000 65.265000  44.400000 ;
      RECT 14.030000  44.330000 65.265000  44.400000 ;
      RECT 14.030000  44.400000 65.335000  44.470000 ;
      RECT 14.030000  44.400000 65.335000  44.470000 ;
      RECT 14.030000  44.470000 65.405000  44.540000 ;
      RECT 14.030000  44.470000 65.405000  44.540000 ;
      RECT 14.030000  44.540000 65.475000  44.610000 ;
      RECT 14.030000  44.540000 65.475000  44.610000 ;
      RECT 14.030000  44.610000 65.545000  44.680000 ;
      RECT 14.030000  44.610000 65.545000  44.680000 ;
      RECT 14.030000  44.680000 65.615000  44.750000 ;
      RECT 14.030000  44.680000 65.615000  44.750000 ;
      RECT 14.030000  44.730000 65.860000  49.895000 ;
      RECT 14.030000  44.750000 65.685000  44.785000 ;
      RECT 14.030000  44.750000 65.685000  44.785000 ;
      RECT 14.030000  44.785000 65.720000  49.840000 ;
      RECT 14.030000  49.840000 65.650000  49.910000 ;
      RECT 14.030000  49.840000 65.650000  49.910000 ;
      RECT 14.030000  49.895000 64.885000  50.870000 ;
      RECT 14.030000  49.910000 65.580000  49.980000 ;
      RECT 14.030000  49.910000 65.580000  49.980000 ;
      RECT 14.030000  49.980000 65.510000  50.050000 ;
      RECT 14.030000  49.980000 65.510000  50.050000 ;
      RECT 14.030000  50.050000 65.440000  50.120000 ;
      RECT 14.030000  50.050000 65.440000  50.120000 ;
      RECT 14.030000  50.120000 65.370000  50.190000 ;
      RECT 14.030000  50.120000 65.370000  50.190000 ;
      RECT 14.030000  50.190000 65.300000  50.260000 ;
      RECT 14.030000  50.190000 65.300000  50.260000 ;
      RECT 14.030000  50.260000 65.230000  50.330000 ;
      RECT 14.030000  50.260000 65.230000  50.330000 ;
      RECT 14.030000  50.330000 65.160000  50.400000 ;
      RECT 14.030000  50.330000 65.160000  50.400000 ;
      RECT 14.030000  50.400000 65.090000  50.470000 ;
      RECT 14.030000  50.400000 65.090000  50.470000 ;
      RECT 14.030000  50.470000 65.020000  50.540000 ;
      RECT 14.030000  50.470000 65.020000  50.540000 ;
      RECT 14.030000  50.540000 64.950000  50.610000 ;
      RECT 14.030000  50.540000 64.950000  50.610000 ;
      RECT 14.030000  50.610000 64.880000  50.680000 ;
      RECT 14.030000  50.610000 64.880000  50.680000 ;
      RECT 14.030000  50.680000 64.830000  50.730000 ;
      RECT 14.030000  50.680000 64.830000  50.730000 ;
      RECT 14.030000  50.730000 15.855000  53.930000 ;
      RECT 14.030000  50.870000 15.995000  53.790000 ;
      RECT 14.030000  53.790000 65.855000  54.745000 ;
      RECT 14.030000  53.930000 64.845000  54.000000 ;
      RECT 14.030000  53.930000 64.845000  54.000000 ;
      RECT 14.030000  54.000000 64.915000  54.070000 ;
      RECT 14.030000  54.000000 64.915000  54.070000 ;
      RECT 14.030000  54.070000 64.985000  54.140000 ;
      RECT 14.030000  54.070000 64.985000  54.140000 ;
      RECT 14.030000  54.140000 65.055000  54.210000 ;
      RECT 14.030000  54.140000 65.055000  54.210000 ;
      RECT 14.030000  54.210000 65.125000  54.280000 ;
      RECT 14.030000  54.210000 65.125000  54.280000 ;
      RECT 14.030000  54.280000 65.195000  54.350000 ;
      RECT 14.030000  54.280000 65.195000  54.350000 ;
      RECT 14.030000  54.350000 65.265000  54.420000 ;
      RECT 14.030000  54.350000 65.265000  54.420000 ;
      RECT 14.030000  54.420000 65.335000  54.490000 ;
      RECT 14.030000  54.420000 65.335000  54.490000 ;
      RECT 14.030000  54.490000 65.405000  54.560000 ;
      RECT 14.030000  54.490000 65.405000  54.560000 ;
      RECT 14.030000  54.560000 65.475000  54.630000 ;
      RECT 14.030000  54.560000 65.475000  54.630000 ;
      RECT 14.030000  54.630000 65.545000  54.700000 ;
      RECT 14.030000  54.630000 65.545000  54.700000 ;
      RECT 14.030000  54.700000 65.615000  54.770000 ;
      RECT 14.030000  54.700000 65.615000  54.770000 ;
      RECT 14.030000  54.745000 65.855000  59.880000 ;
      RECT 14.030000  54.770000 65.685000  54.800000 ;
      RECT 14.030000  54.770000 65.685000  54.800000 ;
      RECT 14.030000  54.800000 65.715000  59.825000 ;
      RECT 14.030000  59.825000 65.645000  59.895000 ;
      RECT 14.030000  59.825000 65.645000  59.895000 ;
      RECT 14.030000  59.880000 64.885000  60.850000 ;
      RECT 14.030000  59.895000 65.575000  59.965000 ;
      RECT 14.030000  59.895000 65.575000  59.965000 ;
      RECT 14.030000  59.965000 65.505000  60.035000 ;
      RECT 14.030000  59.965000 65.505000  60.035000 ;
      RECT 14.030000  60.035000 65.435000  60.105000 ;
      RECT 14.030000  60.035000 65.435000  60.105000 ;
      RECT 14.030000  60.105000 65.365000  60.175000 ;
      RECT 14.030000  60.105000 65.365000  60.175000 ;
      RECT 14.030000  60.175000 65.295000  60.245000 ;
      RECT 14.030000  60.175000 65.295000  60.245000 ;
      RECT 14.030000  60.245000 65.225000  60.315000 ;
      RECT 14.030000  60.245000 65.225000  60.315000 ;
      RECT 14.030000  60.315000 65.155000  60.385000 ;
      RECT 14.030000  60.315000 65.155000  60.385000 ;
      RECT 14.030000  60.385000 65.085000  60.455000 ;
      RECT 14.030000  60.385000 65.085000  60.455000 ;
      RECT 14.030000  60.455000 65.015000  60.525000 ;
      RECT 14.030000  60.455000 65.015000  60.525000 ;
      RECT 14.030000  60.525000 64.945000  60.595000 ;
      RECT 14.030000  60.525000 64.945000  60.595000 ;
      RECT 14.030000  60.595000 64.875000  60.665000 ;
      RECT 14.030000  60.595000 64.875000  60.665000 ;
      RECT 14.030000  60.665000 64.830000  60.710000 ;
      RECT 14.030000  60.665000 64.830000  60.710000 ;
      RECT 14.030000  60.710000 15.855000  63.910000 ;
      RECT 14.030000  60.850000 15.995000  63.770000 ;
      RECT 14.030000  63.770000 65.855000  64.735000 ;
      RECT 14.030000  63.910000 64.830000  63.980000 ;
      RECT 14.030000  63.910000 64.830000  63.980000 ;
      RECT 14.030000  63.980000 64.900000  64.050000 ;
      RECT 14.030000  63.980000 64.900000  64.050000 ;
      RECT 14.030000  64.050000 64.970000  64.120000 ;
      RECT 14.030000  64.050000 64.970000  64.120000 ;
      RECT 14.030000  64.120000 65.040000  64.190000 ;
      RECT 14.030000  64.120000 65.040000  64.190000 ;
      RECT 14.030000  64.190000 65.110000  64.260000 ;
      RECT 14.030000  64.190000 65.110000  64.260000 ;
      RECT 14.030000  64.260000 65.180000  64.330000 ;
      RECT 14.030000  64.260000 65.180000  64.330000 ;
      RECT 14.030000  64.330000 65.250000  64.400000 ;
      RECT 14.030000  64.330000 65.250000  64.400000 ;
      RECT 14.030000  64.400000 65.320000  64.470000 ;
      RECT 14.030000  64.400000 65.320000  64.470000 ;
      RECT 14.030000  64.470000 65.390000  64.540000 ;
      RECT 14.030000  64.470000 65.390000  64.540000 ;
      RECT 14.030000  64.540000 65.460000  64.610000 ;
      RECT 14.030000  64.540000 65.460000  64.610000 ;
      RECT 14.030000  64.610000 65.530000  64.680000 ;
      RECT 14.030000  64.610000 65.530000  64.680000 ;
      RECT 14.030000  64.680000 65.600000  64.750000 ;
      RECT 14.030000  64.680000 65.600000  64.750000 ;
      RECT 14.030000  64.735000 65.855000  69.880000 ;
      RECT 14.030000  64.750000 65.670000  64.795000 ;
      RECT 14.030000  64.750000 65.670000  64.795000 ;
      RECT 14.030000  64.795000 65.715000  69.825000 ;
      RECT 14.030000  69.825000 65.645000  69.895000 ;
      RECT 14.030000  69.825000 65.645000  69.895000 ;
      RECT 14.030000  69.880000 64.885000  70.850000 ;
      RECT 14.030000  69.895000 65.575000  69.965000 ;
      RECT 14.030000  69.895000 65.575000  69.965000 ;
      RECT 14.030000  69.965000 65.505000  70.035000 ;
      RECT 14.030000  69.965000 65.505000  70.035000 ;
      RECT 14.030000  70.035000 65.435000  70.105000 ;
      RECT 14.030000  70.035000 65.435000  70.105000 ;
      RECT 14.030000  70.105000 65.365000  70.175000 ;
      RECT 14.030000  70.105000 65.365000  70.175000 ;
      RECT 14.030000  70.175000 65.295000  70.245000 ;
      RECT 14.030000  70.175000 65.295000  70.245000 ;
      RECT 14.030000  70.245000 65.225000  70.315000 ;
      RECT 14.030000  70.245000 65.225000  70.315000 ;
      RECT 14.030000  70.315000 65.155000  70.385000 ;
      RECT 14.030000  70.315000 65.155000  70.385000 ;
      RECT 14.030000  70.385000 65.085000  70.455000 ;
      RECT 14.030000  70.385000 65.085000  70.455000 ;
      RECT 14.030000  70.455000 65.015000  70.525000 ;
      RECT 14.030000  70.455000 65.015000  70.525000 ;
      RECT 14.030000  70.525000 64.945000  70.595000 ;
      RECT 14.030000  70.525000 64.945000  70.595000 ;
      RECT 14.030000  70.595000 64.875000  70.665000 ;
      RECT 14.030000  70.595000 64.875000  70.665000 ;
      RECT 14.030000  70.665000 64.830000  70.710000 ;
      RECT 14.030000  70.665000 64.830000  70.710000 ;
      RECT 14.030000  70.710000 15.855000  73.910000 ;
      RECT 14.030000  70.850000 15.995000  73.770000 ;
      RECT 14.030000  73.770000 65.550000  74.180000 ;
      RECT 14.030000  73.910000 65.085000  73.980000 ;
      RECT 14.030000  73.980000 65.155000  74.050000 ;
      RECT 14.030000  74.050000 65.225000  74.120000 ;
      RECT 14.030000  74.120000 65.295000  74.180000 ;
      RECT 14.030000  74.180000 65.760000  74.390000 ;
      RECT 14.065000  25.265000 65.430000  25.300000 ;
      RECT 14.065000  25.265000 65.430000  25.300000 ;
      RECT 14.100000  74.180000 65.350000  74.250000 ;
      RECT 14.135000  25.195000 65.360000  25.265000 ;
      RECT 14.135000  25.195000 65.360000  25.265000 ;
      RECT 14.170000  74.250000 65.425000  74.320000 ;
      RECT 14.205000  25.125000 65.290000  25.195000 ;
      RECT 14.205000  25.125000 65.290000  25.195000 ;
      RECT 14.240000  73.910000 65.085000  73.980000 ;
      RECT 14.240000  73.910000 65.085000  73.980000 ;
      RECT 14.240000  73.980000 65.155000  74.050000 ;
      RECT 14.240000  73.980000 65.155000  74.050000 ;
      RECT 14.240000  74.050000 65.225000  74.120000 ;
      RECT 14.240000  74.050000 65.225000  74.120000 ;
      RECT 14.240000  74.120000 65.295000  74.180000 ;
      RECT 14.240000  74.120000 65.295000  74.180000 ;
      RECT 14.240000  74.180000 65.350000  74.250000 ;
      RECT 14.240000  74.180000 65.350000  74.250000 ;
      RECT 14.240000  74.250000 65.425000  74.320000 ;
      RECT 14.240000  74.250000 65.425000  74.320000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.390000 65.565000  74.460000 ;
      RECT 14.240000  74.390000 65.565000  74.460000 ;
      RECT 14.240000  74.390000 65.860000  74.490000 ;
      RECT 14.240000  74.460000 65.635000  74.530000 ;
      RECT 14.240000  74.460000 65.635000  74.530000 ;
      RECT 14.240000  74.490000 65.860000  98.700000 ;
      RECT 14.240000  74.530000 65.705000  74.545000 ;
      RECT 14.240000  74.530000 65.705000  74.545000 ;
      RECT 14.240000  74.545000 65.720000  98.840000 ;
      RECT 14.240000  98.700000 75.000000 129.820000 ;
      RECT 14.240000  98.840000 75.000000 129.820000 ;
      RECT 14.240000 129.820000 75.000000 130.705000 ;
      RECT 14.240000 134.795000 75.000000 139.825000 ;
      RECT 14.240000 134.795000 75.000000 139.825000 ;
      RECT 14.240000 139.825000 75.000000 140.710000 ;
      RECT 14.240000 144.795000 75.000000 149.825000 ;
      RECT 14.240000 144.795000 75.000000 149.825000 ;
      RECT 14.240000 149.825000 75.000000 150.710000 ;
      RECT 14.240000 154.795000 75.000000 159.825000 ;
      RECT 14.240000 154.795000 75.000000 159.825000 ;
      RECT 14.240000 159.825000 75.000000 160.710000 ;
      RECT 14.240000 164.795000 75.000000 169.825000 ;
      RECT 14.240000 164.795000 75.000000 169.825000 ;
      RECT 14.240000 169.825000 75.000000 170.710000 ;
      RECT 14.240000 174.795000 75.000000 179.825000 ;
      RECT 14.240000 174.795000 75.000000 179.825000 ;
      RECT 14.240000 179.825000 75.000000 180.710000 ;
      RECT 14.240000 184.795000 75.000000 189.825000 ;
      RECT 14.240000 184.795000 75.000000 189.825000 ;
      RECT 14.240000 189.825000 75.000000 190.710000 ;
      RECT 14.275000  25.055000 65.220000  25.125000 ;
      RECT 14.275000  25.055000 65.220000  25.125000 ;
      RECT 14.285000 134.750000 75.000000 134.795000 ;
      RECT 14.285000 134.750000 75.000000 134.795000 ;
      RECT 14.285000 144.750000 75.000000 144.795000 ;
      RECT 14.285000 144.750000 75.000000 144.795000 ;
      RECT 14.285000 154.750000 75.000000 154.795000 ;
      RECT 14.285000 154.750000 75.000000 154.795000 ;
      RECT 14.285000 164.750000 75.000000 164.795000 ;
      RECT 14.285000 164.750000 75.000000 164.795000 ;
      RECT 14.285000 174.750000 75.000000 174.795000 ;
      RECT 14.285000 174.750000 75.000000 174.795000 ;
      RECT 14.285000 184.750000 75.000000 184.795000 ;
      RECT 14.285000 184.750000 75.000000 184.795000 ;
      RECT 14.310000 129.820000 75.000000 129.890000 ;
      RECT 14.310000 129.820000 75.000000 129.890000 ;
      RECT 14.310000 139.825000 75.000000 139.895000 ;
      RECT 14.310000 139.825000 75.000000 139.895000 ;
      RECT 14.310000 149.825000 75.000000 149.895000 ;
      RECT 14.310000 149.825000 75.000000 149.895000 ;
      RECT 14.310000 159.825000 75.000000 159.895000 ;
      RECT 14.310000 159.825000 75.000000 159.895000 ;
      RECT 14.310000 169.825000 75.000000 169.895000 ;
      RECT 14.310000 169.825000 75.000000 169.895000 ;
      RECT 14.310000 179.825000 75.000000 179.895000 ;
      RECT 14.310000 179.825000 75.000000 179.895000 ;
      RECT 14.310000 189.825000 75.000000 189.895000 ;
      RECT 14.310000 189.825000 75.000000 189.895000 ;
      RECT 14.345000  24.985000 65.150000  25.055000 ;
      RECT 14.345000  24.985000 65.150000  25.055000 ;
      RECT 14.355000 134.680000 75.000000 134.750000 ;
      RECT 14.355000 134.680000 75.000000 134.750000 ;
      RECT 14.355000 144.680000 75.000000 144.750000 ;
      RECT 14.355000 144.680000 75.000000 144.750000 ;
      RECT 14.355000 154.680000 75.000000 154.750000 ;
      RECT 14.355000 154.680000 75.000000 154.750000 ;
      RECT 14.355000 164.680000 75.000000 164.750000 ;
      RECT 14.355000 164.680000 75.000000 164.750000 ;
      RECT 14.355000 174.680000 75.000000 174.750000 ;
      RECT 14.355000 174.680000 75.000000 174.750000 ;
      RECT 14.355000 184.680000 75.000000 184.750000 ;
      RECT 14.355000 184.680000 75.000000 184.750000 ;
      RECT 14.380000 129.890000 75.000000 129.960000 ;
      RECT 14.380000 129.890000 75.000000 129.960000 ;
      RECT 14.380000 139.895000 75.000000 139.965000 ;
      RECT 14.380000 139.895000 75.000000 139.965000 ;
      RECT 14.380000 149.895000 75.000000 149.965000 ;
      RECT 14.380000 149.895000 75.000000 149.965000 ;
      RECT 14.380000 159.895000 75.000000 159.965000 ;
      RECT 14.380000 159.895000 75.000000 159.965000 ;
      RECT 14.380000 169.895000 75.000000 169.965000 ;
      RECT 14.380000 169.895000 75.000000 169.965000 ;
      RECT 14.380000 179.895000 75.000000 179.965000 ;
      RECT 14.380000 179.895000 75.000000 179.965000 ;
      RECT 14.380000 189.895000 75.000000 189.965000 ;
      RECT 14.380000 189.895000 75.000000 189.965000 ;
      RECT 14.415000  24.915000 65.080000  24.985000 ;
      RECT 14.415000  24.915000 65.080000  24.985000 ;
      RECT 14.425000 134.610000 75.000000 134.680000 ;
      RECT 14.425000 134.610000 75.000000 134.680000 ;
      RECT 14.425000 144.610000 75.000000 144.680000 ;
      RECT 14.425000 144.610000 75.000000 144.680000 ;
      RECT 14.425000 154.610000 75.000000 154.680000 ;
      RECT 14.425000 154.610000 75.000000 154.680000 ;
      RECT 14.425000 164.610000 75.000000 164.680000 ;
      RECT 14.425000 164.610000 75.000000 164.680000 ;
      RECT 14.425000 174.610000 75.000000 174.680000 ;
      RECT 14.425000 174.610000 75.000000 174.680000 ;
      RECT 14.425000 184.610000 75.000000 184.680000 ;
      RECT 14.425000 184.610000 75.000000 184.680000 ;
      RECT 14.450000 129.960000 75.000000 130.030000 ;
      RECT 14.450000 129.960000 75.000000 130.030000 ;
      RECT 14.450000 139.965000 75.000000 140.035000 ;
      RECT 14.450000 139.965000 75.000000 140.035000 ;
      RECT 14.450000 149.965000 75.000000 150.035000 ;
      RECT 14.450000 149.965000 75.000000 150.035000 ;
      RECT 14.450000 159.965000 75.000000 160.035000 ;
      RECT 14.450000 159.965000 75.000000 160.035000 ;
      RECT 14.450000 169.965000 75.000000 170.035000 ;
      RECT 14.450000 169.965000 75.000000 170.035000 ;
      RECT 14.450000 179.965000 75.000000 180.035000 ;
      RECT 14.450000 179.965000 75.000000 180.035000 ;
      RECT 14.450000 189.965000 75.000000 190.035000 ;
      RECT 14.450000 189.965000 75.000000 190.035000 ;
      RECT 14.485000  24.845000 65.010000  24.915000 ;
      RECT 14.485000  24.845000 65.010000  24.915000 ;
      RECT 14.495000 134.540000 75.000000 134.610000 ;
      RECT 14.495000 134.540000 75.000000 134.610000 ;
      RECT 14.495000 144.540000 75.000000 144.610000 ;
      RECT 14.495000 144.540000 75.000000 144.610000 ;
      RECT 14.495000 154.540000 75.000000 154.610000 ;
      RECT 14.495000 154.540000 75.000000 154.610000 ;
      RECT 14.495000 164.540000 75.000000 164.610000 ;
      RECT 14.495000 164.540000 75.000000 164.610000 ;
      RECT 14.495000 174.540000 75.000000 174.610000 ;
      RECT 14.495000 174.540000 75.000000 174.610000 ;
      RECT 14.495000 184.540000 75.000000 184.610000 ;
      RECT 14.495000 184.540000 75.000000 184.610000 ;
      RECT 14.520000 130.030000 75.000000 130.100000 ;
      RECT 14.520000 130.030000 75.000000 130.100000 ;
      RECT 14.520000 140.035000 75.000000 140.105000 ;
      RECT 14.520000 140.035000 75.000000 140.105000 ;
      RECT 14.520000 150.035000 75.000000 150.105000 ;
      RECT 14.520000 150.035000 75.000000 150.105000 ;
      RECT 14.520000 160.035000 75.000000 160.105000 ;
      RECT 14.520000 160.035000 75.000000 160.105000 ;
      RECT 14.520000 170.035000 75.000000 170.105000 ;
      RECT 14.520000 170.035000 75.000000 170.105000 ;
      RECT 14.520000 180.035000 75.000000 180.105000 ;
      RECT 14.520000 180.035000 75.000000 180.105000 ;
      RECT 14.520000 190.035000 75.000000 190.105000 ;
      RECT 14.520000 190.035000 75.000000 190.105000 ;
      RECT 14.555000  24.775000 64.940000  24.845000 ;
      RECT 14.555000  24.775000 64.940000  24.845000 ;
      RECT 14.565000 134.470000 75.000000 134.540000 ;
      RECT 14.565000 134.470000 75.000000 134.540000 ;
      RECT 14.565000 144.470000 75.000000 144.540000 ;
      RECT 14.565000 144.470000 75.000000 144.540000 ;
      RECT 14.565000 154.470000 75.000000 154.540000 ;
      RECT 14.565000 154.470000 75.000000 154.540000 ;
      RECT 14.565000 164.470000 75.000000 164.540000 ;
      RECT 14.565000 164.470000 75.000000 164.540000 ;
      RECT 14.565000 174.470000 75.000000 174.540000 ;
      RECT 14.565000 174.470000 75.000000 174.540000 ;
      RECT 14.565000 184.470000 75.000000 184.540000 ;
      RECT 14.565000 184.470000 75.000000 184.540000 ;
      RECT 14.590000 130.100000 75.000000 130.170000 ;
      RECT 14.590000 130.100000 75.000000 130.170000 ;
      RECT 14.590000 140.105000 75.000000 140.175000 ;
      RECT 14.590000 140.105000 75.000000 140.175000 ;
      RECT 14.590000 150.105000 75.000000 150.175000 ;
      RECT 14.590000 150.105000 75.000000 150.175000 ;
      RECT 14.590000 160.105000 75.000000 160.175000 ;
      RECT 14.590000 160.105000 75.000000 160.175000 ;
      RECT 14.590000 170.105000 75.000000 170.175000 ;
      RECT 14.590000 170.105000 75.000000 170.175000 ;
      RECT 14.590000 180.105000 75.000000 180.175000 ;
      RECT 14.590000 180.105000 75.000000 180.175000 ;
      RECT 14.590000 190.105000 75.000000 190.175000 ;
      RECT 14.590000 190.105000 75.000000 190.175000 ;
      RECT 14.625000  24.705000 64.870000  24.775000 ;
      RECT 14.625000  24.705000 64.870000  24.775000 ;
      RECT 14.635000 134.400000 75.000000 134.470000 ;
      RECT 14.635000 134.400000 75.000000 134.470000 ;
      RECT 14.635000 144.400000 75.000000 144.470000 ;
      RECT 14.635000 144.400000 75.000000 144.470000 ;
      RECT 14.635000 154.400000 75.000000 154.470000 ;
      RECT 14.635000 154.400000 75.000000 154.470000 ;
      RECT 14.635000 164.400000 75.000000 164.470000 ;
      RECT 14.635000 164.400000 75.000000 164.470000 ;
      RECT 14.635000 174.400000 75.000000 174.470000 ;
      RECT 14.635000 174.400000 75.000000 174.470000 ;
      RECT 14.635000 184.400000 75.000000 184.470000 ;
      RECT 14.635000 184.400000 75.000000 184.470000 ;
      RECT 14.660000 130.170000 75.000000 130.240000 ;
      RECT 14.660000 130.170000 75.000000 130.240000 ;
      RECT 14.660000 140.175000 75.000000 140.245000 ;
      RECT 14.660000 140.175000 75.000000 140.245000 ;
      RECT 14.660000 150.175000 75.000000 150.245000 ;
      RECT 14.660000 150.175000 75.000000 150.245000 ;
      RECT 14.660000 160.175000 75.000000 160.245000 ;
      RECT 14.660000 160.175000 75.000000 160.245000 ;
      RECT 14.660000 170.175000 75.000000 170.245000 ;
      RECT 14.660000 170.175000 75.000000 170.245000 ;
      RECT 14.660000 180.175000 75.000000 180.245000 ;
      RECT 14.660000 180.175000 75.000000 180.245000 ;
      RECT 14.660000 190.175000 75.000000 190.245000 ;
      RECT 14.660000 190.175000 75.000000 190.245000 ;
      RECT 14.695000  24.635000 64.800000  24.705000 ;
      RECT 14.695000  24.635000 64.800000  24.705000 ;
      RECT 14.705000 134.330000 75.000000 134.400000 ;
      RECT 14.705000 134.330000 75.000000 134.400000 ;
      RECT 14.705000 144.330000 75.000000 144.400000 ;
      RECT 14.705000 144.330000 75.000000 144.400000 ;
      RECT 14.705000 154.330000 75.000000 154.400000 ;
      RECT 14.705000 154.330000 75.000000 154.400000 ;
      RECT 14.705000 164.330000 75.000000 164.400000 ;
      RECT 14.705000 164.330000 75.000000 164.400000 ;
      RECT 14.705000 174.330000 75.000000 174.400000 ;
      RECT 14.705000 174.330000 75.000000 174.400000 ;
      RECT 14.705000 184.330000 75.000000 184.400000 ;
      RECT 14.705000 184.330000 75.000000 184.400000 ;
      RECT 14.730000 130.240000 75.000000 130.310000 ;
      RECT 14.730000 130.240000 75.000000 130.310000 ;
      RECT 14.730000 140.245000 75.000000 140.315000 ;
      RECT 14.730000 140.245000 75.000000 140.315000 ;
      RECT 14.730000 150.245000 75.000000 150.315000 ;
      RECT 14.730000 150.245000 75.000000 150.315000 ;
      RECT 14.730000 160.245000 75.000000 160.315000 ;
      RECT 14.730000 160.245000 75.000000 160.315000 ;
      RECT 14.730000 170.245000 75.000000 170.315000 ;
      RECT 14.730000 170.245000 75.000000 170.315000 ;
      RECT 14.730000 180.245000 75.000000 180.315000 ;
      RECT 14.730000 180.245000 75.000000 180.315000 ;
      RECT 14.730000 190.245000 75.000000 190.315000 ;
      RECT 14.730000 190.245000 75.000000 190.315000 ;
      RECT 14.765000  24.565000 64.730000  24.635000 ;
      RECT 14.765000  24.565000 64.730000  24.635000 ;
      RECT 14.775000 134.260000 75.000000 134.330000 ;
      RECT 14.775000 134.260000 75.000000 134.330000 ;
      RECT 14.775000 144.260000 75.000000 144.330000 ;
      RECT 14.775000 144.260000 75.000000 144.330000 ;
      RECT 14.775000 154.260000 75.000000 154.330000 ;
      RECT 14.775000 154.260000 75.000000 154.330000 ;
      RECT 14.775000 164.260000 75.000000 164.330000 ;
      RECT 14.775000 164.260000 75.000000 164.330000 ;
      RECT 14.775000 174.260000 75.000000 174.330000 ;
      RECT 14.775000 174.260000 75.000000 174.330000 ;
      RECT 14.775000 184.260000 75.000000 184.330000 ;
      RECT 14.775000 184.260000 75.000000 184.330000 ;
      RECT 14.800000 130.310000 75.000000 130.380000 ;
      RECT 14.800000 130.310000 75.000000 130.380000 ;
      RECT 14.800000 140.315000 75.000000 140.385000 ;
      RECT 14.800000 140.315000 75.000000 140.385000 ;
      RECT 14.800000 150.315000 75.000000 150.385000 ;
      RECT 14.800000 150.315000 75.000000 150.385000 ;
      RECT 14.800000 160.315000 75.000000 160.385000 ;
      RECT 14.800000 160.315000 75.000000 160.385000 ;
      RECT 14.800000 170.315000 75.000000 170.385000 ;
      RECT 14.800000 170.315000 75.000000 170.385000 ;
      RECT 14.800000 180.315000 75.000000 180.385000 ;
      RECT 14.800000 180.315000 75.000000 180.385000 ;
      RECT 14.800000 190.315000 75.000000 190.385000 ;
      RECT 14.800000 190.315000 75.000000 190.385000 ;
      RECT 14.835000  24.495000 64.660000  24.565000 ;
      RECT 14.835000  24.495000 64.660000  24.565000 ;
      RECT 14.845000 134.190000 75.000000 134.260000 ;
      RECT 14.845000 134.190000 75.000000 134.260000 ;
      RECT 14.845000 144.190000 75.000000 144.260000 ;
      RECT 14.845000 144.190000 75.000000 144.260000 ;
      RECT 14.845000 154.190000 75.000000 154.260000 ;
      RECT 14.845000 154.190000 75.000000 154.260000 ;
      RECT 14.845000 164.190000 75.000000 164.260000 ;
      RECT 14.845000 164.190000 75.000000 164.260000 ;
      RECT 14.845000 174.190000 75.000000 174.260000 ;
      RECT 14.845000 174.190000 75.000000 174.260000 ;
      RECT 14.845000 184.190000 75.000000 184.260000 ;
      RECT 14.845000 184.190000 75.000000 184.260000 ;
      RECT 14.870000 130.380000 75.000000 130.450000 ;
      RECT 14.870000 130.380000 75.000000 130.450000 ;
      RECT 14.870000 140.385000 75.000000 140.455000 ;
      RECT 14.870000 140.385000 75.000000 140.455000 ;
      RECT 14.870000 150.385000 75.000000 150.455000 ;
      RECT 14.870000 150.385000 75.000000 150.455000 ;
      RECT 14.870000 160.385000 75.000000 160.455000 ;
      RECT 14.870000 160.385000 75.000000 160.455000 ;
      RECT 14.870000 170.385000 75.000000 170.455000 ;
      RECT 14.870000 170.385000 75.000000 170.455000 ;
      RECT 14.870000 180.385000 75.000000 180.455000 ;
      RECT 14.870000 180.385000 75.000000 180.455000 ;
      RECT 14.870000 190.385000 75.000000 190.455000 ;
      RECT 14.870000 190.385000 75.000000 190.455000 ;
      RECT 14.905000  24.425000 64.590000  24.495000 ;
      RECT 14.905000  24.425000 64.590000  24.495000 ;
      RECT 14.915000 134.120000 75.000000 134.190000 ;
      RECT 14.915000 134.120000 75.000000 134.190000 ;
      RECT 14.915000 144.120000 75.000000 144.190000 ;
      RECT 14.915000 144.120000 75.000000 144.190000 ;
      RECT 14.915000 154.120000 75.000000 154.190000 ;
      RECT 14.915000 154.120000 75.000000 154.190000 ;
      RECT 14.915000 164.120000 75.000000 164.190000 ;
      RECT 14.915000 164.120000 75.000000 164.190000 ;
      RECT 14.915000 174.120000 75.000000 174.190000 ;
      RECT 14.915000 174.120000 75.000000 174.190000 ;
      RECT 14.915000 184.120000 75.000000 184.190000 ;
      RECT 14.915000 184.120000 75.000000 184.190000 ;
      RECT 14.940000 130.450000 75.000000 130.520000 ;
      RECT 14.940000 130.450000 75.000000 130.520000 ;
      RECT 14.940000 140.455000 75.000000 140.525000 ;
      RECT 14.940000 140.455000 75.000000 140.525000 ;
      RECT 14.940000 150.455000 75.000000 150.525000 ;
      RECT 14.940000 150.455000 75.000000 150.525000 ;
      RECT 14.940000 160.455000 75.000000 160.525000 ;
      RECT 14.940000 160.455000 75.000000 160.525000 ;
      RECT 14.940000 170.455000 75.000000 170.525000 ;
      RECT 14.940000 170.455000 75.000000 170.525000 ;
      RECT 14.940000 180.455000 75.000000 180.525000 ;
      RECT 14.940000 180.455000 75.000000 180.525000 ;
      RECT 14.940000 190.455000 75.000000 190.525000 ;
      RECT 14.940000 190.455000 75.000000 190.525000 ;
      RECT 14.975000  24.355000 64.520000  24.425000 ;
      RECT 14.975000  24.355000 64.520000  24.425000 ;
      RECT 14.985000 134.050000 75.000000 134.120000 ;
      RECT 14.985000 134.050000 75.000000 134.120000 ;
      RECT 14.985000 144.050000 75.000000 144.120000 ;
      RECT 14.985000 144.050000 75.000000 144.120000 ;
      RECT 14.985000 154.050000 75.000000 154.120000 ;
      RECT 14.985000 154.050000 75.000000 154.120000 ;
      RECT 14.985000 164.050000 75.000000 164.120000 ;
      RECT 14.985000 164.050000 75.000000 164.120000 ;
      RECT 14.985000 174.050000 75.000000 174.120000 ;
      RECT 14.985000 174.050000 75.000000 174.120000 ;
      RECT 14.985000 184.050000 75.000000 184.120000 ;
      RECT 14.985000 184.050000 75.000000 184.120000 ;
      RECT 15.010000 130.520000 75.000000 130.590000 ;
      RECT 15.010000 130.520000 75.000000 130.590000 ;
      RECT 15.010000 140.525000 75.000000 140.595000 ;
      RECT 15.010000 140.525000 75.000000 140.595000 ;
      RECT 15.010000 150.525000 75.000000 150.595000 ;
      RECT 15.010000 150.525000 75.000000 150.595000 ;
      RECT 15.010000 160.525000 75.000000 160.595000 ;
      RECT 15.010000 160.525000 75.000000 160.595000 ;
      RECT 15.010000 170.525000 75.000000 170.595000 ;
      RECT 15.010000 170.525000 75.000000 170.595000 ;
      RECT 15.010000 180.525000 75.000000 180.595000 ;
      RECT 15.010000 180.525000 75.000000 180.595000 ;
      RECT 15.010000 190.525000 75.000000 190.595000 ;
      RECT 15.010000 190.525000 75.000000 190.595000 ;
      RECT 15.045000  24.285000 64.450000  24.355000 ;
      RECT 15.045000  24.285000 64.450000  24.355000 ;
      RECT 15.055000 133.980000 75.000000 134.050000 ;
      RECT 15.055000 133.980000 75.000000 134.050000 ;
      RECT 15.055000 143.980000 75.000000 144.050000 ;
      RECT 15.055000 143.980000 75.000000 144.050000 ;
      RECT 15.055000 153.980000 75.000000 154.050000 ;
      RECT 15.055000 153.980000 75.000000 154.050000 ;
      RECT 15.055000 163.980000 75.000000 164.050000 ;
      RECT 15.055000 163.980000 75.000000 164.050000 ;
      RECT 15.055000 173.980000 75.000000 174.050000 ;
      RECT 15.055000 173.980000 75.000000 174.050000 ;
      RECT 15.055000 183.980000 75.000000 184.050000 ;
      RECT 15.055000 183.980000 75.000000 184.050000 ;
      RECT 15.080000 130.590000 75.000000 130.660000 ;
      RECT 15.080000 130.590000 75.000000 130.660000 ;
      RECT 15.080000 140.595000 75.000000 140.665000 ;
      RECT 15.080000 140.595000 75.000000 140.665000 ;
      RECT 15.080000 150.595000 75.000000 150.665000 ;
      RECT 15.080000 150.595000 75.000000 150.665000 ;
      RECT 15.080000 160.595000 75.000000 160.665000 ;
      RECT 15.080000 160.595000 75.000000 160.665000 ;
      RECT 15.080000 170.595000 75.000000 170.665000 ;
      RECT 15.080000 170.595000 75.000000 170.665000 ;
      RECT 15.080000 180.595000 75.000000 180.665000 ;
      RECT 15.080000 180.595000 75.000000 180.665000 ;
      RECT 15.080000 190.595000 75.000000 190.665000 ;
      RECT 15.080000 190.595000 75.000000 190.665000 ;
      RECT 15.115000  24.215000 64.380000  24.285000 ;
      RECT 15.115000  24.215000 64.380000  24.285000 ;
      RECT 15.125000 130.660000 75.000000 130.705000 ;
      RECT 15.125000 130.660000 75.000000 130.705000 ;
      RECT 15.125000 133.910000 75.000000 133.980000 ;
      RECT 15.125000 133.910000 75.000000 133.980000 ;
      RECT 15.125000 133.910000 75.000000 134.795000 ;
      RECT 15.125000 140.665000 75.000000 140.710000 ;
      RECT 15.125000 140.665000 75.000000 140.710000 ;
      RECT 15.125000 143.910000 75.000000 143.980000 ;
      RECT 15.125000 143.910000 75.000000 143.980000 ;
      RECT 15.125000 143.910000 75.000000 144.795000 ;
      RECT 15.125000 150.665000 75.000000 150.710000 ;
      RECT 15.125000 150.665000 75.000000 150.710000 ;
      RECT 15.125000 153.910000 75.000000 153.980000 ;
      RECT 15.125000 153.910000 75.000000 153.980000 ;
      RECT 15.125000 153.910000 75.000000 154.795000 ;
      RECT 15.125000 160.665000 75.000000 160.710000 ;
      RECT 15.125000 160.665000 75.000000 160.710000 ;
      RECT 15.125000 163.910000 75.000000 163.980000 ;
      RECT 15.125000 163.910000 75.000000 163.980000 ;
      RECT 15.125000 163.910000 75.000000 164.795000 ;
      RECT 15.125000 170.665000 75.000000 170.710000 ;
      RECT 15.125000 170.665000 75.000000 170.710000 ;
      RECT 15.125000 173.910000 75.000000 173.980000 ;
      RECT 15.125000 173.910000 75.000000 173.980000 ;
      RECT 15.125000 173.910000 75.000000 174.795000 ;
      RECT 15.125000 180.665000 75.000000 180.710000 ;
      RECT 15.125000 180.665000 75.000000 180.710000 ;
      RECT 15.125000 183.910000 75.000000 183.980000 ;
      RECT 15.125000 183.910000 75.000000 183.980000 ;
      RECT 15.125000 183.910000 75.000000 184.795000 ;
      RECT 15.125000 190.665000 75.000000 190.710000 ;
      RECT 15.125000 190.665000 75.000000 190.710000 ;
      RECT 15.185000  24.145000 64.310000  24.215000 ;
      RECT 15.185000  24.145000 64.310000  24.215000 ;
      RECT 15.255000  24.075000 64.240000  24.145000 ;
      RECT 15.255000  24.075000 64.240000  24.145000 ;
      RECT 15.325000  24.005000 64.170000  24.075000 ;
      RECT 15.325000  24.005000 64.170000  24.075000 ;
      RECT 15.395000  23.935000 64.100000  24.005000 ;
      RECT 15.395000  23.935000 64.100000  24.005000 ;
      RECT 15.465000  23.865000 64.030000  23.935000 ;
      RECT 15.465000  23.865000 64.030000  23.935000 ;
      RECT 15.520000 130.705000 75.000000 130.845000 ;
      RECT 15.520000 140.710000 75.000000 140.850000 ;
      RECT 15.520000 150.710000 75.000000 150.850000 ;
      RECT 15.520000 160.710000 75.000000 160.850000 ;
      RECT 15.520000 170.710000 75.000000 170.850000 ;
      RECT 15.520000 180.710000 75.000000 180.850000 ;
      RECT 15.520000 190.710000 75.000000 190.850000 ;
      RECT 15.535000  23.795000 63.960000  23.865000 ;
      RECT 15.535000  23.795000 63.960000  23.865000 ;
      RECT 15.605000  23.725000 63.890000  23.795000 ;
      RECT 15.605000  23.725000 63.890000  23.795000 ;
      RECT 15.660000 133.770000 75.000000 133.910000 ;
      RECT 15.660000 143.770000 75.000000 143.910000 ;
      RECT 15.660000 153.770000 75.000000 153.910000 ;
      RECT 15.660000 163.770000 75.000000 163.910000 ;
      RECT 15.660000 173.770000 75.000000 173.910000 ;
      RECT 15.660000 183.770000 75.000000 183.910000 ;
      RECT 15.675000  23.655000 63.820000  23.725000 ;
      RECT 15.675000  23.655000 63.820000  23.725000 ;
      RECT 15.745000  23.585000 63.750000  23.655000 ;
      RECT 15.745000  23.585000 63.750000  23.655000 ;
      RECT 15.815000  23.515000 63.680000  23.585000 ;
      RECT 15.815000  23.515000 63.680000  23.585000 ;
      RECT 15.885000  23.445000 63.610000  23.515000 ;
      RECT 15.885000  23.445000 63.610000  23.515000 ;
      RECT 15.955000  23.375000 63.540000  23.445000 ;
      RECT 15.955000  23.375000 63.540000  23.445000 ;
      RECT 16.025000  23.305000 63.470000  23.375000 ;
      RECT 16.025000  23.305000 63.470000  23.375000 ;
      RECT 16.095000  23.235000 63.400000  23.305000 ;
      RECT 16.095000  23.235000 63.400000  23.305000 ;
      RECT 16.165000  23.165000 63.330000  23.235000 ;
      RECT 16.165000  23.165000 63.330000  23.235000 ;
      RECT 16.235000  23.095000 63.260000  23.165000 ;
      RECT 16.235000  23.095000 63.260000  23.165000 ;
      RECT 16.305000  23.025000 63.190000  23.095000 ;
      RECT 16.305000  23.025000 63.190000  23.095000 ;
      RECT 16.375000  22.955000 63.120000  23.025000 ;
      RECT 16.375000  22.955000 63.120000  23.025000 ;
      RECT 16.445000  22.885000 63.050000  22.955000 ;
      RECT 16.445000  22.885000 63.050000  22.955000 ;
      RECT 16.515000  22.815000 62.980000  22.885000 ;
      RECT 16.515000  22.815000 62.980000  22.885000 ;
      RECT 16.585000  22.745000 62.910000  22.815000 ;
      RECT 16.585000  22.745000 62.910000  22.815000 ;
      RECT 16.655000  22.675000 62.840000  22.745000 ;
      RECT 16.655000  22.675000 62.840000  22.745000 ;
      RECT 16.725000  22.605000 62.770000  22.675000 ;
      RECT 16.725000  22.605000 62.770000  22.675000 ;
      RECT 16.795000  22.535000 62.700000  22.605000 ;
      RECT 16.795000  22.535000 62.700000  22.605000 ;
      RECT 16.865000  22.465000 62.630000  22.535000 ;
      RECT 16.865000  22.465000 62.630000  22.535000 ;
      RECT 16.935000  22.395000 62.560000  22.465000 ;
      RECT 16.935000  22.395000 62.560000  22.465000 ;
      RECT 17.005000  22.325000 62.490000  22.395000 ;
      RECT 17.005000  22.325000 62.490000  22.395000 ;
      RECT 17.075000  22.255000 62.420000  22.325000 ;
      RECT 17.075000  22.255000 62.420000  22.325000 ;
      RECT 17.140000   5.235000 17.350000   9.250000 ;
      RECT 17.140000   5.235000 17.490000   9.250000 ;
      RECT 17.140000   9.250000 17.490000   9.600000 ;
      RECT 17.145000  22.185000 62.350000  22.255000 ;
      RECT 17.145000  22.185000 62.350000  22.255000 ;
      RECT 17.210000   5.165000 17.350000   5.235000 ;
      RECT 17.210000   9.250000 17.350000   9.320000 ;
      RECT 17.215000  22.115000 62.280000  22.185000 ;
      RECT 17.215000  22.115000 62.280000  22.185000 ;
      RECT 17.280000   5.095000 17.350000   5.165000 ;
      RECT 17.280000   9.320000 17.350000   9.390000 ;
      RECT 17.285000  22.045000 62.210000  22.115000 ;
      RECT 17.285000  22.045000 62.210000  22.115000 ;
      RECT 17.320000   5.055000 17.490000   5.235000 ;
      RECT 17.355000  21.975000 62.140000  22.045000 ;
      RECT 17.355000  21.975000 62.140000  22.045000 ;
      RECT 17.425000  21.905000 53.815000  21.975000 ;
      RECT 17.425000  21.905000 53.815000  21.975000 ;
      RECT 17.495000  21.835000 53.815000  21.905000 ;
      RECT 17.495000  21.835000 53.815000  21.905000 ;
      RECT 17.495000  21.835000 65.660000  25.300000 ;
      RECT 17.565000  21.765000 53.815000  21.835000 ;
      RECT 17.565000  21.765000 53.815000  21.835000 ;
      RECT 17.570000   9.680000 55.880000   9.800000 ;
      RECT 17.635000  21.695000 53.815000  21.765000 ;
      RECT 17.635000  21.695000 53.815000  21.765000 ;
      RECT 17.705000  21.625000 53.815000  21.695000 ;
      RECT 17.705000  21.625000 53.815000  21.695000 ;
      RECT 17.775000  21.555000 53.815000  21.625000 ;
      RECT 17.775000  21.555000 53.815000  21.625000 ;
      RECT 17.845000  21.485000 53.815000  21.555000 ;
      RECT 17.845000  21.485000 53.815000  21.555000 ;
      RECT 17.915000  21.415000 53.815000  21.485000 ;
      RECT 17.915000  21.415000 53.815000  21.485000 ;
      RECT 17.985000  21.345000 53.815000  21.415000 ;
      RECT 17.985000  21.345000 53.815000  21.415000 ;
      RECT 18.055000  21.275000 53.815000  21.345000 ;
      RECT 18.055000  21.275000 53.815000  21.345000 ;
      RECT 18.125000  21.205000 53.815000  21.275000 ;
      RECT 18.125000  21.205000 53.815000  21.275000 ;
      RECT 18.195000  21.135000 53.815000  21.205000 ;
      RECT 18.195000  21.135000 53.815000  21.205000 ;
      RECT 18.265000  21.065000 53.815000  21.135000 ;
      RECT 18.265000  21.065000 53.815000  21.135000 ;
      RECT 18.335000  20.995000 53.815000  21.065000 ;
      RECT 18.335000  20.995000 53.815000  21.065000 ;
      RECT 18.405000  20.925000 53.815000  20.995000 ;
      RECT 18.405000  20.925000 53.815000  20.995000 ;
      RECT 18.475000  20.855000 53.815000  20.925000 ;
      RECT 18.475000  20.855000 53.815000  20.925000 ;
      RECT 18.545000  20.785000 53.815000  20.855000 ;
      RECT 18.545000  20.785000 53.815000  20.855000 ;
      RECT 18.580000 193.770000 75.000000 193.910000 ;
      RECT 18.615000  20.715000 53.815000  20.785000 ;
      RECT 18.615000  20.715000 53.815000  20.785000 ;
      RECT 18.685000  20.645000 53.815000  20.715000 ;
      RECT 18.685000  20.645000 53.815000  20.715000 ;
      RECT 18.755000  20.575000 53.815000  20.645000 ;
      RECT 18.755000  20.575000 53.815000  20.645000 ;
      RECT 18.825000  20.505000 53.815000  20.575000 ;
      RECT 18.825000  20.505000 53.815000  20.575000 ;
      RECT 18.895000  20.435000 53.815000  20.505000 ;
      RECT 18.895000  20.435000 53.815000  20.505000 ;
      RECT 18.965000  20.365000 53.815000  20.435000 ;
      RECT 18.965000  20.365000 53.815000  20.435000 ;
      RECT 19.035000  20.295000 53.815000  20.365000 ;
      RECT 19.035000  20.295000 53.815000  20.365000 ;
      RECT 19.105000  20.225000 53.815000  20.295000 ;
      RECT 19.105000  20.225000 53.815000  20.295000 ;
      RECT 19.175000  20.155000 53.815000  20.225000 ;
      RECT 19.175000  20.155000 53.815000  20.225000 ;
      RECT 19.245000  20.085000 53.815000  20.155000 ;
      RECT 19.245000  20.085000 53.815000  20.155000 ;
      RECT 19.315000  20.015000 53.815000  20.085000 ;
      RECT 19.315000  20.015000 53.815000  20.085000 ;
      RECT 19.385000  19.945000 53.815000  20.015000 ;
      RECT 19.385000  19.945000 53.815000  20.015000 ;
      RECT 19.400000  19.930000 53.955000  21.835000 ;
      RECT 19.455000  19.875000 53.815000  19.945000 ;
      RECT 19.455000  19.875000 53.815000  19.945000 ;
      RECT 19.510000  19.820000 53.815000  19.875000 ;
      RECT 19.510000  19.820000 53.815000  19.875000 ;
      RECT 19.580000  19.750000 53.870000  19.820000 ;
      RECT 19.580000  19.750000 53.870000  19.820000 ;
      RECT 19.650000  19.680000 53.940000  19.750000 ;
      RECT 19.650000  19.680000 53.940000  19.750000 ;
      RECT 19.720000  19.610000 54.010000  19.680000 ;
      RECT 19.720000  19.610000 54.010000  19.680000 ;
      RECT 19.790000  19.540000 54.080000  19.610000 ;
      RECT 19.790000  19.540000 54.080000  19.610000 ;
      RECT 19.860000  19.470000 54.150000  19.540000 ;
      RECT 19.860000  19.470000 54.150000  19.540000 ;
      RECT 19.930000  19.400000 54.220000  19.470000 ;
      RECT 19.930000  19.400000 54.220000  19.470000 ;
      RECT 20.000000  19.330000 54.290000  19.400000 ;
      RECT 20.000000  19.330000 54.290000  19.400000 ;
      RECT 20.070000  19.260000 54.360000  19.330000 ;
      RECT 20.070000  19.260000 54.360000  19.330000 ;
      RECT 20.140000  19.190000 54.430000  19.260000 ;
      RECT 20.140000  19.190000 54.430000  19.260000 ;
      RECT 20.210000  19.120000 54.500000  19.190000 ;
      RECT 20.210000  19.120000 54.500000  19.190000 ;
      RECT 20.280000  19.050000 54.570000  19.120000 ;
      RECT 20.280000  19.050000 54.570000  19.120000 ;
      RECT 20.350000  18.980000 54.640000  19.050000 ;
      RECT 20.350000  18.980000 54.640000  19.050000 ;
      RECT 20.420000  18.910000 54.710000  18.980000 ;
      RECT 20.420000  18.910000 54.710000  18.980000 ;
      RECT 20.490000  18.840000 54.780000  18.910000 ;
      RECT 20.490000  18.840000 54.780000  18.910000 ;
      RECT 20.560000  18.770000 54.850000  18.840000 ;
      RECT 20.560000  18.770000 54.850000  18.840000 ;
      RECT 20.630000  18.700000 54.920000  18.770000 ;
      RECT 20.630000  18.700000 54.920000  18.770000 ;
      RECT 20.700000  18.630000 54.990000  18.700000 ;
      RECT 20.700000  18.630000 54.990000  18.700000 ;
      RECT 20.770000  18.560000 55.060000  18.630000 ;
      RECT 20.770000  18.560000 55.060000  18.630000 ;
      RECT 20.775000   0.000000 20.785000   1.600000 ;
      RECT 20.775000   1.600000 20.785000   1.760000 ;
      RECT 20.840000  18.490000 55.130000  18.560000 ;
      RECT 20.840000  18.490000 55.130000  18.560000 ;
      RECT 20.910000  18.420000 55.200000  18.490000 ;
      RECT 20.910000  18.420000 55.200000  18.490000 ;
      RECT 20.980000  18.350000 55.270000  18.420000 ;
      RECT 20.980000  18.350000 55.270000  18.420000 ;
      RECT 21.050000  18.280000 55.340000  18.350000 ;
      RECT 21.050000  18.280000 55.340000  18.350000 ;
      RECT 21.120000  18.210000 55.410000  18.280000 ;
      RECT 21.120000  18.210000 55.410000  18.280000 ;
      RECT 21.190000  18.140000 55.480000  18.210000 ;
      RECT 21.190000  18.140000 55.480000  18.210000 ;
      RECT 21.260000  18.070000 55.550000  18.140000 ;
      RECT 21.260000  18.070000 55.550000  18.140000 ;
      RECT 21.330000  18.000000 55.620000  18.070000 ;
      RECT 21.330000  18.000000 55.620000  18.070000 ;
      RECT 21.400000  17.930000 55.690000  18.000000 ;
      RECT 21.400000  17.930000 55.690000  18.000000 ;
      RECT 21.470000  17.860000 55.760000  17.930000 ;
      RECT 21.470000  17.860000 55.760000  17.930000 ;
      RECT 21.540000  17.790000 55.830000  17.860000 ;
      RECT 21.540000  17.790000 55.830000  17.860000 ;
      RECT 21.555000  17.775000 53.955000  19.930000 ;
      RECT 21.610000  17.720000 55.900000  17.790000 ;
      RECT 21.610000  17.720000 55.900000  17.790000 ;
      RECT 21.620000  17.710000 55.970000  17.720000 ;
      RECT 21.620000  17.710000 55.970000  17.720000 ;
      RECT 21.690000  17.640000 55.970000  17.710000 ;
      RECT 21.690000  17.640000 55.970000  17.710000 ;
      RECT 21.760000  17.570000 55.970000  17.640000 ;
      RECT 21.760000  17.570000 55.970000  17.640000 ;
      RECT 21.830000  17.500000 55.970000  17.570000 ;
      RECT 21.830000  17.500000 55.970000  17.570000 ;
      RECT 21.900000  17.430000 55.970000  17.500000 ;
      RECT 21.900000  17.430000 55.970000  17.500000 ;
      RECT 21.970000  17.360000 55.970000  17.430000 ;
      RECT 21.970000  17.360000 55.970000  17.430000 ;
      RECT 21.970000  17.360000 56.110000  17.775000 ;
      RECT 53.675000   0.000000 53.955000   7.875000 ;
      RECT 53.675000   7.875000 55.760000   9.680000 ;
      RECT 53.815000   8.000000 53.885000   8.070000 ;
      RECT 53.815000   8.070000 53.955000   8.140000 ;
      RECT 53.815000   8.140000 54.025000   8.210000 ;
      RECT 53.815000   8.210000 54.095000   8.280000 ;
      RECT 53.815000   8.280000 54.165000   8.350000 ;
      RECT 53.815000   8.350000 54.235000   8.420000 ;
      RECT 53.815000   8.420000 54.305000   8.490000 ;
      RECT 53.815000   8.490000 54.375000   8.560000 ;
      RECT 53.815000   8.560000 54.445000   8.630000 ;
      RECT 53.815000   8.630000 54.515000   8.700000 ;
      RECT 53.815000   8.700000 54.585000   8.770000 ;
      RECT 53.815000   8.770000 54.655000   8.840000 ;
      RECT 53.815000   8.840000 54.725000   8.910000 ;
      RECT 53.815000   8.910000 54.795000   8.980000 ;
      RECT 53.815000   8.980000 54.865000   9.050000 ;
      RECT 53.815000   9.050000 54.935000   9.120000 ;
      RECT 53.815000   9.120000 55.005000   9.190000 ;
      RECT 53.815000   9.190000 55.075000   9.260000 ;
      RECT 53.815000   9.260000 55.145000   9.330000 ;
      RECT 53.815000   9.330000 55.215000   9.400000 ;
      RECT 53.815000   9.400000 55.285000   9.470000 ;
      RECT 53.815000   9.470000 55.355000   9.540000 ;
      RECT 53.815000   9.540000 55.425000   9.610000 ;
      RECT 53.815000   9.610000 55.495000   9.680000 ;
      RECT 53.815000   9.680000 55.565000   9.750000 ;
      RECT 53.815000   9.750000 55.635000   9.800000 ;
      RECT 55.875000   9.800000 56.110000  10.030000 ;
      RECT 55.875000  10.030000 56.110000  17.360000 ;
      RECT 68.150000  74.490000 75.000000  98.700000 ;
      RECT 68.150000 130.845000 75.000000 133.770000 ;
      RECT 68.150000 140.850000 75.000000 143.770000 ;
      RECT 68.150000 150.850000 75.000000 153.770000 ;
      RECT 68.150000 160.850000 75.000000 163.770000 ;
      RECT 68.150000 170.850000 75.000000 173.770000 ;
      RECT 68.150000 180.850000 75.000000 183.770000 ;
      RECT 68.150000 190.850000 75.000000 193.770000 ;
      RECT 68.290000  74.545000 75.000000  98.840000 ;
      RECT 68.290000 130.705000 75.000000 133.910000 ;
      RECT 68.290000 140.710000 75.000000 143.910000 ;
      RECT 68.290000 150.710000 75.000000 153.910000 ;
      RECT 68.290000 160.710000 75.000000 163.910000 ;
      RECT 68.290000 170.710000 75.000000 173.910000 ;
      RECT 68.290000 180.710000 75.000000 183.910000 ;
      RECT 68.290000 190.710000 75.000000 193.910000 ;
      RECT 68.295000  74.540000 75.000000  74.545000 ;
      RECT 68.295000  74.540000 75.000000  74.545000 ;
      RECT 68.365000  74.470000 75.000000  74.540000 ;
      RECT 68.365000  74.470000 75.000000  74.540000 ;
      RECT 68.435000  74.400000 75.000000  74.470000 ;
      RECT 68.435000  74.400000 75.000000  74.470000 ;
      RECT 68.505000  74.330000 75.000000  74.400000 ;
      RECT 68.505000  74.330000 75.000000  74.400000 ;
      RECT 68.575000  74.260000 75.000000  74.330000 ;
      RECT 68.575000  74.260000 75.000000  74.330000 ;
      RECT 68.645000  74.190000 75.000000  74.260000 ;
      RECT 68.645000  74.190000 75.000000  74.260000 ;
      RECT 68.715000  74.120000 75.000000  74.190000 ;
      RECT 68.715000  74.120000 75.000000  74.190000 ;
      RECT 68.785000  74.050000 75.000000  74.120000 ;
      RECT 68.785000  74.050000 75.000000  74.120000 ;
      RECT 68.855000  73.980000 75.000000  74.050000 ;
      RECT 68.855000  73.980000 75.000000  74.050000 ;
      RECT 68.865000  73.770000 75.000000  74.490000 ;
      RECT 68.925000  73.910000 75.000000  73.980000 ;
      RECT 68.925000  73.910000 75.000000  73.980000 ;
      RECT 74.840000   0.000000 75.000000  73.770000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.200000 171.495000 ;
      RECT  0.000000 171.495000 15.205000 189.915000 ;
      RECT  0.000000 171.595000 15.205000 189.915000 ;
      RECT  0.000000 189.915000 75.000000 198.000000 ;
      RECT  0.000000 189.915000 75.000000 198.000000 ;
      RECT 13.200000  94.385000 15.205000 171.495000 ;
      RECT 13.300000  94.425000 15.205000 171.595000 ;
      RECT 13.440000  94.145000 15.205000  94.385000 ;
      RECT 13.440000  94.285000 15.205000  94.425000 ;
      RECT 13.580000  94.145000 15.205000  94.285000 ;
      RECT 13.725000  94.000000 15.205000  94.145000 ;
      RECT 13.875000  93.850000 15.350000  94.000000 ;
      RECT 14.025000  93.700000 15.500000  93.850000 ;
      RECT 14.175000  93.550000 15.650000  93.700000 ;
      RECT 14.325000  93.400000 15.800000  93.550000 ;
      RECT 14.475000  93.250000 15.950000  93.400000 ;
      RECT 14.625000  93.100000 16.100000  93.250000 ;
      RECT 14.775000  92.950000 16.250000  93.100000 ;
      RECT 14.925000  92.800000 16.400000  92.950000 ;
      RECT 15.075000  92.650000 16.550000  92.800000 ;
      RECT 15.225000  92.500000 16.700000  92.650000 ;
      RECT 15.375000  92.350000 16.850000  92.500000 ;
      RECT 15.525000  92.200000 17.000000  92.350000 ;
      RECT 15.675000  92.050000 17.150000  92.200000 ;
      RECT 15.825000  91.900000 17.300000  92.050000 ;
      RECT 15.975000  91.750000 17.450000  91.900000 ;
      RECT 16.125000  91.600000 17.600000  91.750000 ;
      RECT 16.275000  91.450000 17.750000  91.600000 ;
      RECT 16.425000  91.300000 17.900000  91.450000 ;
      RECT 16.575000  91.150000 18.050000  91.300000 ;
      RECT 16.725000  91.000000 18.200000  91.150000 ;
      RECT 16.875000  90.850000 18.350000  91.000000 ;
      RECT 17.025000  90.700000 18.500000  90.850000 ;
      RECT 17.175000  90.550000 18.650000  90.700000 ;
      RECT 17.325000  90.400000 18.800000  90.550000 ;
      RECT 17.475000  90.250000 18.950000  90.400000 ;
      RECT 17.625000  90.100000 19.100000  90.250000 ;
      RECT 17.775000  89.950000 19.250000  90.100000 ;
      RECT 17.925000  89.800000 19.400000  89.950000 ;
      RECT 18.075000  89.650000 19.550000  89.800000 ;
      RECT 18.225000  89.500000 19.700000  89.650000 ;
      RECT 18.375000  89.350000 19.850000  89.500000 ;
      RECT 18.525000  89.200000 20.000000  89.350000 ;
      RECT 18.675000  89.050000 20.150000  89.200000 ;
      RECT 18.825000  88.900000 20.300000  89.050000 ;
      RECT 18.975000  88.750000 20.450000  88.900000 ;
      RECT 19.125000  88.600000 20.600000  88.750000 ;
      RECT 19.275000  88.450000 20.750000  88.600000 ;
      RECT 19.425000  88.300000 20.900000  88.450000 ;
      RECT 19.575000  88.150000 21.050000  88.300000 ;
      RECT 19.725000  88.000000 21.200000  88.150000 ;
      RECT 19.875000  87.850000 21.350000  88.000000 ;
      RECT 20.025000  87.700000 21.500000  87.850000 ;
      RECT 20.175000  87.550000 21.650000  87.700000 ;
      RECT 20.325000  87.400000 21.800000  87.550000 ;
      RECT 20.475000  87.250000 21.950000  87.400000 ;
      RECT 20.625000  87.100000 22.100000  87.250000 ;
      RECT 20.775000  86.950000 22.250000  87.100000 ;
      RECT 20.925000  86.800000 22.400000  86.950000 ;
      RECT 21.075000  86.650000 22.550000  86.800000 ;
      RECT 21.225000  86.500000 22.700000  86.650000 ;
      RECT 21.375000  86.350000 22.850000  86.500000 ;
      RECT 21.525000  86.200000 23.000000  86.350000 ;
      RECT 21.675000  86.050000 23.150000  86.200000 ;
      RECT 21.825000  85.900000 23.300000  86.050000 ;
      RECT 21.950000  85.775000 23.450000  85.900000 ;
      RECT 22.005000  96.955000 25.635000 166.935000 ;
      RECT 22.005000  96.955000 25.635000 166.935000 ;
      RECT 22.005000 166.935000 25.635000 170.445000 ;
      RECT 22.075000  96.885000 25.635000  96.955000 ;
      RECT 22.100000  85.625000 23.450000  85.775000 ;
      RECT 22.155000 166.935000 25.635000 167.085000 ;
      RECT 22.225000  96.735000 25.635000  96.885000 ;
      RECT 22.250000  85.475000 23.450000  85.625000 ;
      RECT 22.305000 167.085000 25.635000 167.235000 ;
      RECT 22.375000  96.585000 25.635000  96.735000 ;
      RECT 22.400000  85.325000 23.450000  85.475000 ;
      RECT 22.455000 167.235000 25.635000 167.385000 ;
      RECT 22.525000  96.435000 25.635000  96.585000 ;
      RECT 22.550000  85.175000 23.450000  85.325000 ;
      RECT 22.605000 167.385000 25.635000 167.535000 ;
      RECT 22.675000  96.285000 25.635000  96.435000 ;
      RECT 22.700000  85.025000 23.450000  85.175000 ;
      RECT 22.755000 167.535000 25.635000 167.685000 ;
      RECT 22.825000  96.135000 25.635000  96.285000 ;
      RECT 22.850000  84.875000 23.450000  85.025000 ;
      RECT 22.905000 167.685000 25.635000 167.835000 ;
      RECT 22.975000  95.985000 25.635000  96.135000 ;
      RECT 23.000000  84.725000 23.450000  84.875000 ;
      RECT 23.055000 167.835000 25.635000 167.985000 ;
      RECT 23.100000  84.485000 23.450000  85.900000 ;
      RECT 23.125000  95.835000 25.635000  95.985000 ;
      RECT 23.150000  84.575000 23.450000  84.725000 ;
      RECT 23.205000 167.985000 25.635000 168.135000 ;
      RECT 23.275000  95.685000 25.635000  95.835000 ;
      RECT 23.300000  84.425000 23.450000  84.575000 ;
      RECT 23.355000 168.135000 25.635000 168.285000 ;
      RECT 23.425000  95.535000 25.635000  95.685000 ;
      RECT 23.505000 168.285000 25.635000 168.435000 ;
      RECT 23.575000  95.385000 25.635000  95.535000 ;
      RECT 23.655000 168.435000 25.635000 168.585000 ;
      RECT 23.725000  95.235000 25.635000  95.385000 ;
      RECT 23.805000 168.585000 25.635000 168.735000 ;
      RECT 23.875000  95.085000 25.635000  95.235000 ;
      RECT 23.955000 168.735000 25.635000 168.885000 ;
      RECT 24.025000  94.935000 25.635000  95.085000 ;
      RECT 24.105000 168.885000 25.635000 169.035000 ;
      RECT 24.175000  94.785000 25.635000  94.935000 ;
      RECT 24.255000 169.035000 25.635000 169.185000 ;
      RECT 24.325000  94.635000 25.635000  94.785000 ;
      RECT 24.405000 169.185000 25.635000 169.335000 ;
      RECT 24.475000  94.485000 25.635000  94.635000 ;
      RECT 24.555000 169.335000 25.635000 169.485000 ;
      RECT 24.625000  94.335000 25.635000  94.485000 ;
      RECT 24.625000  94.335000 25.635000  96.955000 ;
      RECT 24.705000 169.485000 25.635000 169.635000 ;
      RECT 24.745000  94.215000 25.635000  94.335000 ;
      RECT 24.800000   0.000000 25.600000  82.335000 ;
      RECT 24.800000  82.335000 25.150000  82.785000 ;
      RECT 24.855000 169.635000 25.635000 169.785000 ;
      RECT 24.895000  94.065000 25.755000  94.215000 ;
      RECT 24.900000   0.000000 25.600000  82.335000 ;
      RECT 24.900000  82.335000 25.450000  82.485000 ;
      RECT 24.900000  82.485000 25.300000  82.635000 ;
      RECT 24.900000  82.635000 25.150000  82.785000 ;
      RECT 24.900000  82.785000 25.000000  82.935000 ;
      RECT 25.005000 169.785000 25.635000 169.935000 ;
      RECT 25.045000  93.915000 25.905000  94.065000 ;
      RECT 25.155000 169.935000 25.635000 170.085000 ;
      RECT 25.195000  93.765000 26.055000  93.915000 ;
      RECT 25.305000 170.085000 25.635000 170.235000 ;
      RECT 25.345000  93.615000 26.205000  93.765000 ;
      RECT 25.455000 170.235000 25.635000 170.385000 ;
      RECT 25.495000  93.465000 26.355000  93.615000 ;
      RECT 25.515000 170.445000 25.635000 189.915000 ;
      RECT 25.605000 170.385000 25.635000 170.535000 ;
      RECT 25.645000  93.315000 26.505000  93.465000 ;
      RECT 25.795000  93.165000 26.655000  93.315000 ;
      RECT 25.945000  93.015000 26.805000  93.165000 ;
      RECT 26.095000  92.865000 26.955000  93.015000 ;
      RECT 26.245000  92.715000 27.105000  92.865000 ;
      RECT 26.395000  92.565000 27.255000  92.715000 ;
      RECT 26.545000  92.415000 27.405000  92.565000 ;
      RECT 26.695000  92.265000 27.555000  92.415000 ;
      RECT 26.845000  92.115000 27.705000  92.265000 ;
      RECT 26.995000  91.965000 27.855000  92.115000 ;
      RECT 27.145000  91.815000 28.005000  91.965000 ;
      RECT 27.295000  91.665000 28.155000  91.815000 ;
      RECT 27.445000  91.515000 28.305000  91.665000 ;
      RECT 27.595000  91.365000 28.455000  91.515000 ;
      RECT 27.745000  91.215000 28.605000  91.365000 ;
      RECT 27.895000  91.065000 28.755000  91.215000 ;
      RECT 28.045000  90.915000 28.905000  91.065000 ;
      RECT 28.195000  90.765000 29.055000  90.915000 ;
      RECT 28.345000  90.615000 29.205000  90.765000 ;
      RECT 28.495000  90.465000 29.355000  90.615000 ;
      RECT 28.645000  90.315000 29.505000  90.465000 ;
      RECT 28.795000  90.165000 29.655000  90.315000 ;
      RECT 28.945000  90.015000 29.805000  90.165000 ;
      RECT 29.095000  89.865000 29.955000  90.015000 ;
      RECT 29.245000  89.715000 30.105000  89.865000 ;
      RECT 29.395000  89.565000 30.255000  89.715000 ;
      RECT 29.545000  89.415000 30.405000  89.565000 ;
      RECT 29.695000  89.265000 30.555000  89.415000 ;
      RECT 29.845000  89.115000 30.705000  89.265000 ;
      RECT 29.995000  88.965000 30.855000  89.115000 ;
      RECT 30.145000  88.815000 31.005000  88.965000 ;
      RECT 30.295000  88.665000 31.155000  88.815000 ;
      RECT 30.445000  88.515000 31.305000  88.665000 ;
      RECT 30.595000  88.365000 31.455000  88.515000 ;
      RECT 30.745000  88.215000 31.605000  88.365000 ;
      RECT 30.895000  88.065000 31.755000  88.215000 ;
      RECT 31.045000  87.915000 31.905000  88.065000 ;
      RECT 31.195000  87.765000 32.055000  87.915000 ;
      RECT 31.345000  87.615000 32.205000  87.765000 ;
      RECT 31.495000  87.465000 32.355000  87.615000 ;
      RECT 31.645000  87.315000 32.505000  87.465000 ;
      RECT 31.795000  87.165000 32.655000  87.315000 ;
      RECT 31.945000  87.015000 32.805000  87.165000 ;
      RECT 32.095000  86.865000 32.955000  87.015000 ;
      RECT 32.245000  86.715000 33.105000  86.865000 ;
      RECT 32.395000  86.565000 33.255000  86.715000 ;
      RECT 32.435000  93.555000 40.410000  93.705000 ;
      RECT 32.435000  93.555000 42.435000  95.580000 ;
      RECT 32.435000  93.705000 40.560000  93.855000 ;
      RECT 32.435000  93.855000 40.710000  94.005000 ;
      RECT 32.435000  94.005000 40.860000  94.155000 ;
      RECT 32.435000  94.155000 41.010000  94.305000 ;
      RECT 32.435000  94.305000 41.160000  94.455000 ;
      RECT 32.435000  94.455000 41.310000  94.605000 ;
      RECT 32.435000  94.605000 41.460000  94.755000 ;
      RECT 32.435000  94.755000 41.610000  94.905000 ;
      RECT 32.435000  94.905000 41.760000  95.055000 ;
      RECT 32.435000  95.055000 41.910000  95.205000 ;
      RECT 32.435000  95.205000 42.060000  95.355000 ;
      RECT 32.435000  95.355000 42.210000  95.505000 ;
      RECT 32.435000  95.505000 42.360000  95.580000 ;
      RECT 32.435000  95.580000 42.435000 162.405000 ;
      RECT 32.435000  95.580000 42.435000 162.405000 ;
      RECT 32.435000 162.405000 42.435000 163.970000 ;
      RECT 32.515000  93.475000 40.330000  93.555000 ;
      RECT 32.545000  84.855000 34.105000  85.865000 ;
      RECT 32.545000  84.855000 34.105000  85.865000 ;
      RECT 32.545000  85.865000 33.555000  86.415000 ;
      RECT 32.545000  85.865000 33.955000  86.015000 ;
      RECT 32.545000  86.015000 33.805000  86.165000 ;
      RECT 32.545000  86.165000 33.655000  86.315000 ;
      RECT 32.545000  86.315000 33.555000  86.415000 ;
      RECT 32.545000  86.415000 33.405000  86.565000 ;
      RECT 32.570000  84.830000 34.080000  84.855000 ;
      RECT 32.585000 162.405000 42.435000 162.555000 ;
      RECT 32.665000  93.325000 40.180000  93.475000 ;
      RECT 32.720000  84.680000 33.930000  84.830000 ;
      RECT 32.735000 162.555000 42.435000 162.705000 ;
      RECT 32.815000  93.175000 40.030000  93.325000 ;
      RECT 32.870000  84.530000 33.780000  84.680000 ;
      RECT 32.885000 162.705000 42.435000 162.855000 ;
      RECT 32.965000  93.025000 39.880000  93.175000 ;
      RECT 33.020000  84.380000 33.630000  84.530000 ;
      RECT 33.020000  84.380000 34.105000  84.855000 ;
      RECT 33.035000 162.855000 42.435000 163.005000 ;
      RECT 33.115000  92.875000 39.730000  93.025000 ;
      RECT 33.185000 163.005000 42.435000 163.155000 ;
      RECT 33.265000  92.725000 39.580000  92.875000 ;
      RECT 33.335000 163.155000 42.435000 163.305000 ;
      RECT 33.415000  92.575000 39.430000  92.725000 ;
      RECT 33.485000 163.305000 42.435000 163.455000 ;
      RECT 33.565000  92.425000 39.280000  92.575000 ;
      RECT 33.635000 163.455000 42.435000 163.605000 ;
      RECT 33.715000  92.275000 39.130000  92.425000 ;
      RECT 33.785000 163.605000 42.435000 163.755000 ;
      RECT 33.865000  92.125000 38.980000  92.275000 ;
      RECT 33.935000 163.755000 42.435000 163.905000 ;
      RECT 34.000000 163.905000 42.435000 163.970000 ;
      RECT 34.000000 163.970000 39.110000 167.295000 ;
      RECT 34.015000  91.975000 38.830000  92.125000 ;
      RECT 34.150000 163.970000 42.285000 164.120000 ;
      RECT 34.165000  91.825000 38.680000  91.975000 ;
      RECT 34.300000 164.120000 42.135000 164.270000 ;
      RECT 34.315000  91.675000 38.530000  91.825000 ;
      RECT 34.450000 164.270000 41.985000 164.420000 ;
      RECT 34.465000  91.525000 38.380000  91.675000 ;
      RECT 34.600000 164.420000 41.835000 164.570000 ;
      RECT 34.615000  91.375000 38.230000  91.525000 ;
      RECT 34.750000 164.570000 41.685000 164.720000 ;
      RECT 34.765000  91.225000 38.080000  91.375000 ;
      RECT 34.900000 164.720000 41.535000 164.870000 ;
      RECT 34.915000  91.075000 37.930000  91.225000 ;
      RECT 35.050000 164.870000 41.385000 165.020000 ;
      RECT 35.065000  90.925000 37.780000  91.075000 ;
      RECT 35.200000 165.020000 41.235000 165.170000 ;
      RECT 35.215000  90.775000 37.630000  90.925000 ;
      RECT 35.215000  90.775000 40.410000  93.555000 ;
      RECT 35.350000 165.170000 41.085000 165.320000 ;
      RECT 35.500000 165.320000 40.935000 165.470000 ;
      RECT 35.650000 165.470000 40.785000 165.620000 ;
      RECT 35.800000 165.620000 40.635000 165.770000 ;
      RECT 35.950000 165.770000 40.485000 165.920000 ;
      RECT 36.100000 165.920000 40.335000 166.070000 ;
      RECT 36.250000 166.070000 40.185000 166.220000 ;
      RECT 36.400000 166.220000 40.035000 166.370000 ;
      RECT 36.550000 166.370000 39.885000 166.520000 ;
      RECT 36.700000 166.520000 39.735000 166.670000 ;
      RECT 36.850000 166.670000 39.585000 166.820000 ;
      RECT 37.000000 166.820000 39.435000 166.970000 ;
      RECT 37.150000 166.970000 39.285000 167.120000 ;
      RECT 37.280000   0.000000 37.980000  69.890000 ;
      RECT 37.280000   0.000000 37.980000  69.890000 ;
      RECT 37.280000  69.890000 50.355000  70.940000 ;
      RECT 37.280000  69.890000 50.455000  70.940000 ;
      RECT 37.280000  70.940000 50.455000  74.340000 ;
      RECT 37.300000 167.120000 39.135000 167.270000 ;
      RECT 37.325000 167.270000 39.110000 167.295000 ;
      RECT 37.325000 167.295000 37.545000 168.860000 ;
      RECT 37.325000 167.295000 38.960000 167.445000 ;
      RECT 37.325000 167.445000 38.810000 167.595000 ;
      RECT 37.325000 167.595000 38.660000 167.745000 ;
      RECT 37.325000 167.745000 38.510000 167.895000 ;
      RECT 37.325000 167.895000 38.360000 168.045000 ;
      RECT 37.325000 168.045000 38.210000 168.195000 ;
      RECT 37.325000 168.195000 38.060000 168.345000 ;
      RECT 37.325000 168.345000 37.910000 168.495000 ;
      RECT 37.325000 168.495000 37.760000 168.645000 ;
      RECT 37.325000 168.645000 37.610000 168.795000 ;
      RECT 37.325000 168.795000 37.460000 168.945000 ;
      RECT 37.325000 168.860000 37.545000 189.915000 ;
      RECT 37.430000  70.940000 50.355000  71.090000 ;
      RECT 37.430000  70.940000 50.355000  71.090000 ;
      RECT 37.580000  71.090000 50.355000  71.240000 ;
      RECT 37.580000  71.090000 50.355000  71.240000 ;
      RECT 37.730000  71.240000 50.355000  71.390000 ;
      RECT 37.730000  71.240000 50.355000  71.390000 ;
      RECT 37.880000  71.390000 50.355000  71.540000 ;
      RECT 37.880000  71.390000 50.355000  71.540000 ;
      RECT 38.030000  71.540000 50.355000  71.690000 ;
      RECT 38.030000  71.540000 50.355000  71.690000 ;
      RECT 38.180000  71.690000 50.355000  71.840000 ;
      RECT 38.180000  71.690000 50.355000  71.840000 ;
      RECT 38.330000  71.840000 50.355000  71.990000 ;
      RECT 38.330000  71.840000 50.355000  71.990000 ;
      RECT 38.480000  71.990000 50.355000  72.140000 ;
      RECT 38.480000  71.990000 50.355000  72.140000 ;
      RECT 38.630000  72.140000 50.355000  72.290000 ;
      RECT 38.630000  72.140000 50.355000  72.290000 ;
      RECT 38.780000  72.290000 50.355000  72.440000 ;
      RECT 38.780000  72.290000 50.355000  72.440000 ;
      RECT 38.930000  72.440000 50.355000  72.590000 ;
      RECT 38.930000  72.440000 50.355000  72.590000 ;
      RECT 39.080000  72.590000 50.355000  72.740000 ;
      RECT 39.080000  72.590000 50.355000  72.740000 ;
      RECT 39.230000  72.740000 50.355000  72.890000 ;
      RECT 39.230000  72.740000 50.355000  72.890000 ;
      RECT 39.380000  72.890000 50.355000  73.040000 ;
      RECT 39.380000  72.890000 50.355000  73.040000 ;
      RECT 39.530000  73.040000 50.355000  73.190000 ;
      RECT 39.530000  73.040000 50.355000  73.190000 ;
      RECT 39.680000  73.190000 50.355000  73.340000 ;
      RECT 39.680000  73.190000 50.355000  73.340000 ;
      RECT 39.785000  84.855000 41.210000  87.195000 ;
      RECT 39.785000  84.855000 41.210000  87.195000 ;
      RECT 39.785000  87.195000 41.210000  87.610000 ;
      RECT 39.810000  84.830000 41.185000  84.855000 ;
      RECT 39.830000  73.340000 50.355000  73.490000 ;
      RECT 39.830000  73.340000 50.355000  73.490000 ;
      RECT 39.935000  87.195000 41.210000  87.345000 ;
      RECT 39.960000  84.680000 41.035000  84.830000 ;
      RECT 39.980000  73.490000 50.355000  73.640000 ;
      RECT 39.980000  73.490000 50.355000  73.640000 ;
      RECT 40.085000  87.345000 41.210000  87.495000 ;
      RECT 40.110000  84.530000 40.885000  84.680000 ;
      RECT 40.130000  73.640000 50.355000  73.790000 ;
      RECT 40.130000  73.640000 50.355000  73.790000 ;
      RECT 40.200000  87.495000 41.210000  87.610000 ;
      RECT 40.200000  87.610000 50.245000  96.645000 ;
      RECT 40.260000  84.380000 40.735000  84.530000 ;
      RECT 40.260000  84.380000 41.210000  84.855000 ;
      RECT 40.280000  73.790000 50.355000  73.940000 ;
      RECT 40.280000  73.790000 50.355000  73.940000 ;
      RECT 40.350000  87.610000 41.210000  87.760000 ;
      RECT 40.430000  73.940000 50.355000  74.090000 ;
      RECT 40.430000  73.940000 50.355000  74.090000 ;
      RECT 40.500000  87.760000 41.360000  87.910000 ;
      RECT 40.580000  74.090000 50.355000  74.240000 ;
      RECT 40.580000  74.090000 50.355000  74.240000 ;
      RECT 40.650000  87.910000 41.510000  88.060000 ;
      RECT 40.680000  74.240000 50.355000  74.340000 ;
      RECT 40.680000  74.240000 50.355000  74.340000 ;
      RECT 40.800000  88.060000 41.660000  88.210000 ;
      RECT 40.950000  88.210000 41.810000  88.360000 ;
      RECT 41.100000  88.360000 41.960000  88.510000 ;
      RECT 41.250000  88.510000 42.110000  88.660000 ;
      RECT 41.400000  88.660000 42.260000  88.810000 ;
      RECT 41.550000  88.810000 42.410000  88.960000 ;
      RECT 41.700000  88.960000 42.560000  89.110000 ;
      RECT 41.850000  89.110000 42.710000  89.260000 ;
      RECT 42.000000  89.260000 42.860000  89.410000 ;
      RECT 42.150000  89.410000 43.010000  89.560000 ;
      RECT 42.300000  89.560000 43.160000  89.710000 ;
      RECT 42.450000  89.710000 43.310000  89.860000 ;
      RECT 42.600000  89.860000 43.460000  90.010000 ;
      RECT 42.750000  90.010000 43.610000  90.160000 ;
      RECT 42.900000  90.160000 43.760000  90.310000 ;
      RECT 43.050000  90.310000 43.910000  90.460000 ;
      RECT 43.200000  90.460000 44.060000  90.610000 ;
      RECT 43.350000  90.610000 44.210000  90.760000 ;
      RECT 43.500000  90.760000 44.360000  90.910000 ;
      RECT 43.650000  90.910000 44.510000  91.060000 ;
      RECT 43.800000  91.060000 44.660000  91.210000 ;
      RECT 43.950000  91.210000 44.810000  91.360000 ;
      RECT 44.100000  91.360000 44.960000  91.510000 ;
      RECT 44.250000  91.510000 45.110000  91.660000 ;
      RECT 44.400000  91.660000 45.260000  91.810000 ;
      RECT 44.550000  91.810000 45.410000  91.960000 ;
      RECT 44.700000  91.960000 45.560000  92.110000 ;
      RECT 44.850000  92.110000 45.710000  92.260000 ;
      RECT 45.000000  92.260000 45.860000  92.410000 ;
      RECT 45.150000  92.410000 46.010000  92.560000 ;
      RECT 45.300000  92.560000 46.160000  92.710000 ;
      RECT 45.450000  92.710000 46.310000  92.860000 ;
      RECT 45.600000  92.860000 46.460000  93.010000 ;
      RECT 45.750000  93.010000 46.610000  93.160000 ;
      RECT 45.900000  93.160000 46.760000  93.310000 ;
      RECT 46.050000  93.310000 46.910000  93.460000 ;
      RECT 46.200000  93.460000 47.060000  93.610000 ;
      RECT 46.350000  93.610000 47.210000  93.760000 ;
      RECT 46.500000  93.760000 47.360000  93.910000 ;
      RECT 46.650000  93.910000 47.510000  94.060000 ;
      RECT 46.800000  94.060000 47.660000  94.210000 ;
      RECT 46.950000  94.210000 47.810000  94.360000 ;
      RECT 46.960000  74.340000 50.455000  76.650000 ;
      RECT 47.100000  94.360000 47.960000  94.510000 ;
      RECT 47.110000  74.340000 50.355000  74.490000 ;
      RECT 47.110000  74.340000 50.355000  74.490000 ;
      RECT 47.250000  94.510000 48.110000  94.660000 ;
      RECT 47.260000  74.490000 50.355000  74.640000 ;
      RECT 47.260000  74.490000 50.355000  74.640000 ;
      RECT 47.400000  94.660000 48.260000  94.810000 ;
      RECT 47.410000  74.640000 50.355000  74.790000 ;
      RECT 47.410000  74.640000 50.355000  74.790000 ;
      RECT 47.550000  94.810000 48.410000  94.960000 ;
      RECT 47.560000  74.790000 50.355000  74.940000 ;
      RECT 47.560000  74.790000 50.355000  74.940000 ;
      RECT 47.700000  94.960000 48.560000  95.110000 ;
      RECT 47.710000  74.940000 50.355000  75.090000 ;
      RECT 47.710000  74.940000 50.355000  75.090000 ;
      RECT 47.850000  95.110000 48.710000  95.260000 ;
      RECT 47.860000  75.090000 50.355000  75.240000 ;
      RECT 47.860000  75.090000 50.355000  75.240000 ;
      RECT 48.000000  95.260000 48.860000  95.410000 ;
      RECT 48.010000  75.240000 50.355000  75.390000 ;
      RECT 48.010000  75.240000 50.355000  75.390000 ;
      RECT 48.150000  95.410000 49.010000  95.560000 ;
      RECT 48.160000  75.390000 50.355000  75.540000 ;
      RECT 48.160000  75.390000 50.355000  75.540000 ;
      RECT 48.300000  95.560000 49.160000  95.710000 ;
      RECT 48.310000  75.540000 50.355000  75.690000 ;
      RECT 48.310000  75.540000 50.355000  75.690000 ;
      RECT 48.450000  95.710000 49.310000  95.860000 ;
      RECT 48.460000  75.690000 50.355000  75.840000 ;
      RECT 48.460000  75.690000 50.355000  75.840000 ;
      RECT 48.600000  95.860000 49.460000  96.010000 ;
      RECT 48.610000  75.840000 50.355000  75.990000 ;
      RECT 48.610000  75.840000 50.355000  75.990000 ;
      RECT 48.750000  96.010000 49.610000  96.160000 ;
      RECT 48.760000  75.990000 50.355000  76.140000 ;
      RECT 48.760000  75.990000 50.355000  76.140000 ;
      RECT 48.900000  96.160000 49.760000  96.310000 ;
      RECT 48.910000  76.140000 50.355000  76.290000 ;
      RECT 48.910000  76.140000 50.355000  76.290000 ;
      RECT 49.050000  96.310000 49.910000  96.460000 ;
      RECT 49.060000  76.290000 50.355000  76.440000 ;
      RECT 49.060000  76.290000 50.355000  76.440000 ;
      RECT 49.200000  96.460000 50.060000  96.610000 ;
      RECT 49.210000  76.440000 50.355000  76.590000 ;
      RECT 49.210000  76.440000 50.355000  76.590000 ;
      RECT 49.235000  96.610000 50.210000  96.645000 ;
      RECT 49.235000  96.645000 50.245000  96.795000 ;
      RECT 49.235000  96.645000 53.930000 100.330000 ;
      RECT 49.235000  96.795000 50.395000  96.945000 ;
      RECT 49.235000  96.945000 50.545000  97.095000 ;
      RECT 49.235000  97.095000 50.695000  97.245000 ;
      RECT 49.235000  97.245000 50.845000  97.395000 ;
      RECT 49.235000  97.395000 50.995000  97.545000 ;
      RECT 49.235000  97.545000 51.145000  97.695000 ;
      RECT 49.235000  97.695000 51.295000  97.845000 ;
      RECT 49.235000  97.845000 51.445000  97.995000 ;
      RECT 49.235000  97.995000 51.595000  98.145000 ;
      RECT 49.235000  98.145000 51.745000  98.295000 ;
      RECT 49.235000  98.295000 51.895000  98.445000 ;
      RECT 49.235000  98.445000 52.045000  98.595000 ;
      RECT 49.235000  98.595000 52.195000  98.745000 ;
      RECT 49.235000  98.745000 52.345000  98.895000 ;
      RECT 49.235000  98.895000 52.495000  99.045000 ;
      RECT 49.235000  99.045000 52.645000  99.195000 ;
      RECT 49.235000  99.195000 52.795000  99.345000 ;
      RECT 49.235000  99.345000 52.945000  99.495000 ;
      RECT 49.235000  99.495000 53.095000  99.645000 ;
      RECT 49.235000  99.645000 53.245000  99.795000 ;
      RECT 49.235000  99.795000 53.395000  99.945000 ;
      RECT 49.235000  99.945000 53.545000 100.095000 ;
      RECT 49.235000 100.095000 53.695000 100.245000 ;
      RECT 49.235000 100.245000 53.845000 100.330000 ;
      RECT 49.235000 100.330000 53.930000 164.295000 ;
      RECT 49.235000 100.330000 53.930000 164.295000 ;
      RECT 49.235000 164.295000 49.470000 168.755000 ;
      RECT 49.235000 164.295000 53.780000 164.445000 ;
      RECT 49.235000 164.445000 53.630000 164.595000 ;
      RECT 49.235000 164.595000 53.480000 164.745000 ;
      RECT 49.235000 164.745000 53.330000 164.895000 ;
      RECT 49.235000 164.895000 53.180000 165.045000 ;
      RECT 49.235000 165.045000 53.030000 165.195000 ;
      RECT 49.235000 165.195000 52.880000 165.345000 ;
      RECT 49.235000 165.345000 52.730000 165.495000 ;
      RECT 49.235000 165.495000 52.580000 165.645000 ;
      RECT 49.235000 165.645000 52.430000 165.795000 ;
      RECT 49.235000 165.795000 52.280000 165.945000 ;
      RECT 49.235000 165.945000 52.130000 166.095000 ;
      RECT 49.235000 166.095000 51.980000 166.245000 ;
      RECT 49.235000 166.245000 51.830000 166.395000 ;
      RECT 49.235000 166.395000 51.680000 166.545000 ;
      RECT 49.235000 166.545000 51.530000 166.695000 ;
      RECT 49.235000 166.695000 51.380000 166.845000 ;
      RECT 49.235000 166.845000 51.230000 166.995000 ;
      RECT 49.235000 166.995000 51.080000 167.145000 ;
      RECT 49.235000 167.145000 50.930000 167.295000 ;
      RECT 49.235000 167.295000 50.780000 167.445000 ;
      RECT 49.235000 167.445000 50.630000 167.595000 ;
      RECT 49.235000 167.595000 50.480000 167.745000 ;
      RECT 49.235000 167.745000 50.330000 167.895000 ;
      RECT 49.235000 167.895000 50.180000 168.045000 ;
      RECT 49.235000 168.045000 50.030000 168.195000 ;
      RECT 49.235000 168.195000 49.880000 168.345000 ;
      RECT 49.235000 168.345000 49.730000 168.495000 ;
      RECT 49.235000 168.495000 49.580000 168.645000 ;
      RECT 49.235000 168.645000 49.430000 168.795000 ;
      RECT 49.235000 168.755000 49.470000 189.915000 ;
      RECT 49.235000 168.795000 49.280000 168.945000 ;
      RECT 49.270000  76.590000 50.355000  76.650000 ;
      RECT 49.270000  76.590000 50.355000  76.650000 ;
      RECT 49.270000  76.650000 50.455000  84.590000 ;
      RECT 49.270000  77.735000 50.355000  84.630000 ;
      RECT 49.270000  84.590000 50.510000  84.645000 ;
      RECT 49.270000  84.630000 50.355000  84.635000 ;
      RECT 49.270000  84.635000 50.360000  84.640000 ;
      RECT 49.270000  84.640000 50.365000  84.645000 ;
      RECT 49.270000  84.645000 52.660000  86.795000 ;
      RECT 49.420000  76.650000 50.355000  76.800000 ;
      RECT 49.420000  76.650000 50.355000  76.800000 ;
      RECT 49.420000  84.645000 50.370000  84.795000 ;
      RECT 49.570000  76.800000 50.355000  76.950000 ;
      RECT 49.570000  76.800000 50.355000  76.950000 ;
      RECT 49.570000  84.795000 50.520000  84.945000 ;
      RECT 49.655000   0.000000 50.355000  69.890000 ;
      RECT 49.655000   0.000000 50.455000  69.890000 ;
      RECT 49.720000  76.950000 50.355000  77.100000 ;
      RECT 49.720000  76.950000 50.355000  77.100000 ;
      RECT 49.720000  84.945000 50.670000  85.095000 ;
      RECT 49.870000  77.100000 50.355000  77.250000 ;
      RECT 49.870000  77.100000 50.355000  77.250000 ;
      RECT 49.870000  85.095000 50.820000  85.245000 ;
      RECT 50.020000  77.250000 50.355000  77.400000 ;
      RECT 50.020000  77.250000 50.355000  77.400000 ;
      RECT 50.020000  85.245000 50.970000  85.395000 ;
      RECT 50.170000  77.400000 50.355000  77.550000 ;
      RECT 50.170000  77.400000 50.355000  77.550000 ;
      RECT 50.170000  85.395000 51.120000  85.545000 ;
      RECT 50.320000  77.550000 50.355000  77.700000 ;
      RECT 50.320000  77.550000 50.355000  77.700000 ;
      RECT 50.320000  85.545000 51.270000  85.695000 ;
      RECT 50.470000  85.695000 51.420000  85.845000 ;
      RECT 50.620000  85.845000 51.570000  85.995000 ;
      RECT 50.770000  85.995000 51.720000  86.145000 ;
      RECT 50.920000  86.145000 51.870000  86.295000 ;
      RECT 51.070000  86.295000 52.020000  86.445000 ;
      RECT 51.220000  86.445000 52.170000  86.595000 ;
      RECT 51.370000  86.595000 52.320000  86.745000 ;
      RECT 51.420000  86.745000 52.470000  86.795000 ;
      RECT 51.420000  86.795000 52.520000  86.945000 ;
      RECT 51.420000  86.795000 54.075000  88.210000 ;
      RECT 51.420000  86.945000 52.670000  87.095000 ;
      RECT 51.420000  87.095000 52.820000  87.245000 ;
      RECT 51.420000  87.245000 52.970000  87.395000 ;
      RECT 51.420000  87.395000 53.120000  87.545000 ;
      RECT 51.420000  87.545000 53.270000  87.695000 ;
      RECT 51.420000  87.695000 53.420000  87.845000 ;
      RECT 51.420000  87.845000 53.570000  87.995000 ;
      RECT 51.420000  87.995000 53.720000  88.145000 ;
      RECT 51.420000  88.145000 53.870000  88.210000 ;
      RECT 51.420000  88.210000 61.745000  95.880000 ;
      RECT 51.570000  88.210000 53.935000  88.360000 ;
      RECT 51.720000  88.360000 54.085000  88.510000 ;
      RECT 51.870000  88.510000 54.235000  88.660000 ;
      RECT 52.020000  88.660000 54.385000  88.810000 ;
      RECT 52.170000  88.810000 54.535000  88.960000 ;
      RECT 52.320000  88.960000 54.685000  89.110000 ;
      RECT 52.470000  89.110000 54.835000  89.260000 ;
      RECT 52.620000  89.260000 54.985000  89.410000 ;
      RECT 52.770000  89.410000 55.135000  89.560000 ;
      RECT 52.920000  89.560000 55.285000  89.710000 ;
      RECT 53.070000  89.710000 55.435000  89.860000 ;
      RECT 53.220000  89.860000 55.585000  90.010000 ;
      RECT 53.370000  90.010000 55.735000  90.160000 ;
      RECT 53.520000  90.160000 55.885000  90.310000 ;
      RECT 53.670000  90.310000 56.035000  90.460000 ;
      RECT 53.820000  90.460000 56.185000  90.610000 ;
      RECT 53.970000  90.610000 56.335000  90.760000 ;
      RECT 54.120000  90.760000 56.485000  90.910000 ;
      RECT 54.270000  90.910000 56.635000  91.060000 ;
      RECT 54.420000  91.060000 56.785000  91.210000 ;
      RECT 54.570000  91.210000 56.935000  91.360000 ;
      RECT 54.720000  91.360000 57.085000  91.510000 ;
      RECT 54.870000  91.510000 57.235000  91.660000 ;
      RECT 55.020000  91.660000 57.385000  91.810000 ;
      RECT 55.170000  91.810000 57.535000  91.960000 ;
      RECT 55.320000  91.960000 57.685000  92.110000 ;
      RECT 55.470000  92.110000 57.835000  92.260000 ;
      RECT 55.620000  92.260000 57.985000  92.410000 ;
      RECT 55.770000  92.410000 58.135000  92.560000 ;
      RECT 55.920000  92.560000 58.285000  92.710000 ;
      RECT 56.070000  92.710000 58.435000  92.860000 ;
      RECT 56.220000  92.860000 58.585000  93.010000 ;
      RECT 56.370000  93.010000 58.735000  93.160000 ;
      RECT 56.520000  93.160000 58.885000  93.310000 ;
      RECT 56.670000  93.310000 59.035000  93.460000 ;
      RECT 56.820000  93.460000 59.185000  93.610000 ;
      RECT 56.970000  93.610000 59.335000  93.760000 ;
      RECT 57.120000  93.760000 59.485000  93.910000 ;
      RECT 57.270000  93.910000 59.635000  94.060000 ;
      RECT 57.420000  94.060000 59.785000  94.210000 ;
      RECT 57.570000  94.210000 59.935000  94.360000 ;
      RECT 57.720000  94.360000 60.085000  94.510000 ;
      RECT 57.870000  94.510000 60.235000  94.660000 ;
      RECT 58.020000  94.660000 60.385000  94.810000 ;
      RECT 58.170000  94.810000 60.535000  94.960000 ;
      RECT 58.320000  94.960000 60.685000  95.110000 ;
      RECT 58.470000  95.110000 60.835000  95.260000 ;
      RECT 58.620000  95.260000 60.985000  95.410000 ;
      RECT 58.770000  95.410000 61.135000  95.560000 ;
      RECT 58.920000  95.560000 61.285000  95.710000 ;
      RECT 59.070000  95.710000 61.435000  95.860000 ;
      RECT 59.090000  95.880000 61.745000  97.520000 ;
      RECT 59.130000  95.860000 61.585000  95.920000 ;
      RECT 59.280000  95.920000 61.645000  96.070000 ;
      RECT 59.430000  96.070000 61.645000  96.220000 ;
      RECT 59.580000  96.220000 61.645000  96.370000 ;
      RECT 59.730000  96.370000 61.645000  96.520000 ;
      RECT 59.880000  96.520000 61.645000  96.670000 ;
      RECT 60.030000  96.670000 61.645000  96.820000 ;
      RECT 60.180000  96.820000 61.645000  96.970000 ;
      RECT 60.330000  96.970000 61.645000  97.120000 ;
      RECT 60.480000  97.120000 61.645000  97.270000 ;
      RECT 60.630000  97.270000 61.645000  97.420000 ;
      RECT 60.730000  97.420000 61.645000  97.520000 ;
      RECT 60.730000  97.520000 61.645000 172.635000 ;
      RECT 60.730000  97.520000 61.745000 172.535000 ;
      RECT 60.730000 172.535000 75.000000 189.915000 ;
      RECT 60.730000 172.635000 75.000000 189.915000 ;
    LAYER met4 ;
      RECT  0.000000   5.885000  1.670000   6.485000 ;
      RECT  0.000000   5.885000 75.000000   6.485000 ;
      RECT  0.000000  11.935000  1.365000  12.535000 ;
      RECT  0.000000  11.935000 75.000000  12.535000 ;
      RECT  0.000000  16.785000  1.365000  17.385000 ;
      RECT  0.000000  16.785000 75.000000  17.385000 ;
      RECT  0.000000  22.835000  1.670000  23.435000 ;
      RECT  0.000000  22.835000 75.000000  23.435000 ;
      RECT  0.000000  28.885000  1.670000  29.485000 ;
      RECT  0.000000  28.885000 75.000000  29.485000 ;
      RECT  0.000000  33.735000  1.670000  34.335000 ;
      RECT  0.000000  33.735000 75.000000  34.335000 ;
      RECT  0.000000  38.585000  1.670000  39.185000 ;
      RECT  0.000000  38.585000 75.000000  39.185000 ;
      RECT  0.000000  44.635000  1.670000  45.335000 ;
      RECT  0.000000  44.635000 75.000000  45.435000 ;
      RECT  0.000000  55.035000 75.000000  55.835000 ;
      RECT  0.000000  55.135000  1.670000  55.835000 ;
      RECT  0.000000  61.085000  1.670000  61.685000 ;
      RECT  0.000000  61.085000 75.000000  61.685000 ;
      RECT  0.000000  66.935000  1.670000  67.635000 ;
      RECT  0.000000  66.935000 75.000000  67.635000 ;
      RECT  0.000000  93.400000 75.000000 173.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.570000  45.435000 73.430000  55.035000 ;
      RECT  1.670000   0.000000 73.330000  11.935000 ;
      RECT  1.670000  17.385000 73.330000  93.400000 ;
      RECT  1.670000 173.385000 73.330000 198.000000 ;
      RECT 73.330000   5.885000 75.000000   6.485000 ;
      RECT 73.330000  22.835000 75.000000  23.435000 ;
      RECT 73.330000  28.885000 75.000000  29.485000 ;
      RECT 73.330000  33.735000 75.000000  34.335000 ;
      RECT 73.330000  38.585000 75.000000  39.185000 ;
      RECT 73.330000  44.635000 75.000000  45.335000 ;
      RECT 73.330000  55.135000 75.000000  55.835000 ;
      RECT 73.330000  61.085000 75.000000  61.685000 ;
      RECT 73.330000  66.935000 75.000000  67.635000 ;
      RECT 73.635000  11.935000 75.000000  12.535000 ;
      RECT 73.635000  16.785000 75.000000  17.385000 ;
    LAYER met5 ;
      RECT  0.000000  94.585000 75.000000 161.165000 ;
      RECT  0.000000 161.165000 30.095000 168.720000 ;
      RECT  0.000000 168.720000 75.000000 172.185000 ;
      RECT  2.565000  13.035000 72.435000  16.285000 ;
      RECT  2.870000   0.000000 72.130000  13.035000 ;
      RECT  2.870000  16.285000 72.130000  94.585000 ;
      RECT  2.870000 172.185000 72.130000 198.000000 ;
      RECT 53.940000 161.165000 75.000000 168.720000 ;
  END
END sky130_fd_io__top_power_lvc_wpad


MACRO sky130_fd_io__overlay_vddio_hvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 24.370000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000  1.270000 70.060000 ;
        RECT 0.000000 70.060000 24.400000 90.435000 ;
        RECT 0.000000 90.435000  1.270000 90.630000 ;
        RECT 0.000000 90.630000 19.740000 94.770000 ;
        RECT 0.000000 94.770000  1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.660000 70.060000 75.000000 90.435000 ;
        RECT 55.320000 90.630000 75.000000 94.770000 ;
        RECT 73.730000 70.035000 75.000000 70.060000 ;
        RECT 73.730000 90.435000 75.000000 90.630000 ;
        RECT 73.730000 94.770000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 24.370000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  68.935000 24.770000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000   0.000000 73.330000  19.385000 ;
      RECT  1.670000   0.000000 73.330000  19.385000 ;
      RECT  1.670000  24.835000 73.330000  63.685000 ;
      RECT  1.670000  24.835000 73.330000  63.685000 ;
      RECT  1.670000  24.835000 73.330000  63.685000 ;
      RECT  1.670000  24.835000 73.330000  63.685000 ;
      RECT  1.670000  24.835000 73.330000  63.685000 ;
      RECT  1.670000  24.835000 73.330000  63.685000 ;
      RECT  1.670000  24.835000 73.330000  63.685000 ;
      RECT  1.670000  69.635000 24.770000  69.660000 ;
      RECT  1.670000  95.170000 73.330000  95.400000 ;
      RECT  1.670000  95.170000 73.330000 200.000000 ;
      RECT  1.670000  95.170000 73.330000 200.000000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT 20.140000  90.835000 54.920000  95.170000 ;
      RECT 20.140000  90.835000 54.920000 200.000000 ;
      RECT 24.770000   0.000000 50.015000  68.935000 ;
      RECT 24.770000   0.000000 50.015000  69.660000 ;
      RECT 24.770000  19.385000 50.015000  24.835000 ;
      RECT 24.770000  63.685000 50.015000  68.935000 ;
      RECT 24.770000  68.935000 50.260000  69.660000 ;
      RECT 24.800000  68.935000 50.260000 200.000000 ;
      RECT 24.800000  69.660000 50.260000  90.835000 ;
      RECT 50.260000  68.935000 75.000000  69.635000 ;
      RECT 50.260000  69.635000 73.330000  69.660000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT 0.000000   0.000000 75.000000   1.335000 ;
      RECT 0.000000  95.785000 75.000000 174.985000 ;
      RECT 1.765000  14.235000 73.235000  19.085000 ;
      RECT 2.070000   1.335000 72.930000  14.235000 ;
      RECT 2.070000  19.085000 72.930000  95.785000 ;
      RECT 2.070000 174.985000 72.930000 200.000000 ;
  END
END sky130_fd_io__overlay_vddio_hvc


MACRO sky130_fd_io__overlay_vdda_lvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.600000 12.940000 24.500000 16.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 12.940000 74.655000 16.380000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 24.475000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.690000 13.020000  0.890000 13.220000 ;
        RECT  0.690000 13.460000  0.890000 13.660000 ;
        RECT  0.690000 13.900000  0.890000 14.100000 ;
        RECT  0.690000 14.340000  0.890000 14.540000 ;
        RECT  0.690000 14.780000  0.890000 14.980000 ;
        RECT  0.690000 15.220000  0.890000 15.420000 ;
        RECT  0.690000 15.660000  0.890000 15.860000 ;
        RECT  0.690000 16.100000  0.890000 16.300000 ;
        RECT  1.100000 13.020000  1.300000 13.220000 ;
        RECT  1.100000 13.460000  1.300000 13.660000 ;
        RECT  1.100000 13.900000  1.300000 14.100000 ;
        RECT  1.100000 14.340000  1.300000 14.540000 ;
        RECT  1.100000 14.780000  1.300000 14.980000 ;
        RECT  1.100000 15.220000  1.300000 15.420000 ;
        RECT  1.100000 15.660000  1.300000 15.860000 ;
        RECT  1.100000 16.100000  1.300000 16.300000 ;
        RECT  1.510000 13.020000  1.710000 13.220000 ;
        RECT  1.510000 13.460000  1.710000 13.660000 ;
        RECT  1.510000 13.900000  1.710000 14.100000 ;
        RECT  1.510000 14.340000  1.710000 14.540000 ;
        RECT  1.510000 14.780000  1.710000 14.980000 ;
        RECT  1.510000 15.220000  1.710000 15.420000 ;
        RECT  1.510000 15.660000  1.710000 15.860000 ;
        RECT  1.510000 16.100000  1.710000 16.300000 ;
        RECT  1.920000 13.020000  2.120000 13.220000 ;
        RECT  1.920000 13.460000  2.120000 13.660000 ;
        RECT  1.920000 13.900000  2.120000 14.100000 ;
        RECT  1.920000 14.340000  2.120000 14.540000 ;
        RECT  1.920000 14.780000  2.120000 14.980000 ;
        RECT  1.920000 15.220000  2.120000 15.420000 ;
        RECT  1.920000 15.660000  2.120000 15.860000 ;
        RECT  1.920000 16.100000  2.120000 16.300000 ;
        RECT  2.330000 13.020000  2.530000 13.220000 ;
        RECT  2.330000 13.460000  2.530000 13.660000 ;
        RECT  2.330000 13.900000  2.530000 14.100000 ;
        RECT  2.330000 14.340000  2.530000 14.540000 ;
        RECT  2.330000 14.780000  2.530000 14.980000 ;
        RECT  2.330000 15.220000  2.530000 15.420000 ;
        RECT  2.330000 15.660000  2.530000 15.860000 ;
        RECT  2.330000 16.100000  2.530000 16.300000 ;
        RECT  2.740000 13.020000  2.940000 13.220000 ;
        RECT  2.740000 13.460000  2.940000 13.660000 ;
        RECT  2.740000 13.900000  2.940000 14.100000 ;
        RECT  2.740000 14.340000  2.940000 14.540000 ;
        RECT  2.740000 14.780000  2.940000 14.980000 ;
        RECT  2.740000 15.220000  2.940000 15.420000 ;
        RECT  2.740000 15.660000  2.940000 15.860000 ;
        RECT  2.740000 16.100000  2.940000 16.300000 ;
        RECT  3.150000 13.020000  3.350000 13.220000 ;
        RECT  3.150000 13.460000  3.350000 13.660000 ;
        RECT  3.150000 13.900000  3.350000 14.100000 ;
        RECT  3.150000 14.340000  3.350000 14.540000 ;
        RECT  3.150000 14.780000  3.350000 14.980000 ;
        RECT  3.150000 15.220000  3.350000 15.420000 ;
        RECT  3.150000 15.660000  3.350000 15.860000 ;
        RECT  3.150000 16.100000  3.350000 16.300000 ;
        RECT  3.555000 13.020000  3.755000 13.220000 ;
        RECT  3.555000 13.460000  3.755000 13.660000 ;
        RECT  3.555000 13.900000  3.755000 14.100000 ;
        RECT  3.555000 14.340000  3.755000 14.540000 ;
        RECT  3.555000 14.780000  3.755000 14.980000 ;
        RECT  3.555000 15.220000  3.755000 15.420000 ;
        RECT  3.555000 15.660000  3.755000 15.860000 ;
        RECT  3.555000 16.100000  3.755000 16.300000 ;
        RECT  3.960000 13.020000  4.160000 13.220000 ;
        RECT  3.960000 13.460000  4.160000 13.660000 ;
        RECT  3.960000 13.900000  4.160000 14.100000 ;
        RECT  3.960000 14.340000  4.160000 14.540000 ;
        RECT  3.960000 14.780000  4.160000 14.980000 ;
        RECT  3.960000 15.220000  4.160000 15.420000 ;
        RECT  3.960000 15.660000  4.160000 15.860000 ;
        RECT  3.960000 16.100000  4.160000 16.300000 ;
        RECT  4.365000 13.020000  4.565000 13.220000 ;
        RECT  4.365000 13.460000  4.565000 13.660000 ;
        RECT  4.365000 13.900000  4.565000 14.100000 ;
        RECT  4.365000 14.340000  4.565000 14.540000 ;
        RECT  4.365000 14.780000  4.565000 14.980000 ;
        RECT  4.365000 15.220000  4.565000 15.420000 ;
        RECT  4.365000 15.660000  4.565000 15.860000 ;
        RECT  4.365000 16.100000  4.565000 16.300000 ;
        RECT  4.770000 13.020000  4.970000 13.220000 ;
        RECT  4.770000 13.460000  4.970000 13.660000 ;
        RECT  4.770000 13.900000  4.970000 14.100000 ;
        RECT  4.770000 14.340000  4.970000 14.540000 ;
        RECT  4.770000 14.780000  4.970000 14.980000 ;
        RECT  4.770000 15.220000  4.970000 15.420000 ;
        RECT  4.770000 15.660000  4.970000 15.860000 ;
        RECT  4.770000 16.100000  4.970000 16.300000 ;
        RECT  5.175000 13.020000  5.375000 13.220000 ;
        RECT  5.175000 13.460000  5.375000 13.660000 ;
        RECT  5.175000 13.900000  5.375000 14.100000 ;
        RECT  5.175000 14.340000  5.375000 14.540000 ;
        RECT  5.175000 14.780000  5.375000 14.980000 ;
        RECT  5.175000 15.220000  5.375000 15.420000 ;
        RECT  5.175000 15.660000  5.375000 15.860000 ;
        RECT  5.175000 16.100000  5.375000 16.300000 ;
        RECT  5.580000 13.020000  5.780000 13.220000 ;
        RECT  5.580000 13.460000  5.780000 13.660000 ;
        RECT  5.580000 13.900000  5.780000 14.100000 ;
        RECT  5.580000 14.340000  5.780000 14.540000 ;
        RECT  5.580000 14.780000  5.780000 14.980000 ;
        RECT  5.580000 15.220000  5.780000 15.420000 ;
        RECT  5.580000 15.660000  5.780000 15.860000 ;
        RECT  5.580000 16.100000  5.780000 16.300000 ;
        RECT  5.985000 13.020000  6.185000 13.220000 ;
        RECT  5.985000 13.460000  6.185000 13.660000 ;
        RECT  5.985000 13.900000  6.185000 14.100000 ;
        RECT  5.985000 14.340000  6.185000 14.540000 ;
        RECT  5.985000 14.780000  6.185000 14.980000 ;
        RECT  5.985000 15.220000  6.185000 15.420000 ;
        RECT  5.985000 15.660000  6.185000 15.860000 ;
        RECT  5.985000 16.100000  6.185000 16.300000 ;
        RECT  6.390000 13.020000  6.590000 13.220000 ;
        RECT  6.390000 13.460000  6.590000 13.660000 ;
        RECT  6.390000 13.900000  6.590000 14.100000 ;
        RECT  6.390000 14.340000  6.590000 14.540000 ;
        RECT  6.390000 14.780000  6.590000 14.980000 ;
        RECT  6.390000 15.220000  6.590000 15.420000 ;
        RECT  6.390000 15.660000  6.590000 15.860000 ;
        RECT  6.390000 16.100000  6.590000 16.300000 ;
        RECT  6.795000 13.020000  6.995000 13.220000 ;
        RECT  6.795000 13.460000  6.995000 13.660000 ;
        RECT  6.795000 13.900000  6.995000 14.100000 ;
        RECT  6.795000 14.340000  6.995000 14.540000 ;
        RECT  6.795000 14.780000  6.995000 14.980000 ;
        RECT  6.795000 15.220000  6.995000 15.420000 ;
        RECT  6.795000 15.660000  6.995000 15.860000 ;
        RECT  6.795000 16.100000  6.995000 16.300000 ;
        RECT  7.200000 13.020000  7.400000 13.220000 ;
        RECT  7.200000 13.460000  7.400000 13.660000 ;
        RECT  7.200000 13.900000  7.400000 14.100000 ;
        RECT  7.200000 14.340000  7.400000 14.540000 ;
        RECT  7.200000 14.780000  7.400000 14.980000 ;
        RECT  7.200000 15.220000  7.400000 15.420000 ;
        RECT  7.200000 15.660000  7.400000 15.860000 ;
        RECT  7.200000 16.100000  7.400000 16.300000 ;
        RECT  7.605000 13.020000  7.805000 13.220000 ;
        RECT  7.605000 13.460000  7.805000 13.660000 ;
        RECT  7.605000 13.900000  7.805000 14.100000 ;
        RECT  7.605000 14.340000  7.805000 14.540000 ;
        RECT  7.605000 14.780000  7.805000 14.980000 ;
        RECT  7.605000 15.220000  7.805000 15.420000 ;
        RECT  7.605000 15.660000  7.805000 15.860000 ;
        RECT  7.605000 16.100000  7.805000 16.300000 ;
        RECT  8.010000 13.020000  8.210000 13.220000 ;
        RECT  8.010000 13.460000  8.210000 13.660000 ;
        RECT  8.010000 13.900000  8.210000 14.100000 ;
        RECT  8.010000 14.340000  8.210000 14.540000 ;
        RECT  8.010000 14.780000  8.210000 14.980000 ;
        RECT  8.010000 15.220000  8.210000 15.420000 ;
        RECT  8.010000 15.660000  8.210000 15.860000 ;
        RECT  8.010000 16.100000  8.210000 16.300000 ;
        RECT  8.415000 13.020000  8.615000 13.220000 ;
        RECT  8.415000 13.460000  8.615000 13.660000 ;
        RECT  8.415000 13.900000  8.615000 14.100000 ;
        RECT  8.415000 14.340000  8.615000 14.540000 ;
        RECT  8.415000 14.780000  8.615000 14.980000 ;
        RECT  8.415000 15.220000  8.615000 15.420000 ;
        RECT  8.415000 15.660000  8.615000 15.860000 ;
        RECT  8.415000 16.100000  8.615000 16.300000 ;
        RECT  8.820000 13.020000  9.020000 13.220000 ;
        RECT  8.820000 13.460000  9.020000 13.660000 ;
        RECT  8.820000 13.900000  9.020000 14.100000 ;
        RECT  8.820000 14.340000  9.020000 14.540000 ;
        RECT  8.820000 14.780000  9.020000 14.980000 ;
        RECT  8.820000 15.220000  9.020000 15.420000 ;
        RECT  8.820000 15.660000  9.020000 15.860000 ;
        RECT  8.820000 16.100000  9.020000 16.300000 ;
        RECT  9.225000 13.020000  9.425000 13.220000 ;
        RECT  9.225000 13.460000  9.425000 13.660000 ;
        RECT  9.225000 13.900000  9.425000 14.100000 ;
        RECT  9.225000 14.340000  9.425000 14.540000 ;
        RECT  9.225000 14.780000  9.425000 14.980000 ;
        RECT  9.225000 15.220000  9.425000 15.420000 ;
        RECT  9.225000 15.660000  9.425000 15.860000 ;
        RECT  9.225000 16.100000  9.425000 16.300000 ;
        RECT  9.630000 13.020000  9.830000 13.220000 ;
        RECT  9.630000 13.460000  9.830000 13.660000 ;
        RECT  9.630000 13.900000  9.830000 14.100000 ;
        RECT  9.630000 14.340000  9.830000 14.540000 ;
        RECT  9.630000 14.780000  9.830000 14.980000 ;
        RECT  9.630000 15.220000  9.830000 15.420000 ;
        RECT  9.630000 15.660000  9.830000 15.860000 ;
        RECT  9.630000 16.100000  9.830000 16.300000 ;
        RECT 10.035000 13.020000 10.235000 13.220000 ;
        RECT 10.035000 13.460000 10.235000 13.660000 ;
        RECT 10.035000 13.900000 10.235000 14.100000 ;
        RECT 10.035000 14.340000 10.235000 14.540000 ;
        RECT 10.035000 14.780000 10.235000 14.980000 ;
        RECT 10.035000 15.220000 10.235000 15.420000 ;
        RECT 10.035000 15.660000 10.235000 15.860000 ;
        RECT 10.035000 16.100000 10.235000 16.300000 ;
        RECT 10.440000 13.020000 10.640000 13.220000 ;
        RECT 10.440000 13.460000 10.640000 13.660000 ;
        RECT 10.440000 13.900000 10.640000 14.100000 ;
        RECT 10.440000 14.340000 10.640000 14.540000 ;
        RECT 10.440000 14.780000 10.640000 14.980000 ;
        RECT 10.440000 15.220000 10.640000 15.420000 ;
        RECT 10.440000 15.660000 10.640000 15.860000 ;
        RECT 10.440000 16.100000 10.640000 16.300000 ;
        RECT 10.845000 13.020000 11.045000 13.220000 ;
        RECT 10.845000 13.460000 11.045000 13.660000 ;
        RECT 10.845000 13.900000 11.045000 14.100000 ;
        RECT 10.845000 14.340000 11.045000 14.540000 ;
        RECT 10.845000 14.780000 11.045000 14.980000 ;
        RECT 10.845000 15.220000 11.045000 15.420000 ;
        RECT 10.845000 15.660000 11.045000 15.860000 ;
        RECT 10.845000 16.100000 11.045000 16.300000 ;
        RECT 11.250000 13.020000 11.450000 13.220000 ;
        RECT 11.250000 13.460000 11.450000 13.660000 ;
        RECT 11.250000 13.900000 11.450000 14.100000 ;
        RECT 11.250000 14.340000 11.450000 14.540000 ;
        RECT 11.250000 14.780000 11.450000 14.980000 ;
        RECT 11.250000 15.220000 11.450000 15.420000 ;
        RECT 11.250000 15.660000 11.450000 15.860000 ;
        RECT 11.250000 16.100000 11.450000 16.300000 ;
        RECT 11.655000 13.020000 11.855000 13.220000 ;
        RECT 11.655000 13.460000 11.855000 13.660000 ;
        RECT 11.655000 13.900000 11.855000 14.100000 ;
        RECT 11.655000 14.340000 11.855000 14.540000 ;
        RECT 11.655000 14.780000 11.855000 14.980000 ;
        RECT 11.655000 15.220000 11.855000 15.420000 ;
        RECT 11.655000 15.660000 11.855000 15.860000 ;
        RECT 11.655000 16.100000 11.855000 16.300000 ;
        RECT 12.060000 13.020000 12.260000 13.220000 ;
        RECT 12.060000 13.460000 12.260000 13.660000 ;
        RECT 12.060000 13.900000 12.260000 14.100000 ;
        RECT 12.060000 14.340000 12.260000 14.540000 ;
        RECT 12.060000 14.780000 12.260000 14.980000 ;
        RECT 12.060000 15.220000 12.260000 15.420000 ;
        RECT 12.060000 15.660000 12.260000 15.860000 ;
        RECT 12.060000 16.100000 12.260000 16.300000 ;
        RECT 12.465000 13.020000 12.665000 13.220000 ;
        RECT 12.465000 13.460000 12.665000 13.660000 ;
        RECT 12.465000 13.900000 12.665000 14.100000 ;
        RECT 12.465000 14.340000 12.665000 14.540000 ;
        RECT 12.465000 14.780000 12.665000 14.980000 ;
        RECT 12.465000 15.220000 12.665000 15.420000 ;
        RECT 12.465000 15.660000 12.665000 15.860000 ;
        RECT 12.465000 16.100000 12.665000 16.300000 ;
        RECT 12.870000 13.020000 13.070000 13.220000 ;
        RECT 12.870000 13.460000 13.070000 13.660000 ;
        RECT 12.870000 13.900000 13.070000 14.100000 ;
        RECT 12.870000 14.340000 13.070000 14.540000 ;
        RECT 12.870000 14.780000 13.070000 14.980000 ;
        RECT 12.870000 15.220000 13.070000 15.420000 ;
        RECT 12.870000 15.660000 13.070000 15.860000 ;
        RECT 12.870000 16.100000 13.070000 16.300000 ;
        RECT 13.275000 13.020000 13.475000 13.220000 ;
        RECT 13.275000 13.460000 13.475000 13.660000 ;
        RECT 13.275000 13.900000 13.475000 14.100000 ;
        RECT 13.275000 14.340000 13.475000 14.540000 ;
        RECT 13.275000 14.780000 13.475000 14.980000 ;
        RECT 13.275000 15.220000 13.475000 15.420000 ;
        RECT 13.275000 15.660000 13.475000 15.860000 ;
        RECT 13.275000 16.100000 13.475000 16.300000 ;
        RECT 13.680000 13.020000 13.880000 13.220000 ;
        RECT 13.680000 13.460000 13.880000 13.660000 ;
        RECT 13.680000 13.900000 13.880000 14.100000 ;
        RECT 13.680000 14.340000 13.880000 14.540000 ;
        RECT 13.680000 14.780000 13.880000 14.980000 ;
        RECT 13.680000 15.220000 13.880000 15.420000 ;
        RECT 13.680000 15.660000 13.880000 15.860000 ;
        RECT 13.680000 16.100000 13.880000 16.300000 ;
        RECT 14.085000 13.020000 14.285000 13.220000 ;
        RECT 14.085000 13.460000 14.285000 13.660000 ;
        RECT 14.085000 13.900000 14.285000 14.100000 ;
        RECT 14.085000 14.340000 14.285000 14.540000 ;
        RECT 14.085000 14.780000 14.285000 14.980000 ;
        RECT 14.085000 15.220000 14.285000 15.420000 ;
        RECT 14.085000 15.660000 14.285000 15.860000 ;
        RECT 14.085000 16.100000 14.285000 16.300000 ;
        RECT 14.490000 13.020000 14.690000 13.220000 ;
        RECT 14.490000 13.460000 14.690000 13.660000 ;
        RECT 14.490000 13.900000 14.690000 14.100000 ;
        RECT 14.490000 14.340000 14.690000 14.540000 ;
        RECT 14.490000 14.780000 14.690000 14.980000 ;
        RECT 14.490000 15.220000 14.690000 15.420000 ;
        RECT 14.490000 15.660000 14.690000 15.860000 ;
        RECT 14.490000 16.100000 14.690000 16.300000 ;
        RECT 14.895000 13.020000 15.095000 13.220000 ;
        RECT 14.895000 13.460000 15.095000 13.660000 ;
        RECT 14.895000 13.900000 15.095000 14.100000 ;
        RECT 14.895000 14.340000 15.095000 14.540000 ;
        RECT 14.895000 14.780000 15.095000 14.980000 ;
        RECT 14.895000 15.220000 15.095000 15.420000 ;
        RECT 14.895000 15.660000 15.095000 15.860000 ;
        RECT 14.895000 16.100000 15.095000 16.300000 ;
        RECT 15.300000 13.020000 15.500000 13.220000 ;
        RECT 15.300000 13.460000 15.500000 13.660000 ;
        RECT 15.300000 13.900000 15.500000 14.100000 ;
        RECT 15.300000 14.340000 15.500000 14.540000 ;
        RECT 15.300000 14.780000 15.500000 14.980000 ;
        RECT 15.300000 15.220000 15.500000 15.420000 ;
        RECT 15.300000 15.660000 15.500000 15.860000 ;
        RECT 15.300000 16.100000 15.500000 16.300000 ;
        RECT 15.705000 13.020000 15.905000 13.220000 ;
        RECT 15.705000 13.460000 15.905000 13.660000 ;
        RECT 15.705000 13.900000 15.905000 14.100000 ;
        RECT 15.705000 14.340000 15.905000 14.540000 ;
        RECT 15.705000 14.780000 15.905000 14.980000 ;
        RECT 15.705000 15.220000 15.905000 15.420000 ;
        RECT 15.705000 15.660000 15.905000 15.860000 ;
        RECT 15.705000 16.100000 15.905000 16.300000 ;
        RECT 16.110000 13.020000 16.310000 13.220000 ;
        RECT 16.110000 13.460000 16.310000 13.660000 ;
        RECT 16.110000 13.900000 16.310000 14.100000 ;
        RECT 16.110000 14.340000 16.310000 14.540000 ;
        RECT 16.110000 14.780000 16.310000 14.980000 ;
        RECT 16.110000 15.220000 16.310000 15.420000 ;
        RECT 16.110000 15.660000 16.310000 15.860000 ;
        RECT 16.110000 16.100000 16.310000 16.300000 ;
        RECT 16.515000 13.020000 16.715000 13.220000 ;
        RECT 16.515000 13.460000 16.715000 13.660000 ;
        RECT 16.515000 13.900000 16.715000 14.100000 ;
        RECT 16.515000 14.340000 16.715000 14.540000 ;
        RECT 16.515000 14.780000 16.715000 14.980000 ;
        RECT 16.515000 15.220000 16.715000 15.420000 ;
        RECT 16.515000 15.660000 16.715000 15.860000 ;
        RECT 16.515000 16.100000 16.715000 16.300000 ;
        RECT 16.920000 13.020000 17.120000 13.220000 ;
        RECT 16.920000 13.460000 17.120000 13.660000 ;
        RECT 16.920000 13.900000 17.120000 14.100000 ;
        RECT 16.920000 14.340000 17.120000 14.540000 ;
        RECT 16.920000 14.780000 17.120000 14.980000 ;
        RECT 16.920000 15.220000 17.120000 15.420000 ;
        RECT 16.920000 15.660000 17.120000 15.860000 ;
        RECT 16.920000 16.100000 17.120000 16.300000 ;
        RECT 17.325000 13.020000 17.525000 13.220000 ;
        RECT 17.325000 13.460000 17.525000 13.660000 ;
        RECT 17.325000 13.900000 17.525000 14.100000 ;
        RECT 17.325000 14.340000 17.525000 14.540000 ;
        RECT 17.325000 14.780000 17.525000 14.980000 ;
        RECT 17.325000 15.220000 17.525000 15.420000 ;
        RECT 17.325000 15.660000 17.525000 15.860000 ;
        RECT 17.325000 16.100000 17.525000 16.300000 ;
        RECT 17.730000 13.020000 17.930000 13.220000 ;
        RECT 17.730000 13.460000 17.930000 13.660000 ;
        RECT 17.730000 13.900000 17.930000 14.100000 ;
        RECT 17.730000 14.340000 17.930000 14.540000 ;
        RECT 17.730000 14.780000 17.930000 14.980000 ;
        RECT 17.730000 15.220000 17.930000 15.420000 ;
        RECT 17.730000 15.660000 17.930000 15.860000 ;
        RECT 17.730000 16.100000 17.930000 16.300000 ;
        RECT 18.135000 13.020000 18.335000 13.220000 ;
        RECT 18.135000 13.460000 18.335000 13.660000 ;
        RECT 18.135000 13.900000 18.335000 14.100000 ;
        RECT 18.135000 14.340000 18.335000 14.540000 ;
        RECT 18.135000 14.780000 18.335000 14.980000 ;
        RECT 18.135000 15.220000 18.335000 15.420000 ;
        RECT 18.135000 15.660000 18.335000 15.860000 ;
        RECT 18.135000 16.100000 18.335000 16.300000 ;
        RECT 18.540000 13.020000 18.740000 13.220000 ;
        RECT 18.540000 13.460000 18.740000 13.660000 ;
        RECT 18.540000 13.900000 18.740000 14.100000 ;
        RECT 18.540000 14.340000 18.740000 14.540000 ;
        RECT 18.540000 14.780000 18.740000 14.980000 ;
        RECT 18.540000 15.220000 18.740000 15.420000 ;
        RECT 18.540000 15.660000 18.740000 15.860000 ;
        RECT 18.540000 16.100000 18.740000 16.300000 ;
        RECT 18.945000 13.020000 19.145000 13.220000 ;
        RECT 18.945000 13.460000 19.145000 13.660000 ;
        RECT 18.945000 13.900000 19.145000 14.100000 ;
        RECT 18.945000 14.340000 19.145000 14.540000 ;
        RECT 18.945000 14.780000 19.145000 14.980000 ;
        RECT 18.945000 15.220000 19.145000 15.420000 ;
        RECT 18.945000 15.660000 19.145000 15.860000 ;
        RECT 18.945000 16.100000 19.145000 16.300000 ;
        RECT 19.350000 13.020000 19.550000 13.220000 ;
        RECT 19.350000 13.460000 19.550000 13.660000 ;
        RECT 19.350000 13.900000 19.550000 14.100000 ;
        RECT 19.350000 14.340000 19.550000 14.540000 ;
        RECT 19.350000 14.780000 19.550000 14.980000 ;
        RECT 19.350000 15.220000 19.550000 15.420000 ;
        RECT 19.350000 15.660000 19.550000 15.860000 ;
        RECT 19.350000 16.100000 19.550000 16.300000 ;
        RECT 19.755000 13.020000 19.955000 13.220000 ;
        RECT 19.755000 13.460000 19.955000 13.660000 ;
        RECT 19.755000 13.900000 19.955000 14.100000 ;
        RECT 19.755000 14.340000 19.955000 14.540000 ;
        RECT 19.755000 14.780000 19.955000 14.980000 ;
        RECT 19.755000 15.220000 19.955000 15.420000 ;
        RECT 19.755000 15.660000 19.955000 15.860000 ;
        RECT 19.755000 16.100000 19.955000 16.300000 ;
        RECT 20.160000 13.020000 20.360000 13.220000 ;
        RECT 20.160000 13.460000 20.360000 13.660000 ;
        RECT 20.160000 13.900000 20.360000 14.100000 ;
        RECT 20.160000 14.340000 20.360000 14.540000 ;
        RECT 20.160000 14.780000 20.360000 14.980000 ;
        RECT 20.160000 15.220000 20.360000 15.420000 ;
        RECT 20.160000 15.660000 20.360000 15.860000 ;
        RECT 20.160000 16.100000 20.360000 16.300000 ;
        RECT 20.565000 13.020000 20.765000 13.220000 ;
        RECT 20.565000 13.460000 20.765000 13.660000 ;
        RECT 20.565000 13.900000 20.765000 14.100000 ;
        RECT 20.565000 14.340000 20.765000 14.540000 ;
        RECT 20.565000 14.780000 20.765000 14.980000 ;
        RECT 20.565000 15.220000 20.765000 15.420000 ;
        RECT 20.565000 15.660000 20.765000 15.860000 ;
        RECT 20.565000 16.100000 20.765000 16.300000 ;
        RECT 20.970000 13.020000 21.170000 13.220000 ;
        RECT 20.970000 13.460000 21.170000 13.660000 ;
        RECT 20.970000 13.900000 21.170000 14.100000 ;
        RECT 20.970000 14.340000 21.170000 14.540000 ;
        RECT 20.970000 14.780000 21.170000 14.980000 ;
        RECT 20.970000 15.220000 21.170000 15.420000 ;
        RECT 20.970000 15.660000 21.170000 15.860000 ;
        RECT 20.970000 16.100000 21.170000 16.300000 ;
        RECT 21.375000 13.020000 21.575000 13.220000 ;
        RECT 21.375000 13.460000 21.575000 13.660000 ;
        RECT 21.375000 13.900000 21.575000 14.100000 ;
        RECT 21.375000 14.340000 21.575000 14.540000 ;
        RECT 21.375000 14.780000 21.575000 14.980000 ;
        RECT 21.375000 15.220000 21.575000 15.420000 ;
        RECT 21.375000 15.660000 21.575000 15.860000 ;
        RECT 21.375000 16.100000 21.575000 16.300000 ;
        RECT 21.780000 13.020000 21.980000 13.220000 ;
        RECT 21.780000 13.460000 21.980000 13.660000 ;
        RECT 21.780000 13.900000 21.980000 14.100000 ;
        RECT 21.780000 14.340000 21.980000 14.540000 ;
        RECT 21.780000 14.780000 21.980000 14.980000 ;
        RECT 21.780000 15.220000 21.980000 15.420000 ;
        RECT 21.780000 15.660000 21.980000 15.860000 ;
        RECT 21.780000 16.100000 21.980000 16.300000 ;
        RECT 22.185000 13.020000 22.385000 13.220000 ;
        RECT 22.185000 13.460000 22.385000 13.660000 ;
        RECT 22.185000 13.900000 22.385000 14.100000 ;
        RECT 22.185000 14.340000 22.385000 14.540000 ;
        RECT 22.185000 14.780000 22.385000 14.980000 ;
        RECT 22.185000 15.220000 22.385000 15.420000 ;
        RECT 22.185000 15.660000 22.385000 15.860000 ;
        RECT 22.185000 16.100000 22.385000 16.300000 ;
        RECT 22.590000 13.020000 22.790000 13.220000 ;
        RECT 22.590000 13.460000 22.790000 13.660000 ;
        RECT 22.590000 13.900000 22.790000 14.100000 ;
        RECT 22.590000 14.340000 22.790000 14.540000 ;
        RECT 22.590000 14.780000 22.790000 14.980000 ;
        RECT 22.590000 15.220000 22.790000 15.420000 ;
        RECT 22.590000 15.660000 22.790000 15.860000 ;
        RECT 22.590000 16.100000 22.790000 16.300000 ;
        RECT 22.995000 13.020000 23.195000 13.220000 ;
        RECT 22.995000 13.460000 23.195000 13.660000 ;
        RECT 22.995000 13.900000 23.195000 14.100000 ;
        RECT 22.995000 14.340000 23.195000 14.540000 ;
        RECT 22.995000 14.780000 23.195000 14.980000 ;
        RECT 22.995000 15.220000 23.195000 15.420000 ;
        RECT 22.995000 15.660000 23.195000 15.860000 ;
        RECT 22.995000 16.100000 23.195000 16.300000 ;
        RECT 23.400000 13.020000 23.600000 13.220000 ;
        RECT 23.400000 13.460000 23.600000 13.660000 ;
        RECT 23.400000 13.900000 23.600000 14.100000 ;
        RECT 23.400000 14.340000 23.600000 14.540000 ;
        RECT 23.400000 14.780000 23.600000 14.980000 ;
        RECT 23.400000 15.220000 23.600000 15.420000 ;
        RECT 23.400000 15.660000 23.600000 15.860000 ;
        RECT 23.400000 16.100000 23.600000 16.300000 ;
        RECT 23.805000 13.020000 24.005000 13.220000 ;
        RECT 23.805000 13.460000 24.005000 13.660000 ;
        RECT 23.805000 13.900000 24.005000 14.100000 ;
        RECT 23.805000 14.340000 24.005000 14.540000 ;
        RECT 23.805000 14.780000 24.005000 14.980000 ;
        RECT 23.805000 15.220000 24.005000 15.420000 ;
        RECT 23.805000 15.660000 24.005000 15.860000 ;
        RECT 23.805000 16.100000 24.005000 16.300000 ;
        RECT 24.210000 13.020000 24.410000 13.220000 ;
        RECT 24.210000 13.460000 24.410000 13.660000 ;
        RECT 24.210000 13.900000 24.410000 14.100000 ;
        RECT 24.210000 14.340000 24.410000 14.540000 ;
        RECT 24.210000 14.780000 24.410000 14.980000 ;
        RECT 24.210000 15.220000 24.410000 15.420000 ;
        RECT 24.210000 15.660000 24.410000 15.860000 ;
        RECT 24.210000 16.100000 24.410000 16.300000 ;
        RECT 50.845000 13.020000 51.045000 13.220000 ;
        RECT 50.845000 13.460000 51.045000 13.660000 ;
        RECT 50.845000 13.900000 51.045000 14.100000 ;
        RECT 50.845000 14.340000 51.045000 14.540000 ;
        RECT 50.845000 14.780000 51.045000 14.980000 ;
        RECT 50.845000 15.220000 51.045000 15.420000 ;
        RECT 50.845000 15.660000 51.045000 15.860000 ;
        RECT 50.845000 16.100000 51.045000 16.300000 ;
        RECT 51.255000 13.020000 51.455000 13.220000 ;
        RECT 51.255000 13.460000 51.455000 13.660000 ;
        RECT 51.255000 13.900000 51.455000 14.100000 ;
        RECT 51.255000 14.340000 51.455000 14.540000 ;
        RECT 51.255000 14.780000 51.455000 14.980000 ;
        RECT 51.255000 15.220000 51.455000 15.420000 ;
        RECT 51.255000 15.660000 51.455000 15.860000 ;
        RECT 51.255000 16.100000 51.455000 16.300000 ;
        RECT 51.665000 13.020000 51.865000 13.220000 ;
        RECT 51.665000 13.460000 51.865000 13.660000 ;
        RECT 51.665000 13.900000 51.865000 14.100000 ;
        RECT 51.665000 14.340000 51.865000 14.540000 ;
        RECT 51.665000 14.780000 51.865000 14.980000 ;
        RECT 51.665000 15.220000 51.865000 15.420000 ;
        RECT 51.665000 15.660000 51.865000 15.860000 ;
        RECT 51.665000 16.100000 51.865000 16.300000 ;
        RECT 52.075000 13.020000 52.275000 13.220000 ;
        RECT 52.075000 13.460000 52.275000 13.660000 ;
        RECT 52.075000 13.900000 52.275000 14.100000 ;
        RECT 52.075000 14.340000 52.275000 14.540000 ;
        RECT 52.075000 14.780000 52.275000 14.980000 ;
        RECT 52.075000 15.220000 52.275000 15.420000 ;
        RECT 52.075000 15.660000 52.275000 15.860000 ;
        RECT 52.075000 16.100000 52.275000 16.300000 ;
        RECT 52.485000 13.020000 52.685000 13.220000 ;
        RECT 52.485000 13.460000 52.685000 13.660000 ;
        RECT 52.485000 13.900000 52.685000 14.100000 ;
        RECT 52.485000 14.340000 52.685000 14.540000 ;
        RECT 52.485000 14.780000 52.685000 14.980000 ;
        RECT 52.485000 15.220000 52.685000 15.420000 ;
        RECT 52.485000 15.660000 52.685000 15.860000 ;
        RECT 52.485000 16.100000 52.685000 16.300000 ;
        RECT 52.895000 13.020000 53.095000 13.220000 ;
        RECT 52.895000 13.460000 53.095000 13.660000 ;
        RECT 52.895000 13.900000 53.095000 14.100000 ;
        RECT 52.895000 14.340000 53.095000 14.540000 ;
        RECT 52.895000 14.780000 53.095000 14.980000 ;
        RECT 52.895000 15.220000 53.095000 15.420000 ;
        RECT 52.895000 15.660000 53.095000 15.860000 ;
        RECT 52.895000 16.100000 53.095000 16.300000 ;
        RECT 53.305000 13.020000 53.505000 13.220000 ;
        RECT 53.305000 13.460000 53.505000 13.660000 ;
        RECT 53.305000 13.900000 53.505000 14.100000 ;
        RECT 53.305000 14.340000 53.505000 14.540000 ;
        RECT 53.305000 14.780000 53.505000 14.980000 ;
        RECT 53.305000 15.220000 53.505000 15.420000 ;
        RECT 53.305000 15.660000 53.505000 15.860000 ;
        RECT 53.305000 16.100000 53.505000 16.300000 ;
        RECT 53.710000 13.020000 53.910000 13.220000 ;
        RECT 53.710000 13.460000 53.910000 13.660000 ;
        RECT 53.710000 13.900000 53.910000 14.100000 ;
        RECT 53.710000 14.340000 53.910000 14.540000 ;
        RECT 53.710000 14.780000 53.910000 14.980000 ;
        RECT 53.710000 15.220000 53.910000 15.420000 ;
        RECT 53.710000 15.660000 53.910000 15.860000 ;
        RECT 53.710000 16.100000 53.910000 16.300000 ;
        RECT 54.115000 13.020000 54.315000 13.220000 ;
        RECT 54.115000 13.460000 54.315000 13.660000 ;
        RECT 54.115000 13.900000 54.315000 14.100000 ;
        RECT 54.115000 14.340000 54.315000 14.540000 ;
        RECT 54.115000 14.780000 54.315000 14.980000 ;
        RECT 54.115000 15.220000 54.315000 15.420000 ;
        RECT 54.115000 15.660000 54.315000 15.860000 ;
        RECT 54.115000 16.100000 54.315000 16.300000 ;
        RECT 54.520000 13.020000 54.720000 13.220000 ;
        RECT 54.520000 13.460000 54.720000 13.660000 ;
        RECT 54.520000 13.900000 54.720000 14.100000 ;
        RECT 54.520000 14.340000 54.720000 14.540000 ;
        RECT 54.520000 14.780000 54.720000 14.980000 ;
        RECT 54.520000 15.220000 54.720000 15.420000 ;
        RECT 54.520000 15.660000 54.720000 15.860000 ;
        RECT 54.520000 16.100000 54.720000 16.300000 ;
        RECT 54.925000 13.020000 55.125000 13.220000 ;
        RECT 54.925000 13.460000 55.125000 13.660000 ;
        RECT 54.925000 13.900000 55.125000 14.100000 ;
        RECT 54.925000 14.340000 55.125000 14.540000 ;
        RECT 54.925000 14.780000 55.125000 14.980000 ;
        RECT 54.925000 15.220000 55.125000 15.420000 ;
        RECT 54.925000 15.660000 55.125000 15.860000 ;
        RECT 54.925000 16.100000 55.125000 16.300000 ;
        RECT 55.330000 13.020000 55.530000 13.220000 ;
        RECT 55.330000 13.460000 55.530000 13.660000 ;
        RECT 55.330000 13.900000 55.530000 14.100000 ;
        RECT 55.330000 14.340000 55.530000 14.540000 ;
        RECT 55.330000 14.780000 55.530000 14.980000 ;
        RECT 55.330000 15.220000 55.530000 15.420000 ;
        RECT 55.330000 15.660000 55.530000 15.860000 ;
        RECT 55.330000 16.100000 55.530000 16.300000 ;
        RECT 55.735000 13.020000 55.935000 13.220000 ;
        RECT 55.735000 13.460000 55.935000 13.660000 ;
        RECT 55.735000 13.900000 55.935000 14.100000 ;
        RECT 55.735000 14.340000 55.935000 14.540000 ;
        RECT 55.735000 14.780000 55.935000 14.980000 ;
        RECT 55.735000 15.220000 55.935000 15.420000 ;
        RECT 55.735000 15.660000 55.935000 15.860000 ;
        RECT 55.735000 16.100000 55.935000 16.300000 ;
        RECT 56.140000 13.020000 56.340000 13.220000 ;
        RECT 56.140000 13.460000 56.340000 13.660000 ;
        RECT 56.140000 13.900000 56.340000 14.100000 ;
        RECT 56.140000 14.340000 56.340000 14.540000 ;
        RECT 56.140000 14.780000 56.340000 14.980000 ;
        RECT 56.140000 15.220000 56.340000 15.420000 ;
        RECT 56.140000 15.660000 56.340000 15.860000 ;
        RECT 56.140000 16.100000 56.340000 16.300000 ;
        RECT 56.545000 13.020000 56.745000 13.220000 ;
        RECT 56.545000 13.460000 56.745000 13.660000 ;
        RECT 56.545000 13.900000 56.745000 14.100000 ;
        RECT 56.545000 14.340000 56.745000 14.540000 ;
        RECT 56.545000 14.780000 56.745000 14.980000 ;
        RECT 56.545000 15.220000 56.745000 15.420000 ;
        RECT 56.545000 15.660000 56.745000 15.860000 ;
        RECT 56.545000 16.100000 56.745000 16.300000 ;
        RECT 56.950000 13.020000 57.150000 13.220000 ;
        RECT 56.950000 13.460000 57.150000 13.660000 ;
        RECT 56.950000 13.900000 57.150000 14.100000 ;
        RECT 56.950000 14.340000 57.150000 14.540000 ;
        RECT 56.950000 14.780000 57.150000 14.980000 ;
        RECT 56.950000 15.220000 57.150000 15.420000 ;
        RECT 56.950000 15.660000 57.150000 15.860000 ;
        RECT 56.950000 16.100000 57.150000 16.300000 ;
        RECT 57.355000 13.020000 57.555000 13.220000 ;
        RECT 57.355000 13.460000 57.555000 13.660000 ;
        RECT 57.355000 13.900000 57.555000 14.100000 ;
        RECT 57.355000 14.340000 57.555000 14.540000 ;
        RECT 57.355000 14.780000 57.555000 14.980000 ;
        RECT 57.355000 15.220000 57.555000 15.420000 ;
        RECT 57.355000 15.660000 57.555000 15.860000 ;
        RECT 57.355000 16.100000 57.555000 16.300000 ;
        RECT 57.760000 13.020000 57.960000 13.220000 ;
        RECT 57.760000 13.460000 57.960000 13.660000 ;
        RECT 57.760000 13.900000 57.960000 14.100000 ;
        RECT 57.760000 14.340000 57.960000 14.540000 ;
        RECT 57.760000 14.780000 57.960000 14.980000 ;
        RECT 57.760000 15.220000 57.960000 15.420000 ;
        RECT 57.760000 15.660000 57.960000 15.860000 ;
        RECT 57.760000 16.100000 57.960000 16.300000 ;
        RECT 58.165000 13.020000 58.365000 13.220000 ;
        RECT 58.165000 13.460000 58.365000 13.660000 ;
        RECT 58.165000 13.900000 58.365000 14.100000 ;
        RECT 58.165000 14.340000 58.365000 14.540000 ;
        RECT 58.165000 14.780000 58.365000 14.980000 ;
        RECT 58.165000 15.220000 58.365000 15.420000 ;
        RECT 58.165000 15.660000 58.365000 15.860000 ;
        RECT 58.165000 16.100000 58.365000 16.300000 ;
        RECT 58.570000 13.020000 58.770000 13.220000 ;
        RECT 58.570000 13.460000 58.770000 13.660000 ;
        RECT 58.570000 13.900000 58.770000 14.100000 ;
        RECT 58.570000 14.340000 58.770000 14.540000 ;
        RECT 58.570000 14.780000 58.770000 14.980000 ;
        RECT 58.570000 15.220000 58.770000 15.420000 ;
        RECT 58.570000 15.660000 58.770000 15.860000 ;
        RECT 58.570000 16.100000 58.770000 16.300000 ;
        RECT 58.975000 13.020000 59.175000 13.220000 ;
        RECT 58.975000 13.460000 59.175000 13.660000 ;
        RECT 58.975000 13.900000 59.175000 14.100000 ;
        RECT 58.975000 14.340000 59.175000 14.540000 ;
        RECT 58.975000 14.780000 59.175000 14.980000 ;
        RECT 58.975000 15.220000 59.175000 15.420000 ;
        RECT 58.975000 15.660000 59.175000 15.860000 ;
        RECT 58.975000 16.100000 59.175000 16.300000 ;
        RECT 59.380000 13.020000 59.580000 13.220000 ;
        RECT 59.380000 13.460000 59.580000 13.660000 ;
        RECT 59.380000 13.900000 59.580000 14.100000 ;
        RECT 59.380000 14.340000 59.580000 14.540000 ;
        RECT 59.380000 14.780000 59.580000 14.980000 ;
        RECT 59.380000 15.220000 59.580000 15.420000 ;
        RECT 59.380000 15.660000 59.580000 15.860000 ;
        RECT 59.380000 16.100000 59.580000 16.300000 ;
        RECT 59.785000 13.020000 59.985000 13.220000 ;
        RECT 59.785000 13.460000 59.985000 13.660000 ;
        RECT 59.785000 13.900000 59.985000 14.100000 ;
        RECT 59.785000 14.340000 59.985000 14.540000 ;
        RECT 59.785000 14.780000 59.985000 14.980000 ;
        RECT 59.785000 15.220000 59.985000 15.420000 ;
        RECT 59.785000 15.660000 59.985000 15.860000 ;
        RECT 59.785000 16.100000 59.985000 16.300000 ;
        RECT 60.190000 13.020000 60.390000 13.220000 ;
        RECT 60.190000 13.460000 60.390000 13.660000 ;
        RECT 60.190000 13.900000 60.390000 14.100000 ;
        RECT 60.190000 14.340000 60.390000 14.540000 ;
        RECT 60.190000 14.780000 60.390000 14.980000 ;
        RECT 60.190000 15.220000 60.390000 15.420000 ;
        RECT 60.190000 15.660000 60.390000 15.860000 ;
        RECT 60.190000 16.100000 60.390000 16.300000 ;
        RECT 60.595000 13.020000 60.795000 13.220000 ;
        RECT 60.595000 13.460000 60.795000 13.660000 ;
        RECT 60.595000 13.900000 60.795000 14.100000 ;
        RECT 60.595000 14.340000 60.795000 14.540000 ;
        RECT 60.595000 14.780000 60.795000 14.980000 ;
        RECT 60.595000 15.220000 60.795000 15.420000 ;
        RECT 60.595000 15.660000 60.795000 15.860000 ;
        RECT 60.595000 16.100000 60.795000 16.300000 ;
        RECT 61.000000 13.020000 61.200000 13.220000 ;
        RECT 61.000000 13.460000 61.200000 13.660000 ;
        RECT 61.000000 13.900000 61.200000 14.100000 ;
        RECT 61.000000 14.340000 61.200000 14.540000 ;
        RECT 61.000000 14.780000 61.200000 14.980000 ;
        RECT 61.000000 15.220000 61.200000 15.420000 ;
        RECT 61.000000 15.660000 61.200000 15.860000 ;
        RECT 61.000000 16.100000 61.200000 16.300000 ;
        RECT 61.405000 13.020000 61.605000 13.220000 ;
        RECT 61.405000 13.460000 61.605000 13.660000 ;
        RECT 61.405000 13.900000 61.605000 14.100000 ;
        RECT 61.405000 14.340000 61.605000 14.540000 ;
        RECT 61.405000 14.780000 61.605000 14.980000 ;
        RECT 61.405000 15.220000 61.605000 15.420000 ;
        RECT 61.405000 15.660000 61.605000 15.860000 ;
        RECT 61.405000 16.100000 61.605000 16.300000 ;
        RECT 61.810000 13.020000 62.010000 13.220000 ;
        RECT 61.810000 13.460000 62.010000 13.660000 ;
        RECT 61.810000 13.900000 62.010000 14.100000 ;
        RECT 61.810000 14.340000 62.010000 14.540000 ;
        RECT 61.810000 14.780000 62.010000 14.980000 ;
        RECT 61.810000 15.220000 62.010000 15.420000 ;
        RECT 61.810000 15.660000 62.010000 15.860000 ;
        RECT 61.810000 16.100000 62.010000 16.300000 ;
        RECT 62.215000 13.020000 62.415000 13.220000 ;
        RECT 62.215000 13.460000 62.415000 13.660000 ;
        RECT 62.215000 13.900000 62.415000 14.100000 ;
        RECT 62.215000 14.340000 62.415000 14.540000 ;
        RECT 62.215000 14.780000 62.415000 14.980000 ;
        RECT 62.215000 15.220000 62.415000 15.420000 ;
        RECT 62.215000 15.660000 62.415000 15.860000 ;
        RECT 62.215000 16.100000 62.415000 16.300000 ;
        RECT 62.620000 13.020000 62.820000 13.220000 ;
        RECT 62.620000 13.460000 62.820000 13.660000 ;
        RECT 62.620000 13.900000 62.820000 14.100000 ;
        RECT 62.620000 14.340000 62.820000 14.540000 ;
        RECT 62.620000 14.780000 62.820000 14.980000 ;
        RECT 62.620000 15.220000 62.820000 15.420000 ;
        RECT 62.620000 15.660000 62.820000 15.860000 ;
        RECT 62.620000 16.100000 62.820000 16.300000 ;
        RECT 63.025000 13.020000 63.225000 13.220000 ;
        RECT 63.025000 13.460000 63.225000 13.660000 ;
        RECT 63.025000 13.900000 63.225000 14.100000 ;
        RECT 63.025000 14.340000 63.225000 14.540000 ;
        RECT 63.025000 14.780000 63.225000 14.980000 ;
        RECT 63.025000 15.220000 63.225000 15.420000 ;
        RECT 63.025000 15.660000 63.225000 15.860000 ;
        RECT 63.025000 16.100000 63.225000 16.300000 ;
        RECT 63.430000 13.020000 63.630000 13.220000 ;
        RECT 63.430000 13.460000 63.630000 13.660000 ;
        RECT 63.430000 13.900000 63.630000 14.100000 ;
        RECT 63.430000 14.340000 63.630000 14.540000 ;
        RECT 63.430000 14.780000 63.630000 14.980000 ;
        RECT 63.430000 15.220000 63.630000 15.420000 ;
        RECT 63.430000 15.660000 63.630000 15.860000 ;
        RECT 63.430000 16.100000 63.630000 16.300000 ;
        RECT 63.835000 13.020000 64.035000 13.220000 ;
        RECT 63.835000 13.460000 64.035000 13.660000 ;
        RECT 63.835000 13.900000 64.035000 14.100000 ;
        RECT 63.835000 14.340000 64.035000 14.540000 ;
        RECT 63.835000 14.780000 64.035000 14.980000 ;
        RECT 63.835000 15.220000 64.035000 15.420000 ;
        RECT 63.835000 15.660000 64.035000 15.860000 ;
        RECT 63.835000 16.100000 64.035000 16.300000 ;
        RECT 64.240000 13.020000 64.440000 13.220000 ;
        RECT 64.240000 13.460000 64.440000 13.660000 ;
        RECT 64.240000 13.900000 64.440000 14.100000 ;
        RECT 64.240000 14.340000 64.440000 14.540000 ;
        RECT 64.240000 14.780000 64.440000 14.980000 ;
        RECT 64.240000 15.220000 64.440000 15.420000 ;
        RECT 64.240000 15.660000 64.440000 15.860000 ;
        RECT 64.240000 16.100000 64.440000 16.300000 ;
        RECT 64.645000 13.020000 64.845000 13.220000 ;
        RECT 64.645000 13.460000 64.845000 13.660000 ;
        RECT 64.645000 13.900000 64.845000 14.100000 ;
        RECT 64.645000 14.340000 64.845000 14.540000 ;
        RECT 64.645000 14.780000 64.845000 14.980000 ;
        RECT 64.645000 15.220000 64.845000 15.420000 ;
        RECT 64.645000 15.660000 64.845000 15.860000 ;
        RECT 64.645000 16.100000 64.845000 16.300000 ;
        RECT 65.050000 13.020000 65.250000 13.220000 ;
        RECT 65.050000 13.460000 65.250000 13.660000 ;
        RECT 65.050000 13.900000 65.250000 14.100000 ;
        RECT 65.050000 14.340000 65.250000 14.540000 ;
        RECT 65.050000 14.780000 65.250000 14.980000 ;
        RECT 65.050000 15.220000 65.250000 15.420000 ;
        RECT 65.050000 15.660000 65.250000 15.860000 ;
        RECT 65.050000 16.100000 65.250000 16.300000 ;
        RECT 65.455000 13.020000 65.655000 13.220000 ;
        RECT 65.455000 13.460000 65.655000 13.660000 ;
        RECT 65.455000 13.900000 65.655000 14.100000 ;
        RECT 65.455000 14.340000 65.655000 14.540000 ;
        RECT 65.455000 14.780000 65.655000 14.980000 ;
        RECT 65.455000 15.220000 65.655000 15.420000 ;
        RECT 65.455000 15.660000 65.655000 15.860000 ;
        RECT 65.455000 16.100000 65.655000 16.300000 ;
        RECT 65.860000 13.020000 66.060000 13.220000 ;
        RECT 65.860000 13.460000 66.060000 13.660000 ;
        RECT 65.860000 13.900000 66.060000 14.100000 ;
        RECT 65.860000 14.340000 66.060000 14.540000 ;
        RECT 65.860000 14.780000 66.060000 14.980000 ;
        RECT 65.860000 15.220000 66.060000 15.420000 ;
        RECT 65.860000 15.660000 66.060000 15.860000 ;
        RECT 65.860000 16.100000 66.060000 16.300000 ;
        RECT 66.265000 13.020000 66.465000 13.220000 ;
        RECT 66.265000 13.460000 66.465000 13.660000 ;
        RECT 66.265000 13.900000 66.465000 14.100000 ;
        RECT 66.265000 14.340000 66.465000 14.540000 ;
        RECT 66.265000 14.780000 66.465000 14.980000 ;
        RECT 66.265000 15.220000 66.465000 15.420000 ;
        RECT 66.265000 15.660000 66.465000 15.860000 ;
        RECT 66.265000 16.100000 66.465000 16.300000 ;
        RECT 66.670000 13.020000 66.870000 13.220000 ;
        RECT 66.670000 13.460000 66.870000 13.660000 ;
        RECT 66.670000 13.900000 66.870000 14.100000 ;
        RECT 66.670000 14.340000 66.870000 14.540000 ;
        RECT 66.670000 14.780000 66.870000 14.980000 ;
        RECT 66.670000 15.220000 66.870000 15.420000 ;
        RECT 66.670000 15.660000 66.870000 15.860000 ;
        RECT 66.670000 16.100000 66.870000 16.300000 ;
        RECT 67.075000 13.020000 67.275000 13.220000 ;
        RECT 67.075000 13.460000 67.275000 13.660000 ;
        RECT 67.075000 13.900000 67.275000 14.100000 ;
        RECT 67.075000 14.340000 67.275000 14.540000 ;
        RECT 67.075000 14.780000 67.275000 14.980000 ;
        RECT 67.075000 15.220000 67.275000 15.420000 ;
        RECT 67.075000 15.660000 67.275000 15.860000 ;
        RECT 67.075000 16.100000 67.275000 16.300000 ;
        RECT 67.480000 13.020000 67.680000 13.220000 ;
        RECT 67.480000 13.460000 67.680000 13.660000 ;
        RECT 67.480000 13.900000 67.680000 14.100000 ;
        RECT 67.480000 14.340000 67.680000 14.540000 ;
        RECT 67.480000 14.780000 67.680000 14.980000 ;
        RECT 67.480000 15.220000 67.680000 15.420000 ;
        RECT 67.480000 15.660000 67.680000 15.860000 ;
        RECT 67.480000 16.100000 67.680000 16.300000 ;
        RECT 67.885000 13.020000 68.085000 13.220000 ;
        RECT 67.885000 13.460000 68.085000 13.660000 ;
        RECT 67.885000 13.900000 68.085000 14.100000 ;
        RECT 67.885000 14.340000 68.085000 14.540000 ;
        RECT 67.885000 14.780000 68.085000 14.980000 ;
        RECT 67.885000 15.220000 68.085000 15.420000 ;
        RECT 67.885000 15.660000 68.085000 15.860000 ;
        RECT 67.885000 16.100000 68.085000 16.300000 ;
        RECT 68.290000 13.020000 68.490000 13.220000 ;
        RECT 68.290000 13.460000 68.490000 13.660000 ;
        RECT 68.290000 13.900000 68.490000 14.100000 ;
        RECT 68.290000 14.340000 68.490000 14.540000 ;
        RECT 68.290000 14.780000 68.490000 14.980000 ;
        RECT 68.290000 15.220000 68.490000 15.420000 ;
        RECT 68.290000 15.660000 68.490000 15.860000 ;
        RECT 68.290000 16.100000 68.490000 16.300000 ;
        RECT 68.695000 13.020000 68.895000 13.220000 ;
        RECT 68.695000 13.460000 68.895000 13.660000 ;
        RECT 68.695000 13.900000 68.895000 14.100000 ;
        RECT 68.695000 14.340000 68.895000 14.540000 ;
        RECT 68.695000 14.780000 68.895000 14.980000 ;
        RECT 68.695000 15.220000 68.895000 15.420000 ;
        RECT 68.695000 15.660000 68.895000 15.860000 ;
        RECT 68.695000 16.100000 68.895000 16.300000 ;
        RECT 69.100000 13.020000 69.300000 13.220000 ;
        RECT 69.100000 13.460000 69.300000 13.660000 ;
        RECT 69.100000 13.900000 69.300000 14.100000 ;
        RECT 69.100000 14.340000 69.300000 14.540000 ;
        RECT 69.100000 14.780000 69.300000 14.980000 ;
        RECT 69.100000 15.220000 69.300000 15.420000 ;
        RECT 69.100000 15.660000 69.300000 15.860000 ;
        RECT 69.100000 16.100000 69.300000 16.300000 ;
        RECT 69.505000 13.020000 69.705000 13.220000 ;
        RECT 69.505000 13.460000 69.705000 13.660000 ;
        RECT 69.505000 13.900000 69.705000 14.100000 ;
        RECT 69.505000 14.340000 69.705000 14.540000 ;
        RECT 69.505000 14.780000 69.705000 14.980000 ;
        RECT 69.505000 15.220000 69.705000 15.420000 ;
        RECT 69.505000 15.660000 69.705000 15.860000 ;
        RECT 69.505000 16.100000 69.705000 16.300000 ;
        RECT 69.910000 13.020000 70.110000 13.220000 ;
        RECT 69.910000 13.460000 70.110000 13.660000 ;
        RECT 69.910000 13.900000 70.110000 14.100000 ;
        RECT 69.910000 14.340000 70.110000 14.540000 ;
        RECT 69.910000 14.780000 70.110000 14.980000 ;
        RECT 69.910000 15.220000 70.110000 15.420000 ;
        RECT 69.910000 15.660000 70.110000 15.860000 ;
        RECT 69.910000 16.100000 70.110000 16.300000 ;
        RECT 70.315000 13.020000 70.515000 13.220000 ;
        RECT 70.315000 13.460000 70.515000 13.660000 ;
        RECT 70.315000 13.900000 70.515000 14.100000 ;
        RECT 70.315000 14.340000 70.515000 14.540000 ;
        RECT 70.315000 14.780000 70.515000 14.980000 ;
        RECT 70.315000 15.220000 70.515000 15.420000 ;
        RECT 70.315000 15.660000 70.515000 15.860000 ;
        RECT 70.315000 16.100000 70.515000 16.300000 ;
        RECT 70.720000 13.020000 70.920000 13.220000 ;
        RECT 70.720000 13.460000 70.920000 13.660000 ;
        RECT 70.720000 13.900000 70.920000 14.100000 ;
        RECT 70.720000 14.340000 70.920000 14.540000 ;
        RECT 70.720000 14.780000 70.920000 14.980000 ;
        RECT 70.720000 15.220000 70.920000 15.420000 ;
        RECT 70.720000 15.660000 70.920000 15.860000 ;
        RECT 70.720000 16.100000 70.920000 16.300000 ;
        RECT 71.125000 13.020000 71.325000 13.220000 ;
        RECT 71.125000 13.460000 71.325000 13.660000 ;
        RECT 71.125000 13.900000 71.325000 14.100000 ;
        RECT 71.125000 14.340000 71.325000 14.540000 ;
        RECT 71.125000 14.780000 71.325000 14.980000 ;
        RECT 71.125000 15.220000 71.325000 15.420000 ;
        RECT 71.125000 15.660000 71.325000 15.860000 ;
        RECT 71.125000 16.100000 71.325000 16.300000 ;
        RECT 71.530000 13.020000 71.730000 13.220000 ;
        RECT 71.530000 13.460000 71.730000 13.660000 ;
        RECT 71.530000 13.900000 71.730000 14.100000 ;
        RECT 71.530000 14.340000 71.730000 14.540000 ;
        RECT 71.530000 14.780000 71.730000 14.980000 ;
        RECT 71.530000 15.220000 71.730000 15.420000 ;
        RECT 71.530000 15.660000 71.730000 15.860000 ;
        RECT 71.530000 16.100000 71.730000 16.300000 ;
        RECT 71.935000 13.020000 72.135000 13.220000 ;
        RECT 71.935000 13.460000 72.135000 13.660000 ;
        RECT 71.935000 13.900000 72.135000 14.100000 ;
        RECT 71.935000 14.340000 72.135000 14.540000 ;
        RECT 71.935000 14.780000 72.135000 14.980000 ;
        RECT 71.935000 15.220000 72.135000 15.420000 ;
        RECT 71.935000 15.660000 72.135000 15.860000 ;
        RECT 71.935000 16.100000 72.135000 16.300000 ;
        RECT 72.340000 13.020000 72.540000 13.220000 ;
        RECT 72.340000 13.460000 72.540000 13.660000 ;
        RECT 72.340000 13.900000 72.540000 14.100000 ;
        RECT 72.340000 14.340000 72.540000 14.540000 ;
        RECT 72.340000 14.780000 72.540000 14.980000 ;
        RECT 72.340000 15.220000 72.540000 15.420000 ;
        RECT 72.340000 15.660000 72.540000 15.860000 ;
        RECT 72.340000 16.100000 72.540000 16.300000 ;
        RECT 72.745000 13.020000 72.945000 13.220000 ;
        RECT 72.745000 13.460000 72.945000 13.660000 ;
        RECT 72.745000 13.900000 72.945000 14.100000 ;
        RECT 72.745000 14.340000 72.945000 14.540000 ;
        RECT 72.745000 14.780000 72.945000 14.980000 ;
        RECT 72.745000 15.220000 72.945000 15.420000 ;
        RECT 72.745000 15.660000 72.945000 15.860000 ;
        RECT 72.745000 16.100000 72.945000 16.300000 ;
        RECT 73.150000 13.020000 73.350000 13.220000 ;
        RECT 73.150000 13.460000 73.350000 13.660000 ;
        RECT 73.150000 13.900000 73.350000 14.100000 ;
        RECT 73.150000 14.340000 73.350000 14.540000 ;
        RECT 73.150000 14.780000 73.350000 14.980000 ;
        RECT 73.150000 15.220000 73.350000 15.420000 ;
        RECT 73.150000 15.660000 73.350000 15.860000 ;
        RECT 73.150000 16.100000 73.350000 16.300000 ;
        RECT 73.555000 13.020000 73.755000 13.220000 ;
        RECT 73.555000 13.460000 73.755000 13.660000 ;
        RECT 73.555000 13.900000 73.755000 14.100000 ;
        RECT 73.555000 14.340000 73.755000 14.540000 ;
        RECT 73.555000 14.780000 73.755000 14.980000 ;
        RECT 73.555000 15.220000 73.755000 15.420000 ;
        RECT 73.555000 15.660000 73.755000 15.860000 ;
        RECT 73.555000 16.100000 73.755000 16.300000 ;
        RECT 73.960000 13.020000 74.160000 13.220000 ;
        RECT 73.960000 13.460000 74.160000 13.660000 ;
        RECT 73.960000 13.900000 74.160000 14.100000 ;
        RECT 73.960000 14.340000 74.160000 14.540000 ;
        RECT 73.960000 14.780000 74.160000 14.980000 ;
        RECT 73.960000 15.220000 74.160000 15.420000 ;
        RECT 73.960000 15.660000 74.160000 15.860000 ;
        RECT 73.960000 16.100000 74.160000 16.300000 ;
        RECT 74.365000 13.020000 74.565000 13.220000 ;
        RECT 74.365000 13.460000 74.565000 13.660000 ;
        RECT 74.365000 13.900000 74.565000 14.100000 ;
        RECT 74.365000 14.340000 74.565000 14.540000 ;
        RECT 74.365000 14.780000 74.565000 14.980000 ;
        RECT 74.365000 15.220000 74.565000 15.420000 ;
        RECT 74.365000 15.660000 74.565000 15.860000 ;
        RECT 74.365000 16.100000 74.565000 16.300000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 75.000000  12.540000 ;
      RECT  0.000000 16.780000 75.000000 198.000000 ;
      RECT 24.900000 12.540000 50.355000  16.780000 ;
    LAYER met4 ;
      RECT  0.000000   5.885000  1.670000   6.485000 ;
      RECT  0.000000  11.935000  1.670000  12.535000 ;
      RECT  0.000000  16.785000  1.670000  17.385000 ;
      RECT  0.000000  22.835000  1.670000  23.435000 ;
      RECT  0.000000  28.885000  1.670000  29.485000 ;
      RECT  0.000000  33.735000  1.670000  34.335000 ;
      RECT  0.000000  38.585000  1.670000  39.185000 ;
      RECT  0.000000  44.635000  1.670000  45.335000 ;
      RECT  0.000000  55.135000  1.670000  55.835000 ;
      RECT  0.000000  61.085000  1.670000  61.685000 ;
      RECT  0.000000  66.935000  1.670000  67.635000 ;
      RECT  0.000000  93.400000 75.000000 173.385000 ;
      RECT  1.670000   0.000000 73.330000  12.535000 ;
      RECT  1.670000  16.785000 73.330000  93.400000 ;
      RECT  1.670000 173.385000 73.330000 198.000000 ;
      RECT 24.875000  12.535000 50.380000  16.785000 ;
      RECT 73.330000   5.885000 75.000000   6.485000 ;
      RECT 73.330000  11.935000 75.000000  12.535000 ;
      RECT 73.330000  16.785000 75.000000  17.385000 ;
      RECT 73.330000  22.835000 75.000000  23.435000 ;
      RECT 73.330000  28.885000 75.000000  29.485000 ;
      RECT 73.330000  33.735000 75.000000  34.335000 ;
      RECT 73.330000  38.585000 75.000000  39.185000 ;
      RECT 73.330000  44.635000 75.000000  45.335000 ;
      RECT 73.330000  55.135000 75.000000  55.835000 ;
      RECT 73.330000  61.085000 75.000000  61.685000 ;
      RECT 73.330000  66.935000 75.000000  67.635000 ;
    LAYER met5 ;
      RECT 0.000000  93.785000 75.000000 172.985000 ;
      RECT 1.765000  12.235000 73.235000  17.085000 ;
      RECT 2.070000   0.000000 72.930000  12.235000 ;
      RECT 2.070000  17.085000 72.930000  93.785000 ;
      RECT 2.070000 172.985000 72.930000 198.000000 ;
  END
END sky130_fd_io__overlay_vdda_lvc


MACRO sky130_fd_io__top_gpiov2
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 80 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  119.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 53.125000 80.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  119.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 48.365000 80.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN ANALOG_EN
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.430000 0.000000 62.690000 1.915000 ;
    END
  END ANALOG_EN
  PIN ANALOG_POL
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.865000  0.000000 46.195000 36.665000 ;
        RECT 45.865000 36.665000 46.195000 36.735000 ;
        RECT 45.865000 36.735000 46.265000 36.805000 ;
        RECT 45.965000 36.805000 46.335000 36.905000 ;
        RECT 46.065000 36.905000 46.435000 37.005000 ;
        RECT 46.070000 37.005000 46.535000 37.010000 ;
        RECT 46.220000 37.010000 48.225000 37.160000 ;
        RECT 46.370000 37.160000 48.075000 37.310000 ;
        RECT 46.400000 37.310000 48.045000 37.340000 ;
        RECT 47.910000 37.005000 48.375000 37.010000 ;
        RECT 47.960000 35.870000 48.740000 36.190000 ;
        RECT 47.975000 36.940000 48.380000 37.005000 ;
        RECT 48.040000 36.875000 48.445000 36.940000 ;
        RECT 48.070000 36.190000 48.630000 36.300000 ;
        RECT 48.110000 36.805000 48.510000 36.875000 ;
        RECT 48.180000 36.300000 48.520000 36.410000 ;
        RECT 48.180000 36.410000 48.515000 36.415000 ;
        RECT 48.180000 36.415000 48.510000 36.420000 ;
        RECT 48.180000 36.420000 48.510000 36.735000 ;
        RECT 48.180000 36.735000 48.510000 36.805000 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.080000 57.360000 24.590000 57.430000 ;
        RECT 23.080000 57.430000 24.520000 57.500000 ;
        RECT 23.080000 57.500000 24.450000 57.570000 ;
        RECT 23.080000 57.570000 24.380000 57.640000 ;
        RECT 24.285000 57.345000 24.660000 57.360000 ;
        RECT 24.355000 57.275000 24.675000 57.345000 ;
        RECT 24.425000 57.205000 24.745000 57.275000 ;
        RECT 24.495000 57.135000 24.815000 57.205000 ;
        RECT 24.565000 57.065000 24.885000 57.135000 ;
        RECT 24.620000 57.010000 24.955000 57.065000 ;
        RECT 24.675000 53.255000 25.010000 53.310000 ;
        RECT 24.675000 53.310000 24.955000 53.365000 ;
        RECT 24.675000 53.365000 24.955000 56.955000 ;
        RECT 24.675000 56.955000 24.955000 57.010000 ;
        RECT 24.740000 53.190000 25.065000 53.255000 ;
        RECT 24.810000 53.120000 25.130000 53.190000 ;
        RECT 24.880000 53.050000 25.200000 53.120000 ;
        RECT 24.950000 52.980000 25.270000 53.050000 ;
        RECT 25.020000 52.910000 25.340000 52.980000 ;
        RECT 25.090000 52.840000 25.410000 52.910000 ;
        RECT 25.160000 52.770000 25.480000 52.840000 ;
        RECT 25.230000 52.700000 25.550000 52.770000 ;
        RECT 25.300000 52.630000 25.620000 52.700000 ;
        RECT 25.370000 52.560000 25.690000 52.630000 ;
        RECT 25.440000 52.490000 25.760000 52.560000 ;
        RECT 25.510000 52.420000 25.830000 52.490000 ;
        RECT 25.580000 52.350000 25.900000 52.420000 ;
        RECT 25.650000 52.280000 25.970000 52.350000 ;
        RECT 25.720000 52.210000 26.040000 52.280000 ;
        RECT 25.790000 52.140000 29.735000 52.210000 ;
        RECT 25.860000 52.070000 29.805000 52.140000 ;
        RECT 25.930000 52.000000 29.875000 52.070000 ;
        RECT 26.000000 51.930000 29.945000 52.000000 ;
        RECT 29.645000 51.910000 30.015000 51.930000 ;
        RECT 29.715000 51.840000 30.035000 51.910000 ;
        RECT 29.785000 51.770000 30.105000 51.840000 ;
        RECT 29.855000 51.700000 30.175000 51.770000 ;
        RECT 29.925000 51.630000 30.245000 51.700000 ;
        RECT 29.995000 51.560000 30.315000 51.630000 ;
        RECT 30.060000 51.495000 30.385000 51.560000 ;
        RECT 30.125000 17.630000 30.440000 17.685000 ;
        RECT 30.125000 17.685000 30.385000 17.740000 ;
        RECT 30.125000 17.740000 30.385000 36.345000 ;
        RECT 30.125000 36.345000 30.385000 36.400000 ;
        RECT 30.125000 36.400000 30.440000 36.455000 ;
        RECT 30.125000 38.010000 30.440000 38.065000 ;
        RECT 30.125000 38.065000 30.385000 38.120000 ;
        RECT 30.125000 38.120000 30.385000 51.430000 ;
        RECT 30.125000 51.430000 30.385000 51.495000 ;
        RECT 30.140000 37.995000 30.495000 38.010000 ;
        RECT 30.180000 17.575000 30.495000 17.630000 ;
        RECT 30.195000 36.455000 30.495000 36.525000 ;
        RECT 30.210000 37.925000 30.510000 37.995000 ;
        RECT 30.250000 17.505000 30.550000 17.575000 ;
        RECT 30.265000 36.525000 30.565000 36.595000 ;
        RECT 30.280000 36.595000 30.635000 36.610000 ;
        RECT 30.280000 37.855000 30.580000 37.925000 ;
        RECT 30.320000 17.435000 30.620000 17.505000 ;
        RECT 30.335000 36.610000 30.650000 36.665000 ;
        RECT 30.335000 37.800000 30.650000 37.855000 ;
        RECT 30.390000 17.365000 30.690000 17.435000 ;
        RECT 30.390000 36.665000 30.650000 36.720000 ;
        RECT 30.390000 36.720000 30.650000 37.745000 ;
        RECT 30.390000 37.745000 30.650000 37.800000 ;
        RECT 30.460000 17.295000 30.760000 17.365000 ;
        RECT 30.530000 17.225000 30.830000 17.295000 ;
        RECT 30.600000 17.155000 30.900000 17.225000 ;
        RECT 30.670000 17.085000 30.970000 17.155000 ;
        RECT 30.740000 17.015000 31.040000 17.085000 ;
        RECT 30.750000  0.000000 31.010000  2.155000 ;
        RECT 30.750000  2.155000 31.010000  2.210000 ;
        RECT 30.750000  2.210000 31.065000  2.265000 ;
        RECT 30.810000 16.945000 31.110000 17.015000 ;
        RECT 30.820000  2.265000 31.120000  2.335000 ;
        RECT 30.880000 16.875000 31.180000 16.945000 ;
        RECT 30.890000  2.335000 31.190000  2.405000 ;
        RECT 30.950000 16.805000 31.250000 16.875000 ;
        RECT 30.960000  2.405000 31.260000  2.475000 ;
        RECT 31.020000 16.735000 31.320000 16.805000 ;
        RECT 31.030000  2.475000 31.330000  2.545000 ;
        RECT 31.090000 16.665000 31.390000 16.735000 ;
        RECT 31.100000  2.545000 31.400000  2.615000 ;
        RECT 31.160000 16.595000 31.460000 16.665000 ;
        RECT 31.170000  2.615000 31.470000  2.685000 ;
        RECT 31.195000  2.685000 31.540000  2.710000 ;
        RECT 31.230000 16.525000 31.530000 16.595000 ;
        RECT 31.250000  2.710000 31.565000  2.765000 ;
        RECT 31.300000 16.455000 31.600000 16.525000 ;
        RECT 31.305000  2.765000 31.565000  2.820000 ;
        RECT 31.305000  2.820000 31.565000  4.335000 ;
        RECT 31.305000  4.335000 31.565000  4.390000 ;
        RECT 31.305000  4.390000 31.620000  4.445000 ;
        RECT 31.370000 16.385000 31.670000 16.455000 ;
        RECT 31.375000  4.445000 31.675000  4.515000 ;
        RECT 31.440000 16.315000 31.740000 16.385000 ;
        RECT 31.445000  4.515000 31.745000  4.585000 ;
        RECT 31.510000 16.245000 31.810000 16.315000 ;
        RECT 31.515000  4.585000 31.815000  4.655000 ;
        RECT 31.580000  4.655000 31.885000  4.720000 ;
        RECT 31.580000 16.175000 31.880000 16.245000 ;
        RECT 31.635000  4.720000 31.950000  4.775000 ;
        RECT 31.635000 16.120000 31.950000 16.175000 ;
        RECT 31.690000  4.775000 31.950000  4.830000 ;
        RECT 31.690000  4.830000 31.950000 16.065000 ;
        RECT 31.690000 16.065000 31.950000 16.120000 ;
    END
  END ANALOG_SEL
  PIN DM[0]
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.590000 0.545000 50.360000 0.825000 ;
        RECT 49.625000 0.510000 50.325000 0.545000 ;
        RECT 49.695000 0.440000 50.255000 0.510000 ;
        RECT 49.765000 0.370000 50.185000 0.440000 ;
        RECT 49.835000 0.300000 50.115000 0.370000 ;
        RECT 49.845000 0.290000 50.115000 0.300000 ;
        RECT 49.855000 0.000000 50.115000 0.280000 ;
        RECT 49.855000 0.280000 50.115000 0.290000 ;
    END
  END DM[0]
  PIN DM[1]
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.540000 1.195000 67.360000 1.475000 ;
        RECT 66.595000 1.140000 67.305000 1.195000 ;
        RECT 66.665000 1.070000 67.235000 1.140000 ;
        RECT 66.735000 1.000000 67.165000 1.070000 ;
        RECT 66.805000 0.930000 67.095000 1.000000 ;
        RECT 66.820000 0.915000 67.095000 0.930000 ;
        RECT 66.835000 0.000000 67.095000 0.900000 ;
        RECT 66.835000 0.900000 67.095000 0.915000 ;
    END
  END DM[1]
  PIN DM[2]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.490000 0.000000 28.750000 3.960000 ;
        RECT 28.490000 3.960000 28.750000 4.015000 ;
        RECT 28.490000 4.015000 28.805000 4.070000 ;
        RECT 28.560000 4.070000 28.860000 4.140000 ;
        RECT 28.630000 4.140000 28.930000 4.210000 ;
        RECT 28.700000 4.210000 29.000000 4.280000 ;
        RECT 28.770000 4.280000 29.070000 4.350000 ;
        RECT 28.840000 4.350000 29.140000 4.420000 ;
        RECT 28.910000 4.420000 29.210000 4.490000 ;
        RECT 28.980000 4.490000 29.280000 4.560000 ;
        RECT 29.050000 4.560000 29.350000 4.630000 ;
        RECT 29.100000 4.630000 29.420000 4.680000 ;
        RECT 29.155000 4.680000 29.470000 4.735000 ;
        RECT 29.210000 4.735000 29.470000 4.790000 ;
        RECT 29.210000 4.790000 29.470000 6.780000 ;
    END
  END DM[2]
  PIN ENABLE_H
    ANTENNAGATEAREA  4.860000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.135000 2.225000 35.450000 2.280000 ;
        RECT 35.135000 2.280000 35.395000 2.335000 ;
        RECT 35.135000 2.335000 35.395000 3.885000 ;
        RECT 35.140000 2.220000 35.505000 2.225000 ;
        RECT 35.210000 2.150000 35.510000 2.220000 ;
        RECT 35.280000 2.080000 35.580000 2.150000 ;
        RECT 35.350000 2.010000 35.650000 2.080000 ;
        RECT 35.405000 1.955000 35.720000 2.010000 ;
        RECT 35.460000 0.000000 35.720000 1.900000 ;
        RECT 35.460000 1.900000 35.720000 1.955000 ;
    END
  END ENABLE_H
  PIN ENABLE_INP_H
    ANTENNAGATEAREA  3.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.390000 0.000000 38.650000 3.715000 ;
    END
  END ENABLE_INP_H
  PIN ENABLE_VDDA_H
    ANTENNAGATEAREA  3.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  7.315000 56.460000  7.630000 56.515000 ;
        RECT  7.315000 56.515000  7.575000 56.570000 ;
        RECT  7.315000 56.570000  7.575000 73.615000 ;
        RECT  7.315000 73.615000  7.575000 73.670000 ;
        RECT  7.315000 73.670000  7.630000 73.725000 ;
        RECT  7.375000 56.400000  7.685000 56.460000 ;
        RECT  7.385000 73.725000  7.685000 73.795000 ;
        RECT  7.445000 56.330000  7.745000 56.400000 ;
        RECT  7.455000 73.795000  7.755000 73.865000 ;
        RECT  7.515000 56.260000  7.815000 56.330000 ;
        RECT  7.525000 73.865000  7.825000 73.935000 ;
        RECT  7.585000 56.190000  7.885000 56.260000 ;
        RECT  7.595000 73.935000  7.895000 74.005000 ;
        RECT  7.655000 56.120000  7.955000 56.190000 ;
        RECT  7.665000 74.005000  7.965000 74.075000 ;
        RECT  7.695000 74.075000  8.035000 74.105000 ;
        RECT  7.725000 56.050000  8.025000 56.120000 ;
        RECT  7.750000 74.105000  8.065000 74.160000 ;
        RECT  7.795000 55.980000  8.095000 56.050000 ;
        RECT  7.805000 74.160000  8.065000 74.215000 ;
        RECT  7.805000 74.215000  8.065000 74.680000 ;
        RECT  7.805000 74.680000  8.065000 74.735000 ;
        RECT  7.805000 74.735000  8.120000 74.790000 ;
        RECT  7.865000 55.910000  8.165000 55.980000 ;
        RECT  7.875000 74.790000  8.175000 74.860000 ;
        RECT  7.920000 55.855000  8.235000 55.910000 ;
        RECT  7.920000 77.285000  8.560000 77.545000 ;
        RECT  7.945000 74.860000  8.245000 74.930000 ;
        RECT  7.975000 53.960000  8.290000 54.015000 ;
        RECT  7.975000 54.015000  8.235000 54.070000 ;
        RECT  7.975000 54.070000  8.235000 55.800000 ;
        RECT  7.975000 55.800000  8.235000 55.855000 ;
        RECT  8.015000 74.930000  8.315000 75.000000 ;
        RECT  8.030000 53.905000  8.345000 53.960000 ;
        RECT  8.085000 53.850000  8.400000 53.905000 ;
        RECT  8.085000 75.000000  8.385000 75.070000 ;
        RECT  8.085000 77.240000  8.515000 77.285000 ;
        RECT  8.100000 75.070000  8.455000 75.085000 ;
        RECT  8.130000 77.195000  8.470000 77.240000 ;
        RECT  8.140000 53.795000  8.455000 53.850000 ;
        RECT  8.155000 75.085000  8.470000 75.140000 ;
        RECT  8.170000 77.155000  8.470000 77.195000 ;
        RECT  8.195000 44.075000  8.510000 44.130000 ;
        RECT  8.195000 44.130000  8.455000 44.185000 ;
        RECT  8.195000 44.185000  8.455000 53.740000 ;
        RECT  8.195000 53.740000  8.455000 53.795000 ;
        RECT  8.210000 44.060000  8.565000 44.075000 ;
        RECT  8.210000 75.140000  8.470000 75.195000 ;
        RECT  8.210000 75.195000  8.470000 77.115000 ;
        RECT  8.210000 77.115000  8.470000 77.155000 ;
        RECT  8.280000 43.990000  8.580000 44.060000 ;
        RECT  8.350000 43.920000  8.650000 43.990000 ;
        RECT  8.420000 43.850000  8.720000 43.920000 ;
        RECT  8.490000 43.780000  8.790000 43.850000 ;
        RECT  8.560000 43.710000  8.860000 43.780000 ;
        RECT  8.630000 43.640000  8.930000 43.710000 ;
        RECT  8.700000 43.570000  9.000000 43.640000 ;
        RECT  8.770000 43.500000  9.070000 43.570000 ;
        RECT  8.840000 43.430000  9.140000 43.500000 ;
        RECT  8.910000 43.360000  9.210000 43.430000 ;
        RECT  8.980000 43.290000  9.280000 43.360000 ;
        RECT  9.050000 43.220000  9.350000 43.290000 ;
        RECT  9.120000 43.150000  9.420000 43.220000 ;
        RECT  9.190000 43.080000  9.490000 43.150000 ;
        RECT  9.260000 43.010000  9.560000 43.080000 ;
        RECT  9.330000 42.940000  9.630000 43.010000 ;
        RECT  9.400000 42.870000  9.700000 42.940000 ;
        RECT  9.470000 42.800000  9.770000 42.870000 ;
        RECT  9.540000 42.730000  9.840000 42.800000 ;
        RECT  9.610000 42.660000  9.910000 42.730000 ;
        RECT  9.680000 42.590000  9.980000 42.660000 ;
        RECT  9.750000 42.520000 10.050000 42.590000 ;
        RECT  9.820000 42.450000 10.120000 42.520000 ;
        RECT  9.890000 42.380000 10.190000 42.450000 ;
        RECT  9.960000 42.310000 10.260000 42.380000 ;
        RECT 10.030000 42.240000 10.330000 42.310000 ;
        RECT 10.100000 42.170000 10.400000 42.240000 ;
        RECT 10.170000 42.100000 10.470000 42.170000 ;
        RECT 10.240000 42.030000 10.540000 42.100000 ;
        RECT 10.310000 41.960000 10.610000 42.030000 ;
        RECT 10.380000 41.890000 10.680000 41.960000 ;
        RECT 10.450000 41.820000 10.750000 41.890000 ;
        RECT 10.520000 41.750000 10.820000 41.820000 ;
        RECT 10.590000 41.680000 10.890000 41.750000 ;
        RECT 10.660000 41.610000 10.960000 41.680000 ;
        RECT 10.730000 41.540000 11.030000 41.610000 ;
        RECT 10.800000 41.470000 11.100000 41.540000 ;
        RECT 10.870000 41.400000 11.170000 41.470000 ;
        RECT 10.940000 41.330000 11.240000 41.400000 ;
        RECT 11.010000 41.260000 11.310000 41.330000 ;
        RECT 11.080000 41.190000 11.380000 41.260000 ;
        RECT 11.150000 41.120000 11.450000 41.190000 ;
        RECT 11.220000 41.050000 11.520000 41.120000 ;
        RECT 11.290000 40.980000 11.590000 41.050000 ;
        RECT 11.360000 40.910000 11.660000 40.980000 ;
        RECT 11.430000 40.840000 11.730000 40.910000 ;
        RECT 11.500000 40.770000 11.800000 40.840000 ;
        RECT 11.570000 40.700000 11.870000 40.770000 ;
        RECT 11.640000 40.630000 11.940000 40.700000 ;
        RECT 11.710000 40.560000 12.010000 40.630000 ;
        RECT 11.780000 40.490000 12.080000 40.560000 ;
        RECT 11.850000 40.420000 12.150000 40.490000 ;
        RECT 11.920000 40.350000 12.220000 40.420000 ;
        RECT 11.990000 40.280000 12.290000 40.350000 ;
        RECT 12.060000 40.210000 12.360000 40.280000 ;
        RECT 12.130000 40.140000 12.430000 40.210000 ;
        RECT 12.200000 40.070000 12.500000 40.140000 ;
        RECT 12.270000 40.000000 12.570000 40.070000 ;
        RECT 12.340000 39.930000 12.640000 40.000000 ;
        RECT 12.410000 39.860000 12.710000 39.930000 ;
        RECT 12.480000 39.790000 12.780000 39.860000 ;
        RECT 12.550000 39.720000 12.850000 39.790000 ;
        RECT 12.620000 39.650000 12.920000 39.720000 ;
        RECT 12.690000 39.580000 12.990000 39.650000 ;
        RECT 12.755000  0.000000 13.015000  5.240000 ;
        RECT 12.755000  5.240000 13.015000  5.295000 ;
        RECT 12.755000  5.295000 13.070000  5.350000 ;
        RECT 12.760000 39.510000 13.060000 39.580000 ;
        RECT 12.825000  5.350000 13.125000  5.420000 ;
        RECT 12.830000 39.440000 13.130000 39.510000 ;
        RECT 12.895000  5.420000 13.195000  5.490000 ;
        RECT 12.900000 39.370000 13.200000 39.440000 ;
        RECT 12.965000  5.490000 13.265000  5.560000 ;
        RECT 12.970000 39.300000 13.270000 39.370000 ;
        RECT 13.035000  5.560000 13.335000  5.630000 ;
        RECT 13.040000 39.230000 13.340000 39.300000 ;
        RECT 13.105000  5.630000 13.405000  5.700000 ;
        RECT 13.110000 39.160000 13.410000 39.230000 ;
        RECT 13.175000  5.700000 13.475000  5.770000 ;
        RECT 13.180000 39.090000 13.480000 39.160000 ;
        RECT 13.245000  5.770000 13.545000  5.840000 ;
        RECT 13.250000 39.020000 13.550000 39.090000 ;
        RECT 13.315000  5.840000 13.615000  5.910000 ;
        RECT 13.320000 38.950000 13.620000 39.020000 ;
        RECT 13.385000  5.910000 13.685000  5.980000 ;
        RECT 13.390000 38.880000 13.690000 38.950000 ;
        RECT 13.455000  5.980000 13.755000  6.050000 ;
        RECT 13.460000 38.810000 13.760000 38.880000 ;
        RECT 13.525000  6.050000 13.825000  6.120000 ;
        RECT 13.530000 38.740000 13.830000 38.810000 ;
        RECT 13.595000  6.120000 13.895000  6.190000 ;
        RECT 13.600000 38.670000 13.900000 38.740000 ;
        RECT 13.665000  6.190000 13.965000  6.260000 ;
        RECT 13.670000 38.600000 13.970000 38.670000 ;
        RECT 13.735000  6.260000 14.035000  6.330000 ;
        RECT 13.740000 38.530000 14.040000 38.600000 ;
        RECT 13.805000  6.330000 14.105000  6.400000 ;
        RECT 13.810000 38.460000 14.110000 38.530000 ;
        RECT 13.860000  6.400000 14.175000  6.455000 ;
        RECT 13.880000 38.390000 14.180000 38.460000 ;
        RECT 13.915000  6.455000 14.230000  6.510000 ;
        RECT 13.950000 38.320000 14.250000 38.390000 ;
        RECT 13.970000  6.510000 14.230000  6.565000 ;
        RECT 13.970000  6.565000 14.230000 18.115000 ;
        RECT 13.970000 18.115000 14.230000 18.170000 ;
        RECT 13.970000 18.170000 14.285000 18.225000 ;
        RECT 14.020000 38.250000 14.320000 38.320000 ;
        RECT 14.040000 18.225000 14.340000 18.295000 ;
        RECT 14.090000 38.180000 14.390000 38.250000 ;
        RECT 14.110000 18.295000 14.410000 18.365000 ;
        RECT 14.160000 38.110000 14.460000 38.180000 ;
        RECT 14.180000 18.365000 14.480000 18.435000 ;
        RECT 14.230000 38.040000 14.530000 38.110000 ;
        RECT 14.250000 18.435000 14.550000 18.505000 ;
        RECT 14.300000 37.970000 14.600000 38.040000 ;
        RECT 14.320000 18.505000 14.620000 18.575000 ;
        RECT 14.370000 37.900000 14.670000 37.970000 ;
        RECT 14.390000 18.575000 14.690000 18.645000 ;
        RECT 14.440000 37.830000 14.740000 37.900000 ;
        RECT 14.460000 18.645000 14.760000 18.715000 ;
        RECT 14.510000 37.760000 14.810000 37.830000 ;
        RECT 14.530000 18.715000 14.830000 18.785000 ;
        RECT 14.580000 37.690000 14.880000 37.760000 ;
        RECT 14.600000 18.785000 14.900000 18.855000 ;
        RECT 14.650000 37.620000 14.950000 37.690000 ;
        RECT 14.670000 18.855000 14.970000 18.925000 ;
        RECT 14.720000 37.550000 15.020000 37.620000 ;
        RECT 14.740000 18.925000 15.040000 18.995000 ;
        RECT 14.790000 37.480000 15.090000 37.550000 ;
        RECT 14.810000 18.995000 15.110000 19.065000 ;
        RECT 14.860000 37.410000 15.160000 37.480000 ;
        RECT 14.880000 19.065000 15.180000 19.135000 ;
        RECT 14.915000 37.355000 15.230000 37.410000 ;
        RECT 14.950000 19.135000 15.250000 19.205000 ;
        RECT 14.970000 31.960000 15.285000 32.015000 ;
        RECT 14.970000 32.015000 15.230000 32.070000 ;
        RECT 14.970000 32.070000 15.230000 37.300000 ;
        RECT 14.970000 37.300000 15.230000 37.355000 ;
        RECT 14.995000 31.935000 15.340000 31.960000 ;
        RECT 15.020000 19.205000 15.320000 19.275000 ;
        RECT 15.065000 31.865000 15.365000 31.935000 ;
        RECT 15.090000 19.275000 15.390000 19.345000 ;
        RECT 15.135000 31.795000 15.435000 31.865000 ;
        RECT 15.160000 19.345000 15.460000 19.415000 ;
        RECT 15.205000 31.725000 15.505000 31.795000 ;
        RECT 15.230000 19.415000 15.530000 19.485000 ;
        RECT 15.275000 19.485000 15.600000 19.530000 ;
        RECT 15.275000 31.655000 15.575000 31.725000 ;
        RECT 15.330000 19.530000 15.645000 19.585000 ;
        RECT 15.330000 31.600000 15.645000 31.655000 ;
        RECT 15.385000 19.585000 15.645000 19.640000 ;
        RECT 15.385000 19.640000 15.645000 31.545000 ;
        RECT 15.385000 31.545000 15.645000 31.600000 ;
    END
  END ENABLE_VDDA_H
  PIN ENABLE_VDDIO
    ANTENNAGATEAREA  3.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.580000 0.000000 78.910000 176.480000 ;
    END
  END ENABLE_VDDIO
  PIN ENABLE_VSWITCH_H
    ANTENNAGATEAREA  3.120000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.250000 43.835000 11.565000 43.890000 ;
        RECT 11.250000 43.890000 11.510000 43.945000 ;
        RECT 11.250000 43.945000 11.510000 47.275000 ;
        RECT 11.250000 47.275000 11.510000 47.330000 ;
        RECT 11.250000 47.330000 11.565000 47.385000 ;
        RECT 11.270000 43.815000 11.620000 43.835000 ;
        RECT 11.320000 47.385000 11.620000 47.455000 ;
        RECT 11.340000 43.745000 11.640000 43.815000 ;
        RECT 11.390000 47.455000 11.690000 47.525000 ;
        RECT 11.410000 43.675000 11.710000 43.745000 ;
        RECT 11.460000 47.525000 11.760000 47.595000 ;
        RECT 11.480000 43.605000 11.780000 43.675000 ;
        RECT 11.530000 47.595000 11.830000 47.665000 ;
        RECT 11.550000 43.535000 11.850000 43.605000 ;
        RECT 11.600000 47.665000 11.900000 47.735000 ;
        RECT 11.620000 43.465000 11.920000 43.535000 ;
        RECT 11.670000 47.735000 11.970000 47.805000 ;
        RECT 11.680000 47.805000 12.040000 47.815000 ;
        RECT 11.690000 43.395000 11.990000 43.465000 ;
        RECT 11.750000 47.815000 13.850000 47.885000 ;
        RECT 11.760000 43.325000 12.060000 43.395000 ;
        RECT 11.820000 47.885000 13.920000 47.955000 ;
        RECT 11.830000 43.255000 12.130000 43.325000 ;
        RECT 11.890000 47.955000 13.990000 48.025000 ;
        RECT 11.900000 43.185000 12.200000 43.255000 ;
        RECT 11.940000 48.025000 14.060000 48.075000 ;
        RECT 11.970000 43.115000 12.270000 43.185000 ;
        RECT 12.040000 43.045000 12.340000 43.115000 ;
        RECT 12.110000 42.975000 12.410000 43.045000 ;
        RECT 12.180000 42.905000 12.480000 42.975000 ;
        RECT 12.250000 42.835000 12.550000 42.905000 ;
        RECT 12.320000 42.765000 12.620000 42.835000 ;
        RECT 12.390000 42.695000 12.690000 42.765000 ;
        RECT 12.460000 42.625000 12.760000 42.695000 ;
        RECT 12.530000 42.555000 12.830000 42.625000 ;
        RECT 12.600000 42.485000 12.900000 42.555000 ;
        RECT 12.670000 42.415000 12.970000 42.485000 ;
        RECT 12.740000 42.345000 13.040000 42.415000 ;
        RECT 12.810000 42.275000 13.110000 42.345000 ;
        RECT 12.880000 42.205000 13.180000 42.275000 ;
        RECT 12.950000 42.135000 13.250000 42.205000 ;
        RECT 13.020000 42.065000 13.320000 42.135000 ;
        RECT 13.090000 41.995000 13.390000 42.065000 ;
        RECT 13.160000 41.925000 13.460000 41.995000 ;
        RECT 13.230000 41.855000 13.530000 41.925000 ;
        RECT 13.300000 41.785000 13.600000 41.855000 ;
        RECT 13.370000 41.715000 13.670000 41.785000 ;
        RECT 13.440000 41.645000 13.740000 41.715000 ;
        RECT 13.510000 41.575000 13.810000 41.645000 ;
        RECT 13.565000 41.520000 13.880000 41.575000 ;
        RECT 13.620000 40.430000 13.935000 40.485000 ;
        RECT 13.620000 40.485000 13.880000 40.540000 ;
        RECT 13.620000 40.540000 13.880000 41.465000 ;
        RECT 13.620000 41.465000 13.880000 41.520000 ;
        RECT 13.640000 40.410000 13.990000 40.430000 ;
        RECT 13.710000 40.340000 14.010000 40.410000 ;
        RECT 13.780000 40.270000 14.080000 40.340000 ;
        RECT 13.810000 48.075000 14.110000 48.145000 ;
        RECT 13.850000 40.200000 14.150000 40.270000 ;
        RECT 13.880000 48.145000 14.180000 48.215000 ;
        RECT 13.920000 40.130000 14.220000 40.200000 ;
        RECT 13.950000 48.215000 14.250000 48.285000 ;
        RECT 13.990000 40.060000 14.290000 40.130000 ;
        RECT 14.020000 48.285000 14.320000 48.355000 ;
        RECT 14.060000 39.990000 14.360000 40.060000 ;
        RECT 14.090000 48.355000 14.390000 48.425000 ;
        RECT 14.130000 39.920000 14.430000 39.990000 ;
        RECT 14.160000 48.425000 14.460000 48.495000 ;
        RECT 14.180000 39.870000 15.420000 39.920000 ;
        RECT 14.195000 58.050000 14.835000 58.310000 ;
        RECT 14.210000 58.035000 14.820000 58.050000 ;
        RECT 14.230000 48.495000 14.530000 48.565000 ;
        RECT 14.240000 48.565000 14.600000 48.575000 ;
        RECT 14.250000 39.800000 15.470000 39.870000 ;
        RECT 14.280000 57.965000 14.750000 58.035000 ;
        RECT 14.295000 48.575000 14.610000 48.630000 ;
        RECT 14.320000 39.730000 15.540000 39.800000 ;
        RECT 14.350000 48.630000 14.610000 48.685000 ;
        RECT 14.350000 48.685000 14.610000 57.825000 ;
        RECT 14.350000 57.825000 14.610000 57.860000 ;
        RECT 14.350000 57.860000 14.645000 57.895000 ;
        RECT 14.350000 57.895000 14.680000 57.965000 ;
        RECT 14.390000 39.660000 15.610000 39.730000 ;
        RECT 15.365000 39.605000 15.680000 39.660000 ;
        RECT 15.435000 39.535000 15.735000 39.605000 ;
        RECT 15.505000 39.465000 15.805000 39.535000 ;
        RECT 15.575000 39.395000 15.875000 39.465000 ;
        RECT 15.645000 39.325000 15.945000 39.395000 ;
        RECT 15.715000 39.255000 16.015000 39.325000 ;
        RECT 15.785000 39.185000 16.085000 39.255000 ;
        RECT 15.855000 39.115000 16.155000 39.185000 ;
        RECT 15.925000 39.045000 16.225000 39.115000 ;
        RECT 15.995000 38.975000 16.295000 39.045000 ;
        RECT 16.065000 38.905000 16.365000 38.975000 ;
        RECT 16.135000 38.835000 16.435000 38.905000 ;
        RECT 16.205000 38.765000 16.505000 38.835000 ;
        RECT 16.275000 38.695000 16.575000 38.765000 ;
        RECT 16.310000  0.000000 16.570000  2.210000 ;
        RECT 16.310000  2.210000 16.570000  2.265000 ;
        RECT 16.310000  2.265000 16.625000  2.320000 ;
        RECT 16.345000 38.625000 16.645000 38.695000 ;
        RECT 16.365000 31.560000 16.680000 31.615000 ;
        RECT 16.365000 31.615000 16.625000 31.670000 ;
        RECT 16.365000 31.670000 16.625000 34.210000 ;
        RECT 16.365000 34.210000 16.625000 34.265000 ;
        RECT 16.365000 34.265000 16.680000 34.320000 ;
        RECT 16.370000 31.555000 16.735000 31.560000 ;
        RECT 16.380000  2.320000 16.680000  2.390000 ;
        RECT 16.415000 38.555000 16.715000 38.625000 ;
        RECT 16.435000 31.490000 16.740000 31.555000 ;
        RECT 16.435000 34.320000 16.735000 34.390000 ;
        RECT 16.450000  2.390000 16.750000  2.460000 ;
        RECT 16.485000 38.485000 16.785000 38.555000 ;
        RECT 16.500000 31.425000 16.805000 31.490000 ;
        RECT 16.505000 34.390000 16.805000 34.460000 ;
        RECT 16.520000  2.460000 16.820000  2.530000 ;
        RECT 16.555000 31.370000 16.870000 31.425000 ;
        RECT 16.555000 38.415000 16.855000 38.485000 ;
        RECT 16.575000 34.460000 16.875000 34.530000 ;
        RECT 16.590000  2.530000 16.890000  2.600000 ;
        RECT 16.610000  7.160000 16.925000  7.215000 ;
        RECT 16.610000  7.215000 16.870000  7.270000 ;
        RECT 16.610000  7.270000 16.870000 11.540000 ;
        RECT 16.610000 12.475000 16.870000 31.315000 ;
        RECT 16.610000 31.315000 16.870000 31.370000 ;
        RECT 16.615000 12.470000 16.870000 12.475000 ;
        RECT 16.625000 38.345000 16.925000 38.415000 ;
        RECT 16.635000  7.135000 16.980000  7.160000 ;
        RECT 16.645000 34.530000 16.945000 34.600000 ;
        RECT 16.655000 11.540000 16.870000 11.585000 ;
        RECT 16.660000  2.600000 16.960000  2.670000 ;
        RECT 16.660000 12.425000 16.870000 12.470000 ;
        RECT 16.695000 38.275000 16.995000 38.345000 ;
        RECT 16.700000 11.585000 16.870000 11.630000 ;
        RECT 16.705000  7.065000 17.005000  7.135000 ;
        RECT 16.705000 11.630000 16.870000 11.635000 ;
        RECT 16.705000 11.635000 16.870000 12.380000 ;
        RECT 16.705000 12.380000 16.870000 12.425000 ;
        RECT 16.715000 34.600000 17.015000 34.670000 ;
        RECT 16.730000  2.670000 17.030000  2.740000 ;
        RECT 16.765000 38.205000 17.065000 38.275000 ;
        RECT 16.775000  6.995000 17.075000  7.065000 ;
        RECT 16.785000 34.670000 17.085000 34.740000 ;
        RECT 16.800000  2.740000 17.100000  2.810000 ;
        RECT 16.835000 38.135000 17.135000 38.205000 ;
        RECT 16.845000  6.925000 17.145000  6.995000 ;
        RECT 16.855000 34.740000 17.155000 34.810000 ;
        RECT 16.870000  2.810000 17.170000  2.880000 ;
        RECT 16.905000 38.065000 17.205000 38.135000 ;
        RECT 16.915000  6.855000 17.215000  6.925000 ;
        RECT 16.925000 34.810000 17.225000 34.880000 ;
        RECT 16.940000  2.880000 17.240000  2.950000 ;
        RECT 16.975000 37.995000 17.275000 38.065000 ;
        RECT 16.985000  2.950000 17.310000  2.995000 ;
        RECT 16.985000  6.785000 17.285000  6.855000 ;
        RECT 16.995000 34.880000 17.295000 34.950000 ;
        RECT 17.040000  2.995000 17.355000  3.050000 ;
        RECT 17.040000  6.730000 17.355000  6.785000 ;
        RECT 17.045000 37.925000 17.345000 37.995000 ;
        RECT 17.065000 34.950000 17.365000 35.020000 ;
        RECT 17.095000  3.050000 17.355000  3.105000 ;
        RECT 17.095000  3.105000 17.355000  6.675000 ;
        RECT 17.095000  6.675000 17.355000  6.730000 ;
        RECT 17.115000 37.855000 17.415000 37.925000 ;
        RECT 17.135000 35.020000 17.435000 35.090000 ;
        RECT 17.185000 37.785000 17.485000 37.855000 ;
        RECT 17.205000 35.090000 17.505000 35.160000 ;
        RECT 17.255000 37.715000 17.555000 37.785000 ;
        RECT 17.275000 35.160000 17.575000 35.230000 ;
        RECT 17.325000 37.645000 17.625000 37.715000 ;
        RECT 17.345000 35.230000 17.645000 35.300000 ;
        RECT 17.395000 37.575000 17.695000 37.645000 ;
        RECT 17.415000 35.300000 17.715000 35.370000 ;
        RECT 17.465000 35.370000 17.785000 35.420000 ;
        RECT 17.465000 37.505000 17.765000 37.575000 ;
        RECT 17.520000 35.420000 17.835000 35.475000 ;
        RECT 17.520000 37.450000 17.835000 37.505000 ;
        RECT 17.575000 35.475000 17.835000 35.530000 ;
        RECT 17.575000 35.530000 17.835000 37.395000 ;
        RECT 17.575000 37.395000 17.835000 37.450000 ;
    END
  END ENABLE_VSWITCH_H
  PIN HLD_H_N
    ANTENNAGATEAREA  1.620000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.815000 0.000000 32.075000 3.965000 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.600000 0.000000 26.860000 1.695000 ;
    END
  END HLD_OVR
  PIN IB_MODE_SEL
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.420000 0.000000 5.650000 4.375000 ;
        RECT 5.420000 4.375000 5.650000 4.425000 ;
        RECT 5.420000 4.425000 5.700000 4.475000 ;
        RECT 5.490000 4.475000 5.750000 4.545000 ;
        RECT 5.560000 4.545000 5.820000 4.615000 ;
        RECT 5.630000 4.615000 5.890000 4.685000 ;
        RECT 5.700000 4.685000 5.960000 4.755000 ;
        RECT 5.770000 4.755000 6.030000 4.825000 ;
        RECT 5.840000 4.825000 6.100000 4.895000 ;
        RECT 5.910000 4.895000 6.170000 4.965000 ;
        RECT 5.910000 6.425000 6.550000 6.685000 ;
        RECT 5.980000 4.965000 6.240000 5.035000 ;
        RECT 6.050000 5.035000 6.310000 5.105000 ;
        RECT 6.120000 5.105000 6.380000 5.175000 ;
        RECT 6.180000 6.390000 6.550000 6.425000 ;
        RECT 6.190000 5.175000 6.450000 5.245000 ;
        RECT 6.220000 5.245000 6.520000 5.275000 ;
        RECT 6.250000 6.320000 6.550000 6.390000 ;
        RECT 6.270000 5.275000 6.550000 5.325000 ;
        RECT 6.320000 5.325000 6.550000 5.375000 ;
        RECT 6.320000 5.375000 6.550000 6.250000 ;
        RECT 6.320000 6.250000 6.550000 6.320000 ;
    END
  END IB_MODE_SEL
  PIN IN
    ANTENNAPARTIALMETALSIDEAREA  303.1200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.240000 0.000000 79.570000 176.480000 ;
    END
  END IN
  PIN INP_DIS
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.245000 0.000000 45.505000 4.980000 ;
        RECT 45.245000 4.980000 45.505000 5.035000 ;
        RECT 45.245000 5.035000 45.560000 5.090000 ;
        RECT 45.315000 5.090000 45.615000 5.160000 ;
        RECT 45.385000 5.160000 45.685000 5.230000 ;
        RECT 45.455000 5.230000 45.755000 5.300000 ;
        RECT 45.525000 5.300000 45.825000 5.370000 ;
        RECT 45.595000 5.370000 45.895000 5.440000 ;
        RECT 45.665000 5.440000 45.965000 5.510000 ;
        RECT 45.735000 5.510000 46.035000 5.580000 ;
        RECT 45.745000 5.580000 46.105000 5.590000 ;
        RECT 45.800000 5.590000 46.115000 5.645000 ;
        RECT 45.855000 5.645000 46.115000 5.700000 ;
        RECT 45.855000 5.700000 46.115000 6.780000 ;
    END
  END INP_DIS
  PIN IN_H
    ANTENNAPARTIALMETALSIDEAREA  291.9480 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.400000   0.000000 1.020000 178.235000 ;
        RECT 0.400000 178.235000 1.020000 178.360000 ;
        RECT 0.400000 178.360000 1.145000 178.485000 ;
        RECT 0.550000 178.485000 1.270000 178.635000 ;
        RECT 0.700000 178.635000 1.420000 178.785000 ;
        RECT 0.850000 178.785000 1.570000 178.935000 ;
        RECT 1.000000 178.935000 1.720000 179.085000 ;
        RECT 1.150000 179.085000 1.870000 179.235000 ;
        RECT 1.300000 179.235000 2.020000 179.385000 ;
        RECT 1.450000 179.385000 2.170000 179.535000 ;
        RECT 1.600000 179.535000 2.320000 179.685000 ;
        RECT 1.750000 179.685000 2.470000 179.835000 ;
        RECT 1.900000 179.835000 2.620000 179.985000 ;
        RECT 2.050000 179.985000 2.770000 180.135000 ;
        RECT 2.200000 180.135000 2.920000 180.285000 ;
        RECT 2.350000 180.285000 3.070000 180.435000 ;
        RECT 2.355000 180.435000 3.220000 180.440000 ;
        RECT 2.505000 180.440000 4.565000 180.590000 ;
        RECT 2.655000 180.590000 4.565000 180.740000 ;
        RECT 2.805000 180.740000 4.565000 180.890000 ;
        RECT 2.955000 180.890000 4.565000 181.040000 ;
        RECT 3.085000 181.040000 4.565000 181.170000 ;
    END
  END IN_H
  PIN OE_N
    ANTENNAGATEAREA  1.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.375000  0.000000 3.605000  4.375000 ;
        RECT 3.375000  4.375000 3.605000  4.425000 ;
        RECT 3.375000  4.425000 3.655000  4.475000 ;
        RECT 3.445000  4.475000 3.705000  4.545000 ;
        RECT 3.515000  4.545000 3.775000  4.615000 ;
        RECT 3.585000  4.615000 3.845000  4.685000 ;
        RECT 3.655000  4.685000 3.915000  4.755000 ;
        RECT 3.725000  4.755000 3.985000  4.825000 ;
        RECT 3.770000  4.825000 4.055000  4.870000 ;
        RECT 3.840000  4.870000 5.225000  4.940000 ;
        RECT 3.910000  4.940000 5.295000  5.010000 ;
        RECT 3.980000  5.010000 5.365000  5.080000 ;
        RECT 4.000000  5.080000 5.435000  5.100000 ;
        RECT 5.195000  5.100000 5.455000  5.170000 ;
        RECT 5.265000  5.170000 5.525000  5.240000 ;
        RECT 5.300000  5.240000 5.595000  5.275000 ;
        RECT 5.350000  5.275000 5.630000  5.325000 ;
        RECT 5.400000  5.325000 5.630000  5.375000 ;
        RECT 5.400000  5.375000 5.630000  8.250000 ;
        RECT 5.400000  8.250000 5.630000  8.300000 ;
        RECT 5.400000  8.300000 5.680000  8.350000 ;
        RECT 5.470000  8.350000 5.730000  8.420000 ;
        RECT 5.540000  8.420000 5.800000  8.490000 ;
        RECT 5.610000  8.490000 5.870000  8.560000 ;
        RECT 5.680000  8.560000 5.940000  8.630000 ;
        RECT 5.750000  8.630000 6.010000  8.700000 ;
        RECT 5.820000  8.700000 6.080000  8.770000 ;
        RECT 5.890000  8.770000 6.150000  8.840000 ;
        RECT 5.960000  8.840000 6.220000  8.910000 ;
        RECT 5.965000 42.985000 6.225000 43.625000 ;
        RECT 5.970000 42.980000 6.220000 42.985000 ;
        RECT 5.975000 39.420000 6.255000 39.470000 ;
        RECT 5.975000 39.470000 6.205000 39.520000 ;
        RECT 5.975000 39.520000 6.205000 42.965000 ;
        RECT 5.975000 42.965000 6.205000 42.970000 ;
        RECT 5.975000 42.970000 6.210000 42.975000 ;
        RECT 5.975000 42.975000 6.215000 42.980000 ;
        RECT 5.985000 39.410000 6.305000 39.420000 ;
        RECT 6.030000  8.910000 6.290000  8.980000 ;
        RECT 6.055000 39.340000 6.315000 39.410000 ;
        RECT 6.100000  8.980000 6.360000  9.050000 ;
        RECT 6.125000 39.270000 6.385000 39.340000 ;
        RECT 6.170000  9.050000 6.430000  9.120000 ;
        RECT 6.195000 39.200000 6.455000 39.270000 ;
        RECT 6.240000  9.120000 6.500000  9.190000 ;
        RECT 6.265000 39.130000 6.525000 39.200000 ;
        RECT 6.310000  9.190000 6.570000  9.260000 ;
        RECT 6.335000 39.060000 6.595000 39.130000 ;
        RECT 6.380000  9.260000 6.640000  9.330000 ;
        RECT 6.405000 38.990000 6.665000 39.060000 ;
        RECT 6.450000  9.330000 6.710000  9.400000 ;
        RECT 6.475000  9.400000 6.780000  9.425000 ;
        RECT 6.475000 38.920000 6.735000 38.990000 ;
        RECT 6.525000  9.425000 6.805000  9.475000 ;
        RECT 6.525000 38.870000 6.805000 38.920000 ;
        RECT 6.575000  9.475000 6.805000  9.525000 ;
        RECT 6.575000  9.525000 6.805000 38.820000 ;
        RECT 6.575000 38.820000 6.805000 38.870000 ;
    END
  END OE_N
  PIN OUT
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.355000  0.000000 22.615000  6.315000 ;
        RECT 22.355000  6.315000 22.615000  6.370000 ;
        RECT 22.355000  6.370000 22.670000  6.425000 ;
        RECT 22.425000  6.425000 22.725000  6.495000 ;
        RECT 22.495000  6.495000 22.795000  6.565000 ;
        RECT 22.565000  6.565000 22.865000  6.635000 ;
        RECT 22.635000  6.635000 22.935000  6.705000 ;
        RECT 22.655000  6.705000 23.005000  6.725000 ;
        RECT 22.710000  6.725000 23.025000  6.780000 ;
        RECT 22.765000  6.780000 23.025000  6.835000 ;
        RECT 22.765000  6.835000 23.025000 14.375000 ;
        RECT 22.765000 14.375000 23.025000 14.430000 ;
        RECT 22.765000 14.430000 23.080000 14.485000 ;
        RECT 22.835000 14.485000 23.135000 14.555000 ;
        RECT 22.905000 14.555000 23.205000 14.625000 ;
        RECT 22.975000 14.625000 23.275000 14.695000 ;
        RECT 23.045000 14.695000 23.345000 14.765000 ;
        RECT 23.095000 38.695000 23.735000 38.955000 ;
        RECT 23.115000 14.765000 23.415000 14.835000 ;
        RECT 23.185000 14.835000 23.485000 14.905000 ;
        RECT 23.255000 14.905000 23.555000 14.975000 ;
        RECT 23.265000 38.625000 23.735000 38.695000 ;
        RECT 23.325000 14.975000 23.625000 15.045000 ;
        RECT 23.335000 38.555000 23.735000 38.625000 ;
        RECT 23.395000 15.045000 23.695000 15.115000 ;
        RECT 23.405000 38.485000 23.735000 38.555000 ;
        RECT 23.465000 15.115000 23.765000 15.185000 ;
        RECT 23.475000 25.180000 23.790000 25.235000 ;
        RECT 23.475000 25.235000 23.735000 25.290000 ;
        RECT 23.475000 25.290000 23.735000 38.415000 ;
        RECT 23.475000 38.415000 23.735000 38.485000 ;
        RECT 23.510000 25.145000 23.845000 25.180000 ;
        RECT 23.535000 15.185000 23.835000 15.255000 ;
        RECT 23.545000 15.255000 23.905000 15.265000 ;
        RECT 23.545000 25.110000 23.880000 25.145000 ;
        RECT 23.600000 15.265000 23.915000 15.320000 ;
        RECT 23.600000 25.055000 23.915000 25.110000 ;
        RECT 23.655000 15.320000 23.915000 15.375000 ;
        RECT 23.655000 15.375000 23.915000 25.000000 ;
        RECT 23.655000 25.000000 23.915000 25.055000 ;
    END
  END OUT
  PIN PAD
    ANTENNAPARTIALMETALSIDEAREA  216.1550 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.115000 125.470000 53.655000 147.015000 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    ANTENNAPARTIALMETALSIDEAREA  3.812250 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.280000 0.000000 76.920000 1.625000 ;
        RECT 76.280000 1.625000 76.920000 1.695000 ;
        RECT 76.280000 1.695000 76.990000 1.765000 ;
        RECT 76.280000 1.765000 77.060000 1.835000 ;
        RECT 76.280000 1.835000 77.130000 1.905000 ;
        RECT 76.280000 1.905000 77.200000 1.975000 ;
        RECT 76.280000 1.975000 77.270000 2.045000 ;
        RECT 76.280000 2.045000 77.340000 2.055000 ;
        RECT 76.350000 2.055000 77.350000 2.125000 ;
        RECT 76.420000 2.125000 77.420000 2.195000 ;
        RECT 76.490000 2.195000 77.490000 2.265000 ;
        RECT 76.560000 2.265000 77.560000 2.335000 ;
        RECT 76.630000 2.335000 77.630000 2.405000 ;
        RECT 76.700000 2.405000 77.700000 2.475000 ;
        RECT 76.770000 2.475000 77.770000 2.545000 ;
        RECT 76.820000 2.545000 77.840000 2.595000 ;
        RECT 76.890000 2.595000 77.890000 2.665000 ;
        RECT 76.960000 2.665000 77.890000 2.735000 ;
        RECT 77.030000 2.735000 77.890000 2.805000 ;
        RECT 77.100000 2.805000 77.890000 2.875000 ;
        RECT 77.150000 2.875000 77.890000 2.925000 ;
        RECT 77.150000 2.925000 77.890000 5.235000 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    ANTENNAPARTIALMETALSIDEAREA  2.618000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.275000 0.000000 68.925000 3.960000 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    ANTENNAPARTIALCUTAREA  4.960000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.600000  7.425000 60.560000   7.575000 ;
        RECT 59.600000  7.575000 60.410000   7.725000 ;
        RECT 59.600000  7.725000 60.385000   7.750000 ;
        RECT 59.600000  7.750000 60.385000  10.610000 ;
        RECT 59.600000 10.610000 60.385000  10.760000 ;
        RECT 59.600000 10.760000 60.535000  10.910000 ;
        RECT 59.600000 10.910000 60.685000  10.935000 ;
        RECT 59.655000  7.370000 60.710000   7.425000 ;
        RECT 59.750000 10.935000 60.710000  11.085000 ;
        RECT 59.805000  7.220000 60.765000   7.370000 ;
        RECT 59.900000 11.085000 60.860000  11.235000 ;
        RECT 59.955000  7.070000 60.915000   7.220000 ;
        RECT 59.985000  7.040000 63.890000   7.070000 ;
        RECT 60.050000 11.235000 61.010000  11.385000 ;
        RECT 60.135000  6.890000 63.890000   7.040000 ;
        RECT 60.200000 11.385000 61.160000  11.535000 ;
        RECT 60.285000  6.740000 63.890000   6.890000 ;
        RECT 60.350000 11.535000 61.310000  11.685000 ;
        RECT 60.435000  6.590000 63.890000   6.740000 ;
        RECT 60.500000 11.685000 61.460000  11.835000 ;
        RECT 60.585000  6.440000 63.890000   6.590000 ;
        RECT 60.610000 19.065000 61.570000  19.215000 ;
        RECT 60.610000 19.215000 61.420000  19.365000 ;
        RECT 60.610000 19.365000 61.395000  19.390000 ;
        RECT 60.610000 19.390000 61.395000  47.360000 ;
        RECT 60.650000 11.835000 61.610000  11.985000 ;
        RECT 60.690000 18.985000 61.720000  19.065000 ;
        RECT 60.735000  6.290000 63.890000   6.440000 ;
        RECT 60.800000 11.985000 61.760000  12.135000 ;
        RECT 60.840000 18.835000 61.800000  18.985000 ;
        RECT 60.950000 12.135000 61.910000  12.285000 ;
        RECT 60.990000 18.685000 61.950000  18.835000 ;
        RECT 61.100000 12.285000 62.060000  12.435000 ;
        RECT 61.140000 12.435000 62.210000  12.475000 ;
        RECT 61.140000 18.535000 62.100000  18.685000 ;
        RECT 61.170000 18.505000 62.250000  18.535000 ;
        RECT 61.290000 12.475000 62.250000  12.625000 ;
        RECT 61.320000 18.355000 62.250000  18.505000 ;
        RECT 61.440000 12.625000 62.250000  12.775000 ;
        RECT 61.470000 12.775000 62.250000  12.805000 ;
        RECT 61.470000 12.805000 62.250000  18.205000 ;
        RECT 61.470000 18.205000 62.250000  18.355000 ;
        RECT 61.710000 35.760000 63.070000  35.910000 ;
        RECT 61.710000 35.910000 62.920000  36.060000 ;
        RECT 61.710000 36.060000 62.780000  36.200000 ;
        RECT 61.710000 36.200000 62.780000  73.005000 ;
        RECT 61.710000 73.005000 62.780000  73.155000 ;
        RECT 61.710000 73.155000 62.930000  73.305000 ;
        RECT 61.710000 73.305000 63.080000  73.455000 ;
        RECT 61.710000 73.455000 63.230000  73.605000 ;
        RECT 61.710000 73.605000 63.380000  73.755000 ;
        RECT 61.710000 73.755000 63.530000  73.905000 ;
        RECT 61.710000 73.905000 63.680000  74.055000 ;
        RECT 61.710000 74.055000 63.830000  74.185000 ;
        RECT 61.735000 35.735000 63.220000  35.760000 ;
        RECT 61.750000 74.185000 63.960000  74.225000 ;
        RECT 61.790000 74.225000 64.000000  74.265000 ;
        RECT 61.885000 35.585000 63.245000  35.735000 ;
        RECT 61.940000 74.265000 68.555000  74.415000 ;
        RECT 62.035000 35.435000 63.395000  35.585000 ;
        RECT 62.090000 74.415000 68.705000  74.565000 ;
        RECT 62.185000 35.285000 63.545000  35.435000 ;
        RECT 62.220000  6.155000 63.890000   6.290000 ;
        RECT 62.235000  7.070000 63.890000   7.220000 ;
        RECT 62.240000 74.565000 68.855000  74.715000 ;
        RECT 62.325000 35.145000 63.695000  35.285000 ;
        RECT 62.370000  6.005000 63.890000   6.155000 ;
        RECT 62.385000  7.220000 63.890000   7.370000 ;
        RECT 62.390000 74.715000 69.005000  74.865000 ;
        RECT 62.475000 34.995000 63.695000  35.145000 ;
        RECT 62.520000  5.855000 63.890000   6.005000 ;
        RECT 62.535000  7.370000 63.890000   7.520000 ;
        RECT 62.540000 74.865000 69.155000  75.015000 ;
        RECT 62.625000 17.825000 63.890000  18.070000 ;
        RECT 62.625000 18.070000 63.795000  18.165000 ;
        RECT 62.625000 18.165000 63.700000  18.260000 ;
        RECT 62.625000 18.260000 63.695000  18.265000 ;
        RECT 62.625000 18.265000 63.695000  34.845000 ;
        RECT 62.625000 34.845000 63.695000  34.995000 ;
        RECT 62.630000 17.820000 63.890000  17.825000 ;
        RECT 62.670000  5.705000 63.890000   5.855000 ;
        RECT 62.685000  7.520000 63.890000   7.670000 ;
        RECT 62.690000 75.015000 69.305000  75.165000 ;
        RECT 62.725000 17.725000 63.890000  17.820000 ;
        RECT 62.820000  0.000000 63.890000   5.555000 ;
        RECT 62.820000  5.555000 63.890000   5.705000 ;
        RECT 62.820000  7.670000 63.890000   7.805000 ;
        RECT 62.820000  7.805000 63.890000  17.630000 ;
        RECT 62.820000 17.630000 63.890000  17.725000 ;
        RECT 62.840000 75.165000 69.455000  75.315000 ;
        RECT 62.860000 75.315000 69.605000  75.335000 ;
        RECT 67.870000 75.335000 69.625000  75.400000 ;
        RECT 67.935000 75.400000 69.690000  75.465000 ;
        RECT 67.940000 75.465000 69.755000  75.470000 ;
        RECT 68.090000 75.470000 69.760000  75.620000 ;
        RECT 68.240000 75.620000 69.760000  75.770000 ;
        RECT 68.390000 75.770000 69.760000  75.920000 ;
        RECT 68.540000 75.920000 69.760000  76.070000 ;
        RECT 68.690000 76.070000 69.760000  76.220000 ;
        RECT 68.690000 76.220000 69.760000 101.910000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.000000 106.585000 12.500000 118.955000 ;
        RECT 7.665000 118.955000 12.500000 119.105000 ;
        RECT 7.815000 119.105000 12.500000 119.255000 ;
        RECT 7.850000 106.565000 12.500000 106.585000 ;
        RECT 7.965000 119.255000 12.500000 119.405000 ;
        RECT 8.000000 106.415000 12.500000 106.565000 ;
        RECT 8.115000 119.405000 12.500000 119.555000 ;
        RECT 8.150000 106.265000 12.500000 106.415000 ;
        RECT 8.265000 119.555000 12.500000 119.705000 ;
        RECT 8.300000 106.115000 12.500000 106.265000 ;
        RECT 8.415000 119.705000 12.500000 119.855000 ;
        RECT 8.450000 105.965000 12.500000 106.115000 ;
        RECT 8.565000 119.855000 12.500000 120.005000 ;
        RECT 8.600000 105.815000 12.500000 105.965000 ;
        RECT 8.715000 120.005000 12.500000 120.155000 ;
        RECT 8.750000 105.665000 12.500000 105.815000 ;
        RECT 8.865000 120.155000 12.500000 120.305000 ;
        RECT 8.900000 105.515000 12.500000 105.665000 ;
        RECT 9.015000 120.305000 12.500000 120.455000 ;
        RECT 9.050000 105.365000 12.500000 105.515000 ;
        RECT 9.165000 120.455000 12.500000 120.605000 ;
        RECT 9.200000 105.215000 12.500000 105.365000 ;
        RECT 9.315000 120.605000 12.500000 120.755000 ;
        RECT 9.350000 105.065000 12.500000 105.215000 ;
        RECT 9.465000 120.755000 12.500000 120.905000 ;
        RECT 9.500000 104.915000 12.500000 105.065000 ;
        RECT 9.615000 120.905000 12.500000 121.055000 ;
        RECT 9.650000 104.765000 12.500000 104.915000 ;
        RECT 9.765000 121.055000 12.500000 121.205000 ;
        RECT 9.800000 104.615000 12.500000 104.765000 ;
        RECT 9.810000 121.205000 12.500000 121.250000 ;
    END
  END PAD_A_NOESD_H
  PIN SLOW
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.390000 1.185000 78.210000 1.465000 ;
        RECT 77.470000 1.125000 78.120000 1.185000 ;
        RECT 77.540000 1.055000 78.050000 1.125000 ;
        RECT 77.610000 0.000000 77.870000 0.875000 ;
        RECT 77.610000 0.875000 77.870000 0.930000 ;
        RECT 77.610000 0.930000 77.925000 0.985000 ;
        RECT 77.610000 0.985000 77.980000 1.055000 ;
    END
  END SLOW
  PIN TIE_HI_ESD
    ANTENNAPARTIALMETALSIDEAREA  85.19250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.230000 50.760000 76.475000 50.805000 ;
        RECT 76.230000 50.805000 76.430000 50.850000 ;
        RECT 76.230000 50.850000 76.430000 52.425000 ;
        RECT 76.230000 52.425000 76.430000 52.470000 ;
        RECT 76.230000 52.470000 76.475000 52.515000 ;
        RECT 76.280000 50.710000 76.520000 50.760000 ;
        RECT 76.300000 52.515000 76.520000 52.585000 ;
        RECT 76.350000 50.640000 76.570000 50.710000 ;
        RECT 76.370000 52.585000 76.590000 52.655000 ;
        RECT 76.420000 50.570000 76.640000 50.640000 ;
        RECT 76.440000 52.655000 76.660000 52.725000 ;
        RECT 76.490000 50.500000 76.710000 50.570000 ;
        RECT 76.510000 52.725000 76.730000 52.795000 ;
        RECT 76.560000 50.430000 76.780000 50.500000 ;
        RECT 76.580000 52.795000 76.800000 52.865000 ;
        RECT 76.630000 50.360000 76.850000 50.430000 ;
        RECT 76.650000 52.865000 76.870000 52.935000 ;
        RECT 76.700000 50.290000 76.920000 50.360000 ;
        RECT 76.720000 52.935000 76.940000 53.005000 ;
        RECT 76.770000 50.220000 76.990000 50.290000 ;
        RECT 76.790000 53.005000 77.010000 53.075000 ;
        RECT 76.825000 53.075000 77.080000 53.110000 ;
        RECT 76.840000 50.150000 77.060000 50.220000 ;
        RECT 76.870000 53.110000 77.115000 53.155000 ;
        RECT 76.900000 96.210000 77.130000 96.225000 ;
        RECT 76.910000 50.080000 77.130000 50.150000 ;
        RECT 76.915000 53.155000 77.115000 53.200000 ;
        RECT 76.915000 53.200000 77.115000 96.195000 ;
        RECT 76.915000 96.195000 77.115000 96.210000 ;
        RECT 76.980000 50.010000 77.200000 50.080000 ;
        RECT 77.050000 49.940000 77.270000 50.010000 ;
        RECT 77.120000 49.870000 77.340000 49.940000 ;
        RECT 77.190000 49.800000 77.410000 49.870000 ;
        RECT 77.260000 49.730000 77.480000 49.800000 ;
        RECT 77.330000 49.660000 77.550000 49.730000 ;
        RECT 77.400000 49.590000 77.620000 49.660000 ;
        RECT 77.470000 49.520000 77.690000 49.590000 ;
        RECT 77.540000 49.450000 77.760000 49.520000 ;
        RECT 77.610000 49.380000 77.830000 49.450000 ;
        RECT 77.680000 49.310000 77.900000 49.380000 ;
        RECT 77.750000 49.240000 77.970000 49.310000 ;
        RECT 77.820000 49.170000 78.040000 49.240000 ;
        RECT 77.890000 49.100000 78.110000 49.170000 ;
        RECT 77.960000 49.030000 78.180000 49.100000 ;
        RECT 78.030000 48.960000 78.250000 49.030000 ;
        RECT 78.100000 48.890000 78.320000 48.960000 ;
        RECT 78.170000 48.820000 78.390000 48.890000 ;
        RECT 78.240000 48.750000 78.460000 48.820000 ;
        RECT 78.310000 48.680000 78.530000 48.750000 ;
        RECT 78.380000 48.610000 78.600000 48.680000 ;
        RECT 78.450000 48.540000 78.670000 48.610000 ;
        RECT 78.520000 48.470000 78.740000 48.540000 ;
        RECT 78.590000 48.400000 78.810000 48.470000 ;
        RECT 78.615000 10.265000 78.910000 10.340000 ;
        RECT 78.615000 10.340000 78.860000 10.390000 ;
        RECT 78.615000 10.390000 78.810000 10.440000 ;
        RECT 78.615000 10.440000 78.805000 10.445000 ;
        RECT 78.615000 10.445000 78.805000 16.245000 ;
        RECT 78.615000 16.245000 78.805000 16.285000 ;
        RECT 78.615000 16.285000 78.845000 16.325000 ;
        RECT 78.620000 10.260000 78.910000 10.265000 ;
        RECT 78.660000 48.330000 78.880000 48.400000 ;
        RECT 78.665000 10.215000 78.910000 10.260000 ;
        RECT 78.685000 16.325000 78.885000 16.395000 ;
        RECT 78.705000  0.000000 78.905000  1.125000 ;
        RECT 78.705000  1.125000 78.905000  1.130000 ;
        RECT 78.705000  1.130000 78.910000  1.215000 ;
        RECT 78.710000  1.215000 78.910000  1.220000 ;
        RECT 78.710000  1.220000 78.910000 10.170000 ;
        RECT 78.710000 10.170000 78.910000 10.215000 ;
        RECT 78.730000 48.260000 78.950000 48.330000 ;
        RECT 78.755000 16.395000 78.955000 16.465000 ;
        RECT 78.800000 48.190000 79.020000 48.260000 ;
        RECT 78.825000 16.465000 79.025000 16.535000 ;
        RECT 78.870000 48.120000 79.090000 48.190000 ;
        RECT 78.895000 16.535000 79.095000 16.605000 ;
        RECT 78.940000 48.050000 79.160000 48.120000 ;
        RECT 78.965000 16.605000 79.165000 16.675000 ;
        RECT 79.010000 47.980000 79.230000 48.050000 ;
        RECT 79.035000 16.675000 79.235000 16.745000 ;
        RECT 79.080000 47.910000 79.300000 47.980000 ;
        RECT 79.105000 16.745000 79.305000 16.815000 ;
        RECT 79.150000 47.840000 79.370000 47.910000 ;
        RECT 79.175000 16.815000 79.375000 16.885000 ;
        RECT 79.220000 47.770000 79.440000 47.840000 ;
        RECT 79.240000 16.885000 79.445000 16.950000 ;
        RECT 79.270000 47.720000 79.510000 47.770000 ;
        RECT 79.280000 16.950000 79.510000 16.990000 ;
        RECT 79.320000 16.990000 79.510000 17.030000 ;
        RECT 79.320000 17.030000 79.510000 47.670000 ;
        RECT 79.320000 47.670000 79.510000 47.720000 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    ANTENNAPARTIALMETALSIDEAREA  165.2660 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.715000 0.000000 79.915000 96.000000 ;
    END
  END TIE_LO_ESD
  PIN VTRIP_SEL
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.130000 0.000000 6.390000 1.440000 ;
        RECT 6.130000 1.440000 6.390000 1.495000 ;
        RECT 6.130000 1.495000 6.445000 1.550000 ;
        RECT 6.200000 1.550000 6.500000 1.620000 ;
        RECT 6.270000 1.620000 6.570000 1.690000 ;
        RECT 6.340000 1.690000 6.640000 1.760000 ;
        RECT 6.410000 1.760000 6.710000 1.830000 ;
        RECT 6.480000 1.830000 6.780000 1.900000 ;
        RECT 6.550000 1.900000 6.850000 1.970000 ;
        RECT 6.620000 1.970000 6.920000 2.040000 ;
        RECT 6.690000 2.040000 6.990000 2.110000 ;
        RECT 6.760000 2.110000 7.060000 2.180000 ;
        RECT 6.830000 2.180000 7.130000 2.250000 ;
        RECT 6.900000 2.250000 7.200000 2.320000 ;
        RECT 6.970000 2.320000 7.270000 2.390000 ;
        RECT 7.040000 2.390000 7.340000 2.460000 ;
        RECT 7.110000 2.460000 7.410000 2.530000 ;
        RECT 7.180000 2.530000 7.480000 2.600000 ;
        RECT 7.250000 2.600000 7.550000 2.670000 ;
        RECT 7.320000 2.670000 7.620000 2.740000 ;
        RECT 7.390000 2.740000 7.690000 2.810000 ;
        RECT 7.460000 2.810000 7.760000 2.880000 ;
        RECT 7.530000 2.880000 7.830000 2.950000 ;
        RECT 7.600000 2.950000 7.900000 3.020000 ;
        RECT 7.670000 3.020000 7.970000 3.090000 ;
        RECT 7.740000 3.090000 8.040000 3.160000 ;
        RECT 7.810000 3.160000 8.110000 3.230000 ;
        RECT 7.880000 3.230000 8.180000 3.300000 ;
        RECT 7.950000 3.300000 8.250000 3.370000 ;
        RECT 8.020000 3.370000 8.320000 3.440000 ;
        RECT 8.090000 3.440000 8.390000 3.510000 ;
        RECT 8.160000 3.510000 8.460000 3.580000 ;
        RECT 8.230000 3.580000 8.530000 3.650000 ;
        RECT 8.300000 3.650000 8.600000 3.720000 ;
        RECT 8.335000 3.720000 8.670000 3.755000 ;
        RECT 8.390000 3.755000 8.705000 3.810000 ;
        RECT 8.445000 3.810000 8.705000 3.865000 ;
        RECT 8.445000 3.865000 8.705000 6.780000 ;
    END
  END VTRIP_SEL
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 8.885000 80.000000 13.535000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 2.035000 80.000000 7.485000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.035000 14.935000 80.000000 18.385000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 19.785000 80.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 70.035000 80.000000 95.000000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 64.085000 80.000000 68.535000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 36.735000 80.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 47.735000 80.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 51.645000 80.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 56.405000 80.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 41.585000 80.000000 46.235000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 175.785000 80.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 25.835000 80.000000 30.485000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 58.235000 80.000000 62.685000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 31.885000 80.000000 35.335000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT -0.115000  95.895000 45.710000  95.955000 ;
      RECT -0.115000  95.955000  4.915000 130.220000 ;
      RECT -0.115000 131.275000  4.915000 140.050000 ;
      RECT -0.115000 140.050000  1.495000 140.150000 ;
      RECT -0.115000 145.155000  1.495000 145.210000 ;
      RECT -0.115000 145.210000  4.915000 170.090000 ;
      RECT -0.085000  93.065000  9.000000  95.255000 ;
      RECT -0.085000  95.255000 45.710000  95.895000 ;
      RECT -0.085000 130.220000  4.915000 130.225000 ;
      RECT -0.085000 130.995000  4.915000 131.275000 ;
      RECT -0.085000 170.090000  4.915000 178.645000 ;
      RECT  0.950000  18.885000  1.310000  19.055000 ;
      RECT  0.980000  21.465000  1.310000  21.635000 ;
      RECT  1.120000  22.325000  1.310000  22.495000 ;
      RECT  1.150000  19.745000  1.310000  19.915000 ;
      RECT  1.150000  20.605000  1.310000  20.775000 ;
      RECT  1.690000  45.545000  4.585000  45.715000 ;
      RECT  2.260000 145.155000  4.700000 145.210000 ;
      RECT  5.875000   5.940000  6.405000   6.465000 ;
      RECT  6.490000  88.950000  9.000000  93.065000 ;
      RECT  7.805000   5.400000 67.100000   6.230000 ;
      RECT  9.300000  32.000000  9.660000  36.750000 ;
      RECT 10.330000  32.000000 10.690000  36.750000 ;
      RECT 11.410000  32.000000 11.665000  37.260000 ;
      RECT 11.940000  31.110000 12.365000  36.765000 ;
      RECT 12.610000  32.000000 13.140000  37.260000 ;
      RECT 13.390000  32.000000 13.920000  36.750000 ;
      RECT 14.170000  32.000000 14.700000  36.750000 ;
      RECT 14.170000  36.750000 14.305000  37.260000 ;
      RECT 14.320000  26.760000 14.500000  29.470000 ;
      RECT 14.320000  29.470000 14.670000  29.570000 ;
      RECT 14.320000  29.570000 14.490000  30.110000 ;
      RECT 14.955000  32.000000 15.485000  37.260000 ;
      RECT 15.105000  26.760000 15.635000  29.690000 ;
      RECT 15.730000  32.000000 16.260000  36.750000 ;
      RECT 15.730000 179.435000 68.925000 179.450000 ;
      RECT 15.730000 179.450000 77.885000 179.980000 ;
      RECT 15.730000 179.980000 68.925000 180.205000 ;
      RECT 15.885000  26.760000 16.415000  29.470000 ;
      RECT 16.510000  32.000000 16.950000  37.260000 ;
      RECT 16.670000  26.760000 17.200000  29.690000 ;
      RECT 17.210000  32.000000 17.650000  36.750000 ;
      RECT 18.035000  26.760000 18.450000  29.470000 ;
      RECT 18.140000  32.060000 18.630000  36.750000 ;
      RECT 19.040000  26.760000 19.455000  29.470000 ;
      RECT 19.050000  32.000000 19.580000  36.750000 ;
      RECT 19.790000  26.760000 20.320000  29.470000 ;
      RECT 20.640000  32.000000 21.170000  36.750000 ;
      RECT 21.690000  26.760000 22.130000  29.470000 ;
      RECT 22.170000  32.000000 22.700000  36.755000 ;
      RECT 23.725000  32.000000 24.255000  36.755000 ;
      RECT 23.800000  26.760000 24.160000  29.470000 ;
      RECT 24.340000  25.580000 26.330000  25.905000 ;
      RECT 24.340000  25.905000 24.835000  29.690000 ;
      RECT 25.015000  26.760000 25.545000  29.470000 ;
      RECT 25.675000  32.250000 26.090000  37.000000 ;
      RECT 25.930000  59.095000 28.100000  60.125000 ;
      RECT 25.935000  57.585000 29.370000  58.865000 ;
      RECT 26.225000  19.595000 26.670000  24.375000 ;
      RECT 26.385000  32.250000 26.865000  37.330000 ;
      RECT 26.390000  26.760000 26.750000  29.690000 ;
      RECT 26.525000  67.105000 29.670000  67.815000 ;
      RECT 26.975000  19.600000 27.420000  24.365000 ;
      RECT 27.045000  32.250000 27.575000  37.000000 ;
      RECT 27.490000  63.970000 29.315000  64.550000 ;
      RECT 27.510000  26.490000 28.090000  30.360000 ;
      RECT 27.675000  68.735000 29.670000  69.445000 ;
      RECT 27.830000  32.245000 28.360000  37.330000 ;
      RECT 28.340000  59.180000 28.510000  59.710000 ;
      RECT 28.605000  32.250000 29.135000  37.005000 ;
      RECT 28.680000  18.995000 29.210000  23.750000 ;
      RECT 28.860000  95.125000 45.710000  95.255000 ;
      RECT 29.035000  56.755000 29.565000  57.285000 ;
      RECT 29.390000  18.965000 30.080000  23.745000 ;
      RECT 29.390000  32.250000 29.920000  37.330000 ;
      RECT 30.165000  32.250000 30.695000  37.000000 ;
      RECT 30.270000  18.995000 30.800000  23.745000 ;
      RECT 30.950000  32.250000 31.375000  37.330000 ;
      RECT 31.660000  32.250000 32.085000  37.005000 ;
      RECT 31.820000  18.995000 32.350000  23.745000 ;
      RECT 32.410000  32.060000 33.070000  36.750000 ;
      RECT 33.500000  31.990000 33.930000  37.080000 ;
      RECT 34.305000  31.975000 34.865000  36.750000 ;
      RECT 35.060000  31.990000 35.490000  37.080000 ;
      RECT 35.865000  31.975000 36.425000  36.750000 ;
      RECT 35.870000  26.885000 36.305000  28.235000 ;
      RECT 36.620000  31.990000 37.050000  37.080000 ;
      RECT 37.425000  31.975000 37.985000  36.750000 ;
      RECT 38.180000  31.990000 38.610000  37.080000 ;
      RECT 38.985000  31.975000 39.545000  36.750000 ;
      RECT 39.270000  26.885000 39.690000  28.235000 ;
      RECT 39.685000  95.955000 45.710000  96.105000 ;
      RECT 39.715000  31.990000 40.090000  36.750000 ;
      RECT 40.580000  32.155000 40.900000  36.710000 ;
      RECT 43.380000  24.850000 43.870000  27.560000 ;
      RECT 43.855000 180.205000 44.500000 180.370000 ;
      RECT 44.200000  33.270000 44.390000  36.510000 ;
      RECT 45.310000  36.340000 46.360000  36.970000 ;
      RECT 49.340000  32.065000 51.760000  32.445000 ;
      RECT 51.105000  32.445000 51.760000  33.690000 ;
      RECT 52.050000  24.855000 52.580000  27.565000 ;
      RECT 53.470000  24.855000 54.000000  27.565000 ;
      RECT 54.870000  24.855000 55.400000  27.565000 ;
      RECT 56.725000 180.205000 57.305000 180.370000 ;
      RECT 59.360000   2.260000 59.720000   3.430000 ;
      RECT 61.115000   5.230000 67.290000   5.345000 ;
      RECT 61.115000   5.345000 67.100000   5.400000 ;
      RECT 61.370000   5.080000 67.290000   5.230000 ;
      RECT 61.560000   4.765000 67.290000   5.080000 ;
      RECT 64.375000   0.250000 66.075000   1.000000 ;
      RECT 65.660000   6.230000 67.100000   9.570000 ;
      RECT 66.390000   9.570000 67.100000   9.575000 ;
      RECT 66.390000   9.575000 69.665000   9.745000 ;
      RECT 66.390000   9.745000 71.650000  10.185000 ;
      RECT 68.290000   1.940000 69.255000   3.960000 ;
      RECT 69.165000 128.445000 79.585000 130.115000 ;
      RECT 69.625000 179.435000 77.885000 179.450000 ;
      RECT 69.625000 179.980000 77.885000 180.205000 ;
      RECT 69.665000  10.185000 71.650000  11.425000 ;
      RECT 72.315000   1.940000 74.335000   4.420000 ;
      RECT 73.080000   8.080000 74.910000   8.830000 ;
      RECT 74.910000   5.170000 76.930000   5.800000 ;
      RECT 74.910000   5.800000 79.430000   7.820000 ;
      RECT 77.195000   3.705000 79.430000   4.420000 ;
      RECT 77.195000   4.420000 77.775000   5.170000 ;
      RECT 77.410000   3.700000 79.430000   3.705000 ;
      RECT 77.410000   7.820000 79.430000   8.080000 ;
      RECT 79.880000  19.485000 80.120000  25.015000 ;
      RECT 79.880000  30.115000 80.120000  35.725000 ;
    LAYER met1 ;
      RECT -0.115000  95.895000  1.495000 130.220000 ;
      RECT -0.115000 131.275000  1.495000 170.090000 ;
      RECT  0.000000   0.000000  5.565000   1.560000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000 62.290000   2.055000 ;
      RECT  0.000000   1.560000  5.565000   1.565000 ;
      RECT  0.000000   1.565000  5.565000   2.055000 ;
      RECT  0.000000   1.565000 35.575000   1.635000 ;
      RECT  0.000000   1.635000 35.505000   1.705000 ;
      RECT  0.000000   1.705000 35.435000   1.775000 ;
      RECT  0.000000   1.775000 35.365000   1.845000 ;
      RECT  0.000000   1.845000 35.295000   1.915000 ;
      RECT  0.000000   1.915000 35.225000   1.985000 ;
      RECT  0.000000   1.985000 35.155000   2.055000 ;
      RECT  0.000000   2.055000  5.565000   2.875000 ;
      RECT  0.000000   2.055000 80.000000 106.585000 ;
      RECT  0.000000   2.875000 11.260000   3.155000 ;
      RECT  0.000000   3.155000 67.995000   4.240000 ;
      RECT  0.000000   3.155000 67.995000  10.335000 ;
      RECT  0.000000   3.155000 67.995000  10.335000 ;
      RECT  0.000000   3.155000 67.995000  10.335000 ;
      RECT  0.000000   4.240000 76.885000   5.515000 ;
      RECT  0.000000   4.240000 76.885000  10.335000 ;
      RECT  0.000000   4.240000 76.885000  10.335000 ;
      RECT  0.000000   4.240000 76.885000  10.335000 ;
      RECT  0.000000   5.515000 80.000000  10.335000 ;
      RECT  0.000000  10.335000  1.340000  11.155000 ;
      RECT  0.000000  11.155000  0.750000  12.425000 ;
      RECT  0.000000  12.425000 80.000000  13.120000 ;
      RECT  0.000000  14.320000 76.495000  23.850000 ;
      RECT  0.000000  14.320000 80.000000  16.455000 ;
      RECT  0.000000  17.275000 78.550000  23.850000 ;
      RECT  0.000000  17.275000 78.550000  29.840000 ;
      RECT  0.000000  17.275000 79.605000  19.205000 ;
      RECT  0.000000  17.275000 79.605000  20.650000 ;
      RECT  0.000000  17.275000 79.605000  20.650000 ;
      RECT  0.000000  19.205000 79.605000  20.650000 ;
      RECT  0.000000  20.650000 78.550000  29.840000 ;
      RECT  0.000000  20.650000 79.535000  20.720000 ;
      RECT  0.000000  20.650000 79.535000  20.720000 ;
      RECT  0.000000  20.720000 79.465000  20.790000 ;
      RECT  0.000000  20.720000 79.465000  20.790000 ;
      RECT  0.000000  20.790000 79.395000  20.860000 ;
      RECT  0.000000  20.790000 79.395000  20.860000 ;
      RECT  0.000000  20.860000 79.325000  20.930000 ;
      RECT  0.000000  20.860000 79.325000  20.930000 ;
      RECT  0.000000  20.930000 79.255000  21.000000 ;
      RECT  0.000000  20.930000 79.255000  21.000000 ;
      RECT  0.000000  21.000000 79.185000  21.070000 ;
      RECT  0.000000  21.000000 79.185000  21.070000 ;
      RECT  0.000000  21.070000 79.160000  21.095000 ;
      RECT  0.000000  21.070000 79.160000  21.095000 ;
      RECT  0.000000  23.405000 79.160000  23.475000 ;
      RECT  0.000000  23.405000 79.160000  23.475000 ;
      RECT  0.000000  23.475000 79.230000  23.545000 ;
      RECT  0.000000  23.475000 79.230000  23.545000 ;
      RECT  0.000000  23.545000 79.300000  23.615000 ;
      RECT  0.000000  23.545000 79.300000  23.615000 ;
      RECT  0.000000  23.615000 79.370000  23.685000 ;
      RECT  0.000000  23.615000 79.370000  23.685000 ;
      RECT  0.000000  23.685000 79.440000  23.755000 ;
      RECT  0.000000  23.685000 79.440000  23.755000 ;
      RECT  0.000000  23.755000 79.510000  23.825000 ;
      RECT  0.000000  23.755000 79.510000  23.825000 ;
      RECT  0.000000  23.825000 79.580000  23.850000 ;
      RECT  0.000000  23.825000 79.580000  23.850000 ;
      RECT  0.000000  23.850000 79.605000  25.295000 ;
      RECT  0.000000  25.295000 78.845000  36.005000 ;
      RECT  0.000000  25.295000 78.845000  42.035000 ;
      RECT  0.000000  25.295000 80.000000  29.840000 ;
      RECT  0.000000  29.840000 78.845000  42.035000 ;
      RECT  0.000000  29.840000 79.605000  31.400000 ;
      RECT  0.000000  31.400000 79.535000  31.470000 ;
      RECT  0.000000  31.400000 79.535000  31.470000 ;
      RECT  0.000000  31.470000 79.465000  31.540000 ;
      RECT  0.000000  31.470000 79.465000  31.540000 ;
      RECT  0.000000  31.540000 79.395000  31.610000 ;
      RECT  0.000000  31.540000 79.395000  31.610000 ;
      RECT  0.000000  31.610000 79.325000  31.680000 ;
      RECT  0.000000  31.610000 79.325000  31.680000 ;
      RECT  0.000000  31.680000 79.280000  31.725000 ;
      RECT  0.000000  31.680000 79.280000  31.725000 ;
      RECT  0.000000  31.725000 78.845000  34.115000 ;
      RECT  0.000000  34.115000 79.280000  34.185000 ;
      RECT  0.000000  34.115000 79.280000  34.185000 ;
      RECT  0.000000  34.185000 79.350000  34.255000 ;
      RECT  0.000000  34.185000 79.350000  34.255000 ;
      RECT  0.000000  34.255000 79.420000  34.325000 ;
      RECT  0.000000  34.255000 79.420000  34.325000 ;
      RECT  0.000000  34.325000 79.490000  34.395000 ;
      RECT  0.000000  34.325000 79.490000  34.395000 ;
      RECT  0.000000  34.395000 79.560000  34.440000 ;
      RECT  0.000000  34.395000 79.560000  34.440000 ;
      RECT  0.000000  34.440000 79.605000  36.005000 ;
      RECT  0.000000  36.005000 80.000000  42.035000 ;
      RECT  0.000000  42.035000 78.635000  42.340000 ;
      RECT  0.000000  42.340000 78.565000  42.410000 ;
      RECT  0.000000  42.340000 78.565000  42.410000 ;
      RECT  0.000000  42.410000 78.495000  42.480000 ;
      RECT  0.000000  42.410000 78.495000  42.480000 ;
      RECT  0.000000  42.480000 78.425000  42.550000 ;
      RECT  0.000000  42.480000 78.425000  42.550000 ;
      RECT  0.000000  42.550000 78.355000  42.620000 ;
      RECT  0.000000  42.550000 78.355000  42.620000 ;
      RECT  0.000000  42.620000 78.285000  42.690000 ;
      RECT  0.000000  42.620000 78.285000  42.690000 ;
      RECT  0.000000  42.690000 78.215000  42.760000 ;
      RECT  0.000000  42.690000 78.215000  42.760000 ;
      RECT  0.000000  42.760000 78.145000  42.830000 ;
      RECT  0.000000  42.760000 78.145000  42.830000 ;
      RECT  0.000000  42.830000 78.075000  42.900000 ;
      RECT  0.000000  42.830000 78.075000  42.900000 ;
      RECT  0.000000  42.900000 78.005000  42.970000 ;
      RECT  0.000000  42.900000 78.005000  42.970000 ;
      RECT  0.000000  42.970000 78.000000  42.975000 ;
      RECT  0.000000  42.970000 78.000000  42.975000 ;
      RECT  0.000000  42.975000 78.635000  43.235000 ;
      RECT  0.000000  43.235000 80.000000  44.355000 ;
      RECT  0.000000  44.355000  1.020000  45.010000 ;
      RECT  0.000000  45.010000  0.965000  45.240000 ;
      RECT  0.000000  45.240000  0.895000  45.310000 ;
      RECT  0.000000  45.310000  0.825000  45.380000 ;
      RECT  0.000000  45.380000  0.755000  45.450000 ;
      RECT  0.000000  45.450000  0.685000  45.520000 ;
      RECT  0.000000  45.520000  0.615000  45.590000 ;
      RECT  0.000000  45.590000  0.545000  45.660000 ;
      RECT  0.000000  45.660000  0.475000  45.730000 ;
      RECT  0.000000  45.730000  0.405000  45.800000 ;
      RECT  0.000000  45.800000  0.335000  45.870000 ;
      RECT  0.000000  45.870000  0.265000  45.940000 ;
      RECT  0.000000  45.940000  0.195000  46.010000 ;
      RECT  0.000000  46.010000  0.125000  46.080000 ;
      RECT  0.000000  46.080000  0.055000  46.150000 ;
      RECT  0.000000  46.445000  0.965000  46.580000 ;
      RECT  0.000000  46.580000  1.050000  47.350000 ;
      RECT  0.000000  47.350000 80.000000  93.020000 ;
      RECT  0.000000  93.020000  1.070000  94.660000 ;
      RECT  0.000000  94.660000 11.550000  94.830000 ;
      RECT  0.000000  94.830000  1.985000  95.615000 ;
      RECT  0.000000 118.955000 80.000000 200.000000 ;
      RECT  0.000000 130.500000  4.530000 130.715000 ;
      RECT  0.000000 130.715000  1.980000 130.995000 ;
      RECT  0.000000 170.370000  1.980000 178.680000 ;
      RECT  0.000000 178.680000 15.445000 198.405000 ;
      RECT  0.000000 178.680000 15.445000 198.405000 ;
      RECT  0.000000 178.680000 80.000000 179.140000 ;
      RECT  0.000000 179.140000 15.445000 180.290000 ;
      RECT  0.000000 180.290000 15.490000 200.000000 ;
      RECT  0.000000 180.290000 80.000000 198.405000 ;
      RECT  0.000000 198.405000 15.490000 200.000000 ;
      RECT  0.210000  13.400000  0.470000  14.040000 ;
      RECT  0.475000  46.125000  5.000000  46.165000 ;
      RECT  0.545000  46.055000  5.000000  46.125000 ;
      RECT  0.615000  45.985000  5.000000  46.055000 ;
      RECT  0.685000  45.915000  5.000000  45.985000 ;
      RECT  0.750000  11.155000 76.825000  12.425000 ;
      RECT  0.750000  13.120000 80.000000  16.125000 ;
      RECT  0.755000  45.845000  5.000000  45.915000 ;
      RECT  0.825000  45.775000  5.000000  45.845000 ;
      RECT  0.895000  45.705000  5.000000  45.775000 ;
      RECT  0.965000  45.635000  5.000000  45.705000 ;
      RECT  1.035000  45.565000  5.000000  45.635000 ;
      RECT  1.105000  45.495000  5.000000  45.565000 ;
      RECT  1.175000  45.425000  5.000000  45.495000 ;
      RECT  1.245000  45.290000  5.000000  45.355000 ;
      RECT  1.245000  45.355000  5.000000  45.425000 ;
      RECT  1.245000  46.165000  5.000000  46.300000 ;
      RECT  1.300000  44.635000  1.730000  45.290000 ;
      RECT  1.330000  46.300000  2.790000  47.070000 ;
      RECT  1.350000  93.300000  8.265000  94.380000 ;
      RECT  1.620000  10.615000  4.025000  10.875000 ;
      RECT  1.775000  95.615000  1.985000 106.585000 ;
      RECT  1.775000 118.955000  1.985000 130.500000 ;
      RECT  1.775000 130.995000  1.980000 140.430000 ;
      RECT  1.775000 140.430000 80.000000 144.875000 ;
      RECT  1.775000 144.875000  1.980000 170.370000 ;
      RECT  2.000000 106.585000 80.000000 118.955000 ;
      RECT  2.010000  44.355000 80.000000  45.010000 ;
      RECT  2.260000 130.995000  4.700000 139.510000 ;
      RECT  2.260000 139.510000  4.855000 140.150000 ;
      RECT  2.260000 145.155000  4.700000 178.400000 ;
      RECT  2.265000  95.110000  8.970000  95.900000 ;
      RECT  2.265000  95.900000  4.250000 130.220000 ;
      RECT  3.070000  46.580000 80.000000  47.350000 ;
      RECT  3.070000  46.580000 80.000000  93.020000 ;
      RECT  3.070000  46.580000 80.000000  93.020000 ;
      RECT  3.070000  46.580000 80.000000  93.020000 ;
      RECT  4.305000   8.145000 80.000000  11.150000 ;
      RECT  4.305000  11.150000 76.825000  11.155000 ;
      RECT  4.530000  96.180000 80.000000 127.980000 ;
      RECT  4.530000 125.130000 70.100000 128.135000 ;
      RECT  4.530000 128.135000 68.825000 130.425000 ;
      RECT  4.530000 130.425000 70.100000 130.500000 ;
      RECT  4.530000 130.500000 80.000000 130.715000 ;
      RECT  4.980000 130.715000 80.000000 139.230000 ;
      RECT  4.980000 144.875000 80.000000 178.680000 ;
      RECT  4.980000 144.875000 80.000000 179.140000 ;
      RECT  4.980000 144.875000 80.000000 179.140000 ;
      RECT  5.135000 139.230000 80.000000 140.430000 ;
      RECT  5.135000 139.230000 80.000000 144.875000 ;
      RECT  5.280000  43.235000 80.000000  46.580000 ;
      RECT  5.280000  43.235000 80.000000  46.580000 ;
      RECT  5.280000  43.235000 80.000000  47.350000 ;
      RECT  5.280000  43.235000 80.000000  93.020000 ;
      RECT  5.280000  43.235000 80.000000  93.020000 ;
      RECT  5.280000  43.235000 80.000000  93.020000 ;
      RECT  5.280000  45.010000 80.000000  46.580000 ;
      RECT  5.565000   0.000000  6.890000   1.560000 ;
      RECT  5.565000   1.560000 22.990000   1.565000 ;
      RECT  5.845000   2.335000 10.120000   2.595000 ;
      RECT  7.170000   0.270000 10.715000   1.280000 ;
      RECT  8.545000  93.020000 11.550000  94.660000 ;
      RECT  9.250000  47.350000 80.000000 127.980000 ;
      RECT  9.250000  47.350000 80.000000 127.980000 ;
      RECT  9.250000  47.350000 80.000000 127.980000 ;
      RECT 10.400000   2.055000 35.085000   2.125000 ;
      RECT 10.400000   2.125000 35.015000   2.195000 ;
      RECT 10.400000   2.195000 34.945000   2.265000 ;
      RECT 10.400000   2.265000 34.880000   2.330000 ;
      RECT 10.400000   2.330000 13.640000   2.335000 ;
      RECT 10.400000   2.335000 11.260000   2.875000 ;
      RECT 10.995000   0.000000 18.955000   1.560000 ;
      RECT 11.540000   2.615000 35.170000   2.685000 ;
      RECT 11.540000   2.685000 35.100000   2.755000 ;
      RECT 11.540000   2.755000 35.070000   2.785000 ;
      RECT 11.540000   2.785000 18.385000   2.790000 ;
      RECT 11.540000   2.790000 13.990000   2.795000 ;
      RECT 11.540000   2.795000 13.985000   2.800000 ;
      RECT 11.540000   2.800000 12.220000   2.835000 ;
      RECT 11.540000   2.835000 12.185000   2.870000 ;
      RECT 11.540000   2.870000 12.180000   2.875000 ;
      RECT 12.300000   3.150000 67.995000   3.155000 ;
      RECT 12.300000   3.150000 67.995000   3.155000 ;
      RECT 12.310000   3.140000 67.995000   3.150000 ;
      RECT 12.310000   3.140000 67.995000   3.150000 ;
      RECT 12.320000   3.130000 67.995000   3.140000 ;
      RECT 12.320000   3.130000 67.995000   3.140000 ;
      RECT 12.345000   3.105000 59.170000   3.130000 ;
      RECT 12.345000   3.105000 59.170000   3.130000 ;
      RECT 12.370000   3.080000 59.170000   3.105000 ;
      RECT 12.370000   3.080000 59.170000   3.105000 ;
      RECT 13.760000   2.610000 35.240000   2.615000 ;
      RECT 14.105000   3.075000 59.170000   3.080000 ;
      RECT 14.105000   3.075000 59.170000   3.080000 ;
      RECT 14.110000   3.070000 59.170000   3.075000 ;
      RECT 14.110000   3.070000 59.170000   3.075000 ;
      RECT 15.725000 179.420000 77.705000 180.010000 ;
      RECT 15.770000 198.685000 56.715000 199.975000 ;
      RECT 18.505000   3.065000 19.370000   3.070000 ;
      RECT 19.235000   0.270000 21.375000   1.280000 ;
      RECT 19.490000   2.785000 28.955000   2.790000 ;
      RECT 21.655000   0.000000 22.990000   1.560000 ;
      RECT 23.270000   0.275000 26.265000   1.285000 ;
      RECT 26.545000   0.000000 33.120000   1.560000 ;
      RECT 26.545000   1.560000 34.265000   1.565000 ;
      RECT 29.075000   3.065000 30.425000   3.070000 ;
      RECT 29.075000   3.065000 30.425000   3.070000 ;
      RECT 30.545000   2.785000 35.065000   2.790000 ;
      RECT 33.400000   0.270000 37.775000   1.280000 ;
      RECT 34.545000   1.280000 37.775000   1.285000 ;
      RECT 35.055000   2.550000 35.245000   2.610000 ;
      RECT 35.125000   2.480000 35.305000   2.550000 ;
      RECT 35.195000   2.410000 35.375000   2.480000 ;
      RECT 35.205000   3.045000 59.170000   3.070000 ;
      RECT 35.205000   3.045000 59.170000   3.070000 ;
      RECT 35.265000   2.340000 35.445000   2.410000 ;
      RECT 35.275000   2.975000 59.170000   3.045000 ;
      RECT 35.275000   2.975000 59.170000   3.045000 ;
      RECT 35.335000   2.270000 35.515000   2.340000 ;
      RECT 35.345000   2.905000 59.170000   2.975000 ;
      RECT 35.345000   2.905000 59.170000   2.975000 ;
      RECT 35.405000   2.200000 35.585000   2.270000 ;
      RECT 35.415000   2.835000 59.170000   2.905000 ;
      RECT 35.415000   2.835000 59.170000   2.905000 ;
      RECT 35.475000   2.130000 35.655000   2.200000 ;
      RECT 35.485000   2.765000 59.170000   2.835000 ;
      RECT 35.485000   2.765000 59.170000   2.835000 ;
      RECT 35.515000   2.090000 43.035000   2.130000 ;
      RECT 35.555000   2.695000 59.170000   2.765000 ;
      RECT 35.555000   2.695000 59.170000   2.765000 ;
      RECT 35.560000   2.690000 42.990000   2.695000 ;
      RECT 35.560000   2.690000 42.990000   2.695000 ;
      RECT 35.585000   2.020000 42.965000   2.090000 ;
      RECT 35.630000   2.620000 42.920000   2.690000 ;
      RECT 35.630000   2.620000 42.920000   2.690000 ;
      RECT 35.655000   1.950000 42.895000   2.020000 ;
      RECT 35.700000   2.550000 42.850000   2.620000 ;
      RECT 35.700000   2.550000 42.850000   2.620000 ;
      RECT 35.770000   2.480000 42.780000   2.550000 ;
      RECT 35.770000   2.480000 42.780000   2.550000 ;
      RECT 35.840000   2.410000 42.710000   2.480000 ;
      RECT 35.840000   2.410000 42.710000   2.480000 ;
      RECT 38.055000   0.000000 40.785000   1.145000 ;
      RECT 38.055000   1.145000 39.110000   1.670000 ;
      RECT 39.390000   1.425000 43.110000   1.495000 ;
      RECT 39.390000   1.495000 43.180000   1.565000 ;
      RECT 39.390000   1.565000 43.250000   1.635000 ;
      RECT 39.390000   1.635000 43.320000   1.685000 ;
      RECT 41.065000   0.270000 41.935000   1.285000 ;
      RECT 42.215000   0.000000 55.320000   1.145000 ;
      RECT 42.875000   2.130000 43.075000   2.180000 ;
      RECT 42.925000   2.180000 43.125000   2.230000 ;
      RECT 42.930000   2.230000 43.175000   2.235000 ;
      RECT 43.000000   2.235000 51.520000   2.305000 ;
      RECT 43.070000   2.305000 51.520000   2.375000 ;
      RECT 43.110000   1.685000 43.370000   1.755000 ;
      RECT 43.110000   2.375000 51.520000   2.415000 ;
      RECT 43.180000   1.755000 43.440000   1.825000 ;
      RECT 43.200000   1.825000 43.510000   1.845000 ;
      RECT 43.270000   1.145000 62.150000   1.190000 ;
      RECT 43.270000   1.845000 47.840000   1.915000 ;
      RECT 43.315000   1.190000 62.150000   1.235000 ;
      RECT 43.340000   1.915000 47.770000   1.985000 ;
      RECT 43.385000   1.235000 47.725000   1.305000 ;
      RECT 43.410000   1.985000 47.700000   2.055000 ;
      RECT 43.430000   2.055000 47.680000   2.075000 ;
      RECT 43.455000   1.305000 47.655000   1.375000 ;
      RECT 43.525000   1.375000 47.585000   1.445000 ;
      RECT 43.595000   1.445000 47.515000   1.515000 ;
      RECT 43.645000   1.515000 47.465000   1.565000 ;
      RECT 47.630000   1.795000 47.910000   1.845000 ;
      RECT 47.680000   1.745000 47.960000   1.795000 ;
      RECT 47.700000   1.725000 55.040000   1.745000 ;
      RECT 47.770000   1.655000 55.040000   1.725000 ;
      RECT 47.840000   1.585000 55.040000   1.655000 ;
      RECT 47.910000   1.515000 55.040000   1.585000 ;
      RECT 50.840000   2.195000 51.520000   2.235000 ;
      RECT 50.880000   2.155000 51.520000   2.195000 ;
      RECT 51.800000   2.025000 54.525000   2.095000 ;
      RECT 51.800000   2.025000 54.525000   2.095000 ;
      RECT 51.800000   2.095000 54.595000   2.165000 ;
      RECT 51.800000   2.095000 54.595000   2.165000 ;
      RECT 51.800000   2.165000 54.665000   2.235000 ;
      RECT 51.800000   2.165000 54.665000   2.235000 ;
      RECT 51.800000   2.235000 54.735000   2.305000 ;
      RECT 51.800000   2.235000 54.735000   2.305000 ;
      RECT 51.800000   2.305000 54.805000   2.375000 ;
      RECT 51.800000   2.305000 54.805000   2.375000 ;
      RECT 51.800000   2.375000 54.875000   2.445000 ;
      RECT 51.800000   2.375000 54.875000   2.445000 ;
      RECT 51.800000   2.445000 54.945000   2.515000 ;
      RECT 51.800000   2.445000 54.945000   2.515000 ;
      RECT 51.800000   2.515000 55.015000   2.585000 ;
      RECT 51.800000   2.515000 55.015000   2.585000 ;
      RECT 51.800000   2.585000 55.085000   2.655000 ;
      RECT 51.800000   2.585000 55.085000   2.655000 ;
      RECT 51.800000   2.655000 59.170000   2.695000 ;
      RECT 54.655000   1.745000 55.040000   1.760000 ;
      RECT 54.670000   1.760000 55.040000   1.775000 ;
      RECT 54.675000   1.775000 55.040000   1.780000 ;
      RECT 54.745000   1.780000 54.875000   1.850000 ;
      RECT 54.815000   1.850000 54.875000   1.920000 ;
      RECT 55.155000   2.060000 59.170000   2.655000 ;
      RECT 55.320000   0.000000 59.170000   1.145000 ;
      RECT 55.320000   1.145000 59.170000   1.235000 ;
      RECT 55.320000   1.235000 59.170000   1.920000 ;
      RECT 55.320000   1.920000 59.170000   2.060000 ;
      RECT 56.995000 180.290000 71.715000 200.000000 ;
      RECT 56.995000 180.290000 71.715000 200.000000 ;
      RECT 56.995000 180.290000 80.000000 198.420000 ;
      RECT 56.995000 180.290000 80.000000 198.420000 ;
      RECT 56.995000 198.405000 80.000000 198.420000 ;
      RECT 56.995000 198.420000 71.715000 200.000000 ;
      RECT 59.170000   0.000000 62.150000   1.145000 ;
      RECT 59.170000   1.235000 62.150000   1.920000 ;
      RECT 59.450000   2.200000 59.710000   2.850000 ;
      RECT 59.990000   1.920000 62.150000   2.195000 ;
      RECT 59.990000   2.195000 67.995000   3.130000 ;
      RECT 62.830000   0.000000 80.000000   2.055000 ;
      RECT 62.970000   0.000000 64.095000   1.190000 ;
      RECT 62.970000   1.190000 67.995000   1.960000 ;
      RECT 62.970000   1.960000 67.995000   2.195000 ;
      RECT 64.375000   0.260000 67.295000   0.910000 ;
      RECT 67.575000   0.000000 69.205000   1.190000 ;
      RECT 67.995000   1.190000 69.205000   1.960000 ;
      RECT 68.275000   2.240000 68.925000   3.960000 ;
      RECT 69.105000 128.415000 80.145000 130.145000 ;
      RECT 69.205000   0.000000 80.000000   1.190000 ;
      RECT 69.205000   1.190000 80.000000   1.960000 ;
      RECT 69.205000   1.960000 80.000000   3.365000 ;
      RECT 69.205000   3.365000 76.885000   4.240000 ;
      RECT 70.380000 128.260000 80.145000 128.415000 ;
      RECT 70.380000 130.145000 80.145000 130.220000 ;
      RECT 71.995000 198.700000 76.855000 200.000000 ;
      RECT 76.775000  16.735000 77.415000  16.995000 ;
      RECT 77.105000  11.430000 77.365000  12.145000 ;
      RECT 77.135000 198.420000 80.000000 200.000000 ;
      RECT 77.165000   3.645000 77.805000   5.235000 ;
      RECT 77.645000  11.150000 80.000000  12.425000 ;
      RECT 77.695000  16.455000 80.000000  17.275000 ;
      RECT 77.985000 179.140000 80.000000 180.290000 ;
      RECT 78.085000   3.365000 80.000000   5.515000 ;
      RECT 78.705000  42.665000 79.175000  42.695000 ;
      RECT 78.775000  42.595000 79.175000  42.665000 ;
      RECT 78.830000  21.375000 80.115000  23.125000 ;
      RECT 78.845000  42.525000 79.175000  42.595000 ;
      RECT 78.915000  42.315000 79.175000  42.455000 ;
      RECT 78.915000  42.455000 79.175000  42.525000 ;
      RECT 78.915000  42.695000 79.175000  42.955000 ;
      RECT 79.125000  32.005000 80.115000  33.835000 ;
      RECT 79.325000  21.325000 80.115000  21.375000 ;
      RECT 79.345000  23.125000 80.115000  23.195000 ;
      RECT 79.395000  21.255000 80.115000  21.325000 ;
      RECT 79.415000  23.195000 80.115000  23.265000 ;
      RECT 79.455000  42.035000 80.000000  43.235000 ;
      RECT 79.465000  21.185000 80.115000  21.255000 ;
      RECT 79.465000  31.935000 80.115000  32.005000 ;
      RECT 79.465000  33.835000 80.115000  33.905000 ;
      RECT 79.485000  23.265000 80.115000  23.335000 ;
      RECT 79.535000  21.115000 80.115000  21.185000 ;
      RECT 79.535000  31.865000 80.115000  31.935000 ;
      RECT 79.535000  33.905000 80.115000  33.975000 ;
      RECT 79.555000  23.335000 80.115000  23.405000 ;
      RECT 79.605000  17.275000 80.000000  19.205000 ;
      RECT 79.605000  21.045000 80.115000  21.115000 ;
      RECT 79.605000  31.795000 80.115000  31.865000 ;
      RECT 79.605000  33.975000 80.115000  34.045000 ;
      RECT 79.625000  23.405000 80.115000  23.475000 ;
      RECT 79.675000  20.975000 80.115000  21.045000 ;
      RECT 79.675000  31.725000 80.115000  31.795000 ;
      RECT 79.675000  34.045000 80.115000  34.115000 ;
      RECT 79.695000  23.475000 80.115000  23.545000 ;
      RECT 79.745000  20.905000 80.115000  20.975000 ;
      RECT 79.745000  31.655000 80.115000  31.725000 ;
      RECT 79.745000  34.115000 80.115000  34.185000 ;
      RECT 79.765000  23.545000 80.115000  23.615000 ;
      RECT 79.815000  20.835000 80.115000  20.905000 ;
      RECT 79.815000  31.585000 80.115000  31.655000 ;
      RECT 79.815000  34.185000 80.115000  34.255000 ;
      RECT 79.835000  23.615000 80.115000  23.685000 ;
      RECT 79.885000  19.485000 80.115000  20.765000 ;
      RECT 79.885000  20.765000 80.115000  20.835000 ;
      RECT 79.885000  23.685000 80.115000  23.735000 ;
      RECT 79.885000  23.735000 80.115000  25.015000 ;
      RECT 79.885000  30.120000 80.115000  31.515000 ;
      RECT 79.885000  31.515000 80.115000  31.585000 ;
      RECT 79.885000  34.255000 80.115000  34.325000 ;
      RECT 79.885000  34.325000 80.115000  35.725000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  3.095000   4.590000 ;
      RECT  0.000000   0.000000  3.235000   4.535000 ;
      RECT  0.000000   4.535000  3.940000   5.240000 ;
      RECT  0.000000   4.590000  3.095000   4.660000 ;
      RECT  0.000000   4.590000  3.095000   4.660000 ;
      RECT  0.000000   4.660000  3.165000   4.730000 ;
      RECT  0.000000   4.660000  3.165000   4.730000 ;
      RECT  0.000000   4.730000  3.235000   4.800000 ;
      RECT  0.000000   4.730000  3.235000   4.800000 ;
      RECT  0.000000   4.800000  3.305000   4.870000 ;
      RECT  0.000000   4.800000  3.305000   4.870000 ;
      RECT  0.000000   4.870000  3.375000   4.940000 ;
      RECT  0.000000   4.870000  3.375000   4.940000 ;
      RECT  0.000000   4.940000  3.445000   5.010000 ;
      RECT  0.000000   4.940000  3.445000   5.010000 ;
      RECT  0.000000   5.010000  3.515000   5.080000 ;
      RECT  0.000000   5.010000  3.515000   5.080000 ;
      RECT  0.000000   5.080000  3.585000   5.150000 ;
      RECT  0.000000   5.080000  3.585000   5.150000 ;
      RECT  0.000000   5.150000  3.655000   5.220000 ;
      RECT  0.000000   5.150000  3.655000   5.220000 ;
      RECT  0.000000   5.220000  3.725000   5.290000 ;
      RECT  0.000000   5.220000  3.725000   5.290000 ;
      RECT  0.000000   5.240000  5.260000   5.435000 ;
      RECT  0.000000   5.290000  3.795000   5.360000 ;
      RECT  0.000000   5.290000  3.795000   5.360000 ;
      RECT  0.000000   5.360000  3.865000   5.380000 ;
      RECT  0.000000   5.360000  3.865000   5.380000 ;
      RECT  0.000000   5.380000  5.010000   5.435000 ;
      RECT  0.000000   5.380000  5.010000   5.435000 ;
      RECT  0.000000   5.435000  5.065000   5.490000 ;
      RECT  0.000000   5.435000  5.065000   5.490000 ;
      RECT  0.000000   5.435000  5.260000   8.410000 ;
      RECT  0.000000   5.490000  5.120000   8.495000 ;
      RECT  0.000000   8.410000  6.435000   9.585000 ;
      RECT  0.000000   8.465000  5.120000   8.535000 ;
      RECT  0.000000   8.465000  5.120000   8.535000 ;
      RECT  0.000000   8.535000  5.190000   8.605000 ;
      RECT  0.000000   8.535000  5.190000   8.605000 ;
      RECT  0.000000   8.605000  5.260000   8.675000 ;
      RECT  0.000000   8.605000  5.260000   8.675000 ;
      RECT  0.000000   8.675000  5.330000   8.745000 ;
      RECT  0.000000   8.675000  5.330000   8.745000 ;
      RECT  0.000000   8.745000  5.400000   8.815000 ;
      RECT  0.000000   8.745000  5.400000   8.815000 ;
      RECT  0.000000   8.815000  5.470000   8.885000 ;
      RECT  0.000000   8.815000  5.470000   8.885000 ;
      RECT  0.000000   8.885000  5.540000   8.955000 ;
      RECT  0.000000   8.885000  5.540000   8.955000 ;
      RECT  0.000000   8.955000  5.610000   9.025000 ;
      RECT  0.000000   8.955000  5.610000   9.025000 ;
      RECT  0.000000   9.025000  5.680000   9.095000 ;
      RECT  0.000000   9.025000  5.680000   9.095000 ;
      RECT  0.000000   9.095000  5.750000   9.165000 ;
      RECT  0.000000   9.095000  5.750000   9.165000 ;
      RECT  0.000000   9.165000  5.820000   9.235000 ;
      RECT  0.000000   9.165000  5.820000   9.235000 ;
      RECT  0.000000   9.235000  5.890000   9.305000 ;
      RECT  0.000000   9.235000  5.890000   9.305000 ;
      RECT  0.000000   9.305000  5.960000   9.375000 ;
      RECT  0.000000   9.305000  5.960000   9.375000 ;
      RECT  0.000000   9.375000  6.030000   9.445000 ;
      RECT  0.000000   9.375000  6.030000   9.445000 ;
      RECT  0.000000   9.445000  6.100000   9.515000 ;
      RECT  0.000000   9.445000  6.100000   9.515000 ;
      RECT  0.000000   9.515000  6.170000   9.585000 ;
      RECT  0.000000   9.515000  6.170000   9.585000 ;
      RECT  0.000000   9.585000  6.240000   9.640000 ;
      RECT  0.000000   9.585000  6.240000   9.640000 ;
      RECT  0.000000   9.585000  6.435000  38.760000 ;
      RECT  0.000000   9.640000  6.295000  38.705000 ;
      RECT  0.000000  38.705000  6.225000  38.775000 ;
      RECT  0.000000  38.705000  6.225000  38.775000 ;
      RECT  0.000000  38.760000  5.835000  39.360000 ;
      RECT  0.000000  38.775000  6.155000  38.845000 ;
      RECT  0.000000  38.775000  6.155000  38.845000 ;
      RECT  0.000000  38.845000  6.085000  38.915000 ;
      RECT  0.000000  38.845000  6.085000  38.915000 ;
      RECT  0.000000  38.915000  6.015000  38.985000 ;
      RECT  0.000000  38.915000  6.015000  38.985000 ;
      RECT  0.000000  38.985000  5.945000  39.055000 ;
      RECT  0.000000  38.985000  5.945000  39.055000 ;
      RECT  0.000000  39.055000  5.875000  39.125000 ;
      RECT  0.000000  39.055000  5.875000  39.125000 ;
      RECT  0.000000  39.125000  5.805000  39.195000 ;
      RECT  0.000000  39.125000  5.805000  39.195000 ;
      RECT  0.000000  39.195000  5.735000  39.265000 ;
      RECT  0.000000  39.195000  5.735000  39.265000 ;
      RECT  0.000000  39.265000  5.695000  39.305000 ;
      RECT  0.000000  39.265000  5.695000  39.305000 ;
      RECT  0.000000  39.305000  5.685000  53.625000 ;
      RECT  0.000000  39.305000  5.695000  42.860000 ;
      RECT  0.000000  39.360000  5.835000  42.915000 ;
      RECT  0.000000  42.860000  5.690000  42.865000 ;
      RECT  0.000000  42.860000  5.690000  42.865000 ;
      RECT  0.000000  42.865000  5.685000  42.870000 ;
      RECT  0.000000  42.865000  5.685000  42.870000 ;
      RECT  0.000000  42.870000  5.685000  43.905000 ;
      RECT  0.000000  42.915000  5.825000  42.925000 ;
      RECT  0.000000  42.925000  5.825000  43.765000 ;
      RECT  0.000000  43.765000  8.055000  44.015000 ;
      RECT  0.000000  43.905000  7.915000  53.625000 ;
      RECT  0.000000  43.905000  7.945000  43.930000 ;
      RECT  0.000000  43.905000  7.945000  43.930000 ;
      RECT  0.000000  43.930000  7.920000  43.955000 ;
      RECT  0.000000  43.930000  7.920000  43.955000 ;
      RECT  0.000000  43.955000  7.915000  43.960000 ;
      RECT  0.000000  43.955000  7.915000  43.960000 ;
      RECT  0.000000  43.960000  7.915000  53.625000 ;
      RECT  0.000000  44.015000  8.055000  53.680000 ;
      RECT  0.000000  53.625000  7.845000  53.695000 ;
      RECT  0.000000  53.625000  7.845000  53.695000 ;
      RECT  0.000000  53.680000  7.835000  53.900000 ;
      RECT  0.000000  53.695000  7.775000  53.765000 ;
      RECT  0.000000  53.695000  7.775000  53.765000 ;
      RECT  0.000000  53.765000  7.705000  53.835000 ;
      RECT  0.000000  53.765000  7.705000  53.835000 ;
      RECT  0.000000  53.835000  7.695000  53.845000 ;
      RECT  0.000000  53.835000  7.695000  53.845000 ;
      RECT  0.000000  53.845000  7.695000  55.685000 ;
      RECT  0.000000  53.900000  7.835000  55.740000 ;
      RECT  0.000000  55.685000  7.035000  73.840000 ;
      RECT  0.000000  55.685000  7.035000  73.840000 ;
      RECT  0.000000  55.685000  7.035000  73.840000 ;
      RECT  0.000000  55.685000  7.035000  73.840000 ;
      RECT  0.000000  55.685000  7.625000  55.755000 ;
      RECT  0.000000  55.685000  7.625000  55.755000 ;
      RECT  0.000000  55.740000  7.175000  56.400000 ;
      RECT  0.000000  55.755000  7.555000  55.825000 ;
      RECT  0.000000  55.755000  7.555000  55.825000 ;
      RECT  0.000000  55.825000  7.485000  55.895000 ;
      RECT  0.000000  55.825000  7.485000  55.895000 ;
      RECT  0.000000  55.895000  7.415000  55.965000 ;
      RECT  0.000000  55.895000  7.415000  55.965000 ;
      RECT  0.000000  55.965000  7.345000  56.035000 ;
      RECT  0.000000  55.965000  7.345000  56.035000 ;
      RECT  0.000000  56.035000  7.275000  56.105000 ;
      RECT  0.000000  56.035000  7.275000  56.105000 ;
      RECT  0.000000  56.105000  7.205000  56.175000 ;
      RECT  0.000000  56.105000  7.205000  56.175000 ;
      RECT  0.000000  56.175000  7.135000  56.245000 ;
      RECT  0.000000  56.175000  7.135000  56.245000 ;
      RECT  0.000000  56.245000  7.065000  56.315000 ;
      RECT  0.000000  56.245000  7.065000  56.315000 ;
      RECT  0.000000  56.315000  7.035000  56.345000 ;
      RECT  0.000000  56.315000  7.035000  56.345000 ;
      RECT  0.000000  56.400000  7.175000  73.785000 ;
      RECT  0.000000  73.785000  7.665000  74.270000 ;
      RECT  0.000000  73.840000  7.035000  73.910000 ;
      RECT  0.000000  73.840000  7.035000  73.910000 ;
      RECT  0.000000  73.910000  7.105000  73.980000 ;
      RECT  0.000000  73.910000  7.105000  73.980000 ;
      RECT  0.000000  73.980000  7.175000  74.050000 ;
      RECT  0.000000  73.980000  7.175000  74.050000 ;
      RECT  0.000000  74.050000  7.245000  74.120000 ;
      RECT  0.000000  74.050000  7.245000  74.120000 ;
      RECT  0.000000  74.120000  7.315000  74.190000 ;
      RECT  0.000000  74.120000  7.315000  74.190000 ;
      RECT  0.000000  74.190000  7.385000  74.260000 ;
      RECT  0.000000  74.190000  7.385000  74.260000 ;
      RECT  0.000000  74.260000  7.455000  74.330000 ;
      RECT  0.000000  74.260000  7.455000  74.330000 ;
      RECT  0.000000  74.270000  7.665000  74.850000 ;
      RECT  0.000000  74.330000  7.525000  74.905000 ;
      RECT  0.000000  74.850000  8.070000  75.255000 ;
      RECT  0.000000  74.905000  7.525000  74.965000 ;
      RECT  0.000000  74.905000  7.525000  74.965000 ;
      RECT  0.000000  74.905000  7.525000  74.975000 ;
      RECT  0.000000  74.965000  7.585000  75.020000 ;
      RECT  0.000000  74.965000  7.585000  75.020000 ;
      RECT  0.000000  74.975000  7.595000  75.045000 ;
      RECT  0.000000  75.020000  7.640000  75.310000 ;
      RECT  0.000000  75.045000  7.665000  75.115000 ;
      RECT  0.000000  75.115000  7.735000  75.185000 ;
      RECT  0.000000  75.185000  7.805000  75.255000 ;
      RECT  0.000000  75.255000  7.875000  75.310000 ;
      RECT  0.000000  75.255000  8.070000  77.055000 ;
      RECT  0.000000  75.310000  7.930000  77.005000 ;
      RECT  0.000000  77.005000  7.640000  78.315000 ;
      RECT  0.000000  77.055000  7.980000  77.145000 ;
      RECT  0.000000  77.145000  7.780000  77.685000 ;
      RECT  0.000000  77.685000 76.775000  96.135000 ;
      RECT  0.000000  77.825000 76.635000  96.080000 ;
      RECT  0.000000  96.080000 76.565000  96.150000 ;
      RECT  0.000000  96.080000 76.565000  96.150000 ;
      RECT  0.000000  96.135000 76.545000  96.365000 ;
      RECT  0.000000  96.150000 76.495000  96.220000 ;
      RECT  0.000000  96.150000 76.495000  96.220000 ;
      RECT  0.000000  96.220000 76.425000  96.290000 ;
      RECT  0.000000  96.220000 76.425000  96.290000 ;
      RECT  0.000000  96.290000 76.355000  96.360000 ;
      RECT  0.000000  96.290000 76.355000  96.360000 ;
      RECT  0.000000  96.360000 76.285000  96.430000 ;
      RECT  0.000000  96.360000 76.285000  96.430000 ;
      RECT  0.000000  96.365000 80.000000 106.585000 ;
      RECT  0.000000  96.430000 76.215000  96.500000 ;
      RECT  0.000000  96.430000 76.215000  96.500000 ;
      RECT  0.000000  96.500000 76.210000  96.505000 ;
      RECT  0.000000  96.500000 76.210000  96.505000 ;
      RECT  0.000000  96.505000 80.000000 106.585000 ;
      RECT  0.000000 118.955000 80.000000 200.000000 ;
      RECT  0.000000 118.955000 80.000000 200.000000 ;
      RECT  0.740000 106.585000 80.000000 118.955000 ;
      RECT  2.000000 106.585000 80.000000 118.955000 ;
      RECT  3.745000   0.000000  5.280000   4.315000 ;
      RECT  3.745000   4.315000  5.280000   4.535000 ;
      RECT  3.885000   0.000000  5.140000   4.260000 ;
      RECT  3.955000   4.260000  5.140000   4.330000 ;
      RECT  3.960000   4.535000  5.475000   4.730000 ;
      RECT  4.025000   4.330000  5.140000   4.400000 ;
      RECT  4.095000   4.400000  5.140000   4.470000 ;
      RECT  4.165000   4.470000  5.140000   4.540000 ;
      RECT  4.215000   4.540000  5.140000   4.590000 ;
      RECT  5.285000   4.730000  5.965000   5.215000 ;
      RECT  5.770000   5.215000  6.180000   5.435000 ;
      RECT  5.770000   5.435000  6.180000   6.190000 ;
      RECT  5.770000   6.190000  6.085000   6.285000 ;
      RECT  5.770000   6.825000  8.305000   6.920000 ;
      RECT  5.770000   6.920000 13.830000   8.190000 ;
      RECT  5.770000   8.190000 13.830000   9.365000 ;
      RECT  5.790000   0.000000  5.990000   1.610000 ;
      RECT  5.790000   1.610000  8.305000   3.925000 ;
      RECT  5.790000   3.925000  8.305000   4.315000 ;
      RECT  5.790000   4.315000  8.305000   5.215000 ;
      RECT  5.845000   2.335000  6.520000   2.405000 ;
      RECT  5.845000   2.405000  6.590000   2.475000 ;
      RECT  5.845000   2.475000  6.660000   2.545000 ;
      RECT  5.845000   2.545000  6.730000   2.595000 ;
      RECT  5.885000   2.595000  6.780000   2.635000 ;
      RECT  5.910000   6.965000  8.165000   7.060000 ;
      RECT  5.910000   7.060000 13.690000   7.345000 ;
      RECT  5.910000   7.345000 13.690000   8.135000 ;
      RECT  5.925000   2.635000  6.820000   2.675000 ;
      RECT  5.930000   1.815000  6.000000   1.885000 ;
      RECT  5.930000   1.885000  6.070000   1.955000 ;
      RECT  5.930000   1.955000  6.140000   2.025000 ;
      RECT  5.930000   2.025000  6.210000   2.095000 ;
      RECT  5.930000   2.095000  6.280000   2.165000 ;
      RECT  5.930000   2.165000  6.350000   2.235000 ;
      RECT  5.930000   2.235000  6.420000   2.305000 ;
      RECT  5.930000   2.305000  6.490000   2.335000 ;
      RECT  5.930000   2.675000  6.860000   2.680000 ;
      RECT  5.930000   2.680000  6.865000   2.750000 ;
      RECT  5.930000   2.750000  6.935000   2.820000 ;
      RECT  5.930000   2.820000  7.005000   2.890000 ;
      RECT  5.930000   2.890000  7.075000   2.960000 ;
      RECT  5.930000   2.960000  7.145000   3.030000 ;
      RECT  5.930000   3.030000  7.215000   3.100000 ;
      RECT  5.930000   3.100000  7.285000   3.170000 ;
      RECT  5.930000   3.170000  7.355000   3.240000 ;
      RECT  5.930000   3.240000  7.425000   3.310000 ;
      RECT  5.930000   3.310000  7.495000   3.380000 ;
      RECT  5.930000   3.380000  7.565000   3.450000 ;
      RECT  5.930000   3.450000  7.635000   3.520000 ;
      RECT  5.930000   3.520000  7.705000   3.590000 ;
      RECT  5.930000   3.590000  7.775000   3.660000 ;
      RECT  5.930000   3.660000  7.845000   3.730000 ;
      RECT  5.930000   3.730000  7.915000   3.800000 ;
      RECT  5.930000   3.800000  7.985000   3.870000 ;
      RECT  5.930000   3.870000  8.055000   3.940000 ;
      RECT  5.930000   3.940000  8.125000   3.980000 ;
      RECT  5.930000   3.980000  8.165000   4.260000 ;
      RECT  5.980000   8.135000 13.690000   8.205000 ;
      RECT  5.980000   8.135000 13.690000   8.205000 ;
      RECT  6.000000   4.260000  8.165000   4.330000 ;
      RECT  6.050000   8.205000 13.690000   8.275000 ;
      RECT  6.050000   8.205000 13.690000   8.275000 ;
      RECT  6.070000   4.330000  8.165000   4.400000 ;
      RECT  6.120000   8.275000 13.690000   8.345000 ;
      RECT  6.120000   8.275000 13.690000   8.345000 ;
      RECT  6.140000   4.400000  8.165000   4.470000 ;
      RECT  6.190000   8.345000 13.690000   8.415000 ;
      RECT  6.190000   8.345000 13.690000   8.415000 ;
      RECT  6.210000   4.470000  8.165000   4.540000 ;
      RECT  6.260000   8.415000 13.690000   8.485000 ;
      RECT  6.260000   8.415000 13.690000   8.485000 ;
      RECT  6.280000   4.540000  8.165000   4.610000 ;
      RECT  6.330000   8.485000 13.690000   8.555000 ;
      RECT  6.330000   8.485000 13.690000   8.555000 ;
      RECT  6.345000  39.580000  9.165000  42.905000 ;
      RECT  6.345000  42.905000  9.145000  42.925000 ;
      RECT  6.350000   4.610000  8.165000   4.680000 ;
      RECT  6.365000  42.925000  8.305000  43.765000 ;
      RECT  6.400000   8.555000 13.690000   8.625000 ;
      RECT  6.400000   8.555000 13.690000   8.625000 ;
      RECT  6.420000   4.680000  8.165000   4.750000 ;
      RECT  6.470000   8.625000 13.690000   8.695000 ;
      RECT  6.470000   8.625000 13.690000   8.695000 ;
      RECT  6.485000  39.635000 12.170000  39.705000 ;
      RECT  6.485000  39.635000 12.170000  39.705000 ;
      RECT  6.485000  39.705000 12.100000  39.775000 ;
      RECT  6.485000  39.705000 12.100000  39.775000 ;
      RECT  6.485000  39.775000 12.030000  39.845000 ;
      RECT  6.485000  39.775000 12.030000  39.845000 ;
      RECT  6.485000  39.845000 11.960000  39.915000 ;
      RECT  6.485000  39.845000 11.960000  39.915000 ;
      RECT  6.485000  39.915000 11.890000  39.985000 ;
      RECT  6.485000  39.915000 11.890000  39.985000 ;
      RECT  6.485000  39.985000 11.820000  40.055000 ;
      RECT  6.485000  39.985000 11.820000  40.055000 ;
      RECT  6.485000  40.055000 11.750000  40.125000 ;
      RECT  6.485000  40.055000 11.750000  40.125000 ;
      RECT  6.485000  40.125000 11.680000  40.195000 ;
      RECT  6.485000  40.125000 11.680000  40.195000 ;
      RECT  6.485000  40.195000 11.610000  40.265000 ;
      RECT  6.485000  40.195000 11.610000  40.265000 ;
      RECT  6.485000  40.265000 11.540000  40.335000 ;
      RECT  6.485000  40.265000 11.540000  40.335000 ;
      RECT  6.485000  40.335000 11.470000  40.405000 ;
      RECT  6.485000  40.335000 11.470000  40.405000 ;
      RECT  6.485000  40.405000 11.400000  40.475000 ;
      RECT  6.485000  40.405000 11.400000  40.475000 ;
      RECT  6.485000  40.475000 11.330000  40.545000 ;
      RECT  6.485000  40.475000 11.330000  40.545000 ;
      RECT  6.485000  40.545000 11.260000  40.615000 ;
      RECT  6.485000  40.545000 11.260000  40.615000 ;
      RECT  6.485000  40.615000 11.190000  40.685000 ;
      RECT  6.485000  40.615000 11.190000  40.685000 ;
      RECT  6.485000  40.685000 11.120000  40.755000 ;
      RECT  6.485000  40.685000 11.120000  40.755000 ;
      RECT  6.485000  40.755000 11.050000  40.825000 ;
      RECT  6.485000  40.755000 11.050000  40.825000 ;
      RECT  6.485000  40.825000 10.980000  40.895000 ;
      RECT  6.485000  40.825000 10.980000  40.895000 ;
      RECT  6.485000  40.895000 10.910000  40.965000 ;
      RECT  6.485000  40.895000 10.910000  40.965000 ;
      RECT  6.485000  40.965000 10.840000  41.035000 ;
      RECT  6.485000  40.965000 10.840000  41.035000 ;
      RECT  6.485000  41.035000 10.770000  41.105000 ;
      RECT  6.485000  41.035000 10.770000  41.105000 ;
      RECT  6.485000  41.105000 10.700000  41.175000 ;
      RECT  6.485000  41.105000 10.700000  41.175000 ;
      RECT  6.485000  41.175000 10.630000  41.245000 ;
      RECT  6.485000  41.175000 10.630000  41.245000 ;
      RECT  6.485000  41.245000 10.560000  41.315000 ;
      RECT  6.485000  41.245000 10.560000  41.315000 ;
      RECT  6.485000  41.315000 10.490000  41.385000 ;
      RECT  6.485000  41.315000 10.490000  41.385000 ;
      RECT  6.485000  41.385000 10.420000  41.455000 ;
      RECT  6.485000  41.385000 10.420000  41.455000 ;
      RECT  6.485000  41.455000 10.350000  41.525000 ;
      RECT  6.485000  41.455000 10.350000  41.525000 ;
      RECT  6.485000  41.525000 10.280000  41.595000 ;
      RECT  6.485000  41.525000 10.280000  41.595000 ;
      RECT  6.485000  41.595000 10.210000  41.665000 ;
      RECT  6.485000  41.595000 10.210000  41.665000 ;
      RECT  6.485000  41.665000 10.140000  41.735000 ;
      RECT  6.485000  41.665000 10.140000  41.735000 ;
      RECT  6.485000  41.735000 10.070000  41.805000 ;
      RECT  6.485000  41.735000 10.070000  41.805000 ;
      RECT  6.485000  41.805000 10.000000  41.875000 ;
      RECT  6.485000  41.805000 10.000000  41.875000 ;
      RECT  6.485000  41.875000  9.930000  41.945000 ;
      RECT  6.485000  41.875000  9.930000  41.945000 ;
      RECT  6.485000  41.945000  9.860000  42.015000 ;
      RECT  6.485000  41.945000  9.860000  42.015000 ;
      RECT  6.485000  42.015000  9.790000  42.085000 ;
      RECT  6.485000  42.015000  9.790000  42.085000 ;
      RECT  6.485000  42.085000  9.720000  42.155000 ;
      RECT  6.485000  42.085000  9.720000  42.155000 ;
      RECT  6.485000  42.155000  9.650000  42.225000 ;
      RECT  6.485000  42.155000  9.650000  42.225000 ;
      RECT  6.485000  42.225000  9.580000  42.295000 ;
      RECT  6.485000  42.225000  9.580000  42.295000 ;
      RECT  6.485000  42.295000  9.510000  42.365000 ;
      RECT  6.485000  42.295000  9.510000  42.365000 ;
      RECT  6.485000  42.365000  9.440000  42.435000 ;
      RECT  6.485000  42.365000  9.440000  42.435000 ;
      RECT  6.485000  42.435000  9.370000  42.505000 ;
      RECT  6.485000  42.435000  9.370000  42.505000 ;
      RECT  6.485000  42.505000  9.300000  42.575000 ;
      RECT  6.485000  42.505000  9.300000  42.575000 ;
      RECT  6.485000  42.575000  9.230000  42.645000 ;
      RECT  6.485000  42.575000  9.230000  42.645000 ;
      RECT  6.485000  42.645000  9.160000  42.715000 ;
      RECT  6.485000  42.645000  9.160000  42.715000 ;
      RECT  6.485000  42.715000  9.090000  42.785000 ;
      RECT  6.485000  42.715000  9.090000  42.785000 ;
      RECT  6.485000  42.785000  9.025000  42.850000 ;
      RECT  6.485000  42.785000  9.025000  42.850000 ;
      RECT  6.490000   4.750000  8.165000   4.820000 ;
      RECT  6.495000  42.850000  9.015000  42.860000 ;
      RECT  6.495000  42.850000  9.015000  42.860000 ;
      RECT  6.505000  42.860000  9.005000  42.870000 ;
      RECT  6.505000  42.860000  9.005000  42.870000 ;
      RECT  6.505000  42.870000  8.935000  42.940000 ;
      RECT  6.505000  42.870000  8.935000  42.940000 ;
      RECT  6.505000  42.940000  8.865000  43.010000 ;
      RECT  6.505000  42.940000  8.865000  43.010000 ;
      RECT  6.505000  43.010000  8.795000  43.080000 ;
      RECT  6.505000  43.010000  8.795000  43.080000 ;
      RECT  6.505000  43.080000  8.725000  43.150000 ;
      RECT  6.505000  43.080000  8.725000  43.150000 ;
      RECT  6.505000  43.150000  8.655000  43.220000 ;
      RECT  6.505000  43.150000  8.655000  43.220000 ;
      RECT  6.505000  43.220000  8.585000  43.290000 ;
      RECT  6.505000  43.220000  8.585000  43.290000 ;
      RECT  6.505000  43.290000  8.515000  43.360000 ;
      RECT  6.505000  43.290000  8.515000  43.360000 ;
      RECT  6.505000  43.360000  8.445000  43.430000 ;
      RECT  6.505000  43.360000  8.445000  43.430000 ;
      RECT  6.505000  43.430000  8.375000  43.500000 ;
      RECT  6.505000  43.430000  8.375000  43.500000 ;
      RECT  6.505000  43.500000  8.305000  43.570000 ;
      RECT  6.505000  43.500000  8.305000  43.570000 ;
      RECT  6.505000  43.570000  8.235000  43.640000 ;
      RECT  6.505000  43.570000  8.235000  43.640000 ;
      RECT  6.505000  43.640000  8.165000  43.710000 ;
      RECT  6.505000  43.640000  8.165000  43.710000 ;
      RECT  6.505000  43.710000  8.095000  43.780000 ;
      RECT  6.505000  43.710000  8.095000  43.780000 ;
      RECT  6.505000  43.780000  8.025000  43.850000 ;
      RECT  6.505000  43.780000  8.025000  43.850000 ;
      RECT  6.505000  43.850000  7.970000  43.905000 ;
      RECT  6.505000  43.850000  7.970000  43.905000 ;
      RECT  6.525000  39.595000 12.240000  39.635000 ;
      RECT  6.525000  39.595000 12.240000  39.635000 ;
      RECT  6.530000   0.000000 12.615000   1.380000 ;
      RECT  6.530000   1.380000 12.615000   3.695000 ;
      RECT  6.540000   8.695000 13.690000   8.765000 ;
      RECT  6.540000   8.695000 13.690000   8.765000 ;
      RECT  6.560000   4.820000  8.165000   4.890000 ;
      RECT  6.595000  39.525000 12.280000  39.595000 ;
      RECT  6.595000  39.525000 12.280000  39.595000 ;
      RECT  6.610000   8.765000 13.690000   8.835000 ;
      RECT  6.610000   8.765000 13.690000   8.835000 ;
      RECT  6.630000   4.890000  8.165000   4.960000 ;
      RECT  6.665000  39.455000 12.350000  39.525000 ;
      RECT  6.665000  39.455000 12.350000  39.525000 ;
      RECT  6.670000   0.000000 12.475000   1.325000 ;
      RECT  6.680000   8.835000 13.690000   8.905000 ;
      RECT  6.680000   8.835000 13.690000   8.905000 ;
      RECT  6.690000   5.215000  8.305000   6.825000 ;
      RECT  6.700000   4.960000  8.165000   5.030000 ;
      RECT  6.735000  39.385000 12.420000  39.455000 ;
      RECT  6.735000  39.385000 12.420000  39.455000 ;
      RECT  6.740000   1.325000 12.475000   1.395000 ;
      RECT  6.740000   1.325000 12.475000   1.395000 ;
      RECT  6.750000   8.905000 13.690000   8.975000 ;
      RECT  6.750000   8.905000 13.690000   8.975000 ;
      RECT  6.770000   5.030000  8.165000   5.100000 ;
      RECT  6.805000  39.315000 12.490000  39.385000 ;
      RECT  6.805000  39.315000 12.490000  39.385000 ;
      RECT  6.810000   1.395000 12.475000   1.465000 ;
      RECT  6.810000   1.395000 12.475000   1.465000 ;
      RECT  6.820000   8.975000 13.690000   9.045000 ;
      RECT  6.820000   8.975000 13.690000   9.045000 ;
      RECT  6.830000   5.100000  8.165000   5.160000 ;
      RECT  6.830000   5.160000  8.165000   6.965000 ;
      RECT  6.875000  39.245000 12.560000  39.315000 ;
      RECT  6.875000  39.245000 12.560000  39.315000 ;
      RECT  6.880000   1.465000 12.475000   1.535000 ;
      RECT  6.880000   1.465000 12.475000   1.535000 ;
      RECT  6.890000   9.045000 13.690000   9.115000 ;
      RECT  6.890000   9.045000 13.690000   9.115000 ;
      RECT  6.945000   9.365000 13.830000  18.285000 ;
      RECT  6.945000  18.285000 15.245000  19.700000 ;
      RECT  6.945000  19.700000 15.245000  31.485000 ;
      RECT  6.945000  31.485000 14.830000  31.900000 ;
      RECT  6.945000  31.900000 14.830000  37.240000 ;
      RECT  6.945000  37.240000 13.095000  38.980000 ;
      RECT  6.945000  38.980000 12.495000  39.580000 ;
      RECT  6.945000  39.175000 12.630000  39.245000 ;
      RECT  6.945000  39.175000 12.630000  39.245000 ;
      RECT  6.950000   1.535000 12.475000   1.605000 ;
      RECT  6.950000   1.535000 12.475000   1.605000 ;
      RECT  6.960000   9.115000 13.690000   9.185000 ;
      RECT  6.960000   9.115000 13.690000   9.185000 ;
      RECT  7.015000  39.105000 12.700000  39.175000 ;
      RECT  7.015000  39.105000 12.700000  39.175000 ;
      RECT  7.020000   1.605000 12.475000   1.675000 ;
      RECT  7.020000   1.605000 12.475000   1.675000 ;
      RECT  7.030000   9.185000 13.690000   9.255000 ;
      RECT  7.030000   9.185000 13.690000   9.255000 ;
      RECT  7.085000   9.255000 13.690000   9.310000 ;
      RECT  7.085000   9.255000 13.690000   9.310000 ;
      RECT  7.085000   9.310000 13.690000  18.340000 ;
      RECT  7.085000  18.340000 13.690000  18.410000 ;
      RECT  7.085000  18.340000 13.690000  18.410000 ;
      RECT  7.085000  18.410000 13.760000  18.480000 ;
      RECT  7.085000  18.410000 13.760000  18.480000 ;
      RECT  7.085000  18.480000 13.830000  18.550000 ;
      RECT  7.085000  18.480000 13.830000  18.550000 ;
      RECT  7.085000  18.550000 13.900000  18.620000 ;
      RECT  7.085000  18.550000 13.900000  18.620000 ;
      RECT  7.085000  18.620000 13.970000  18.690000 ;
      RECT  7.085000  18.620000 13.970000  18.690000 ;
      RECT  7.085000  18.690000 14.040000  18.760000 ;
      RECT  7.085000  18.690000 14.040000  18.760000 ;
      RECT  7.085000  18.760000 14.110000  18.830000 ;
      RECT  7.085000  18.760000 14.110000  18.830000 ;
      RECT  7.085000  18.830000 14.180000  18.900000 ;
      RECT  7.085000  18.830000 14.180000  18.900000 ;
      RECT  7.085000  18.900000 14.250000  18.970000 ;
      RECT  7.085000  18.900000 14.250000  18.970000 ;
      RECT  7.085000  18.970000 14.320000  19.040000 ;
      RECT  7.085000  18.970000 14.320000  19.040000 ;
      RECT  7.085000  19.040000 14.390000  19.110000 ;
      RECT  7.085000  19.040000 14.390000  19.110000 ;
      RECT  7.085000  19.110000 14.460000  19.180000 ;
      RECT  7.085000  19.110000 14.460000  19.180000 ;
      RECT  7.085000  19.180000 14.530000  19.250000 ;
      RECT  7.085000  19.180000 14.530000  19.250000 ;
      RECT  7.085000  19.250000 14.600000  19.320000 ;
      RECT  7.085000  19.250000 14.600000  19.320000 ;
      RECT  7.085000  19.320000 14.670000  19.390000 ;
      RECT  7.085000  19.320000 14.670000  19.390000 ;
      RECT  7.085000  19.390000 14.740000  19.460000 ;
      RECT  7.085000  19.390000 14.740000  19.460000 ;
      RECT  7.085000  19.460000 14.810000  19.530000 ;
      RECT  7.085000  19.460000 14.810000  19.530000 ;
      RECT  7.085000  19.530000 14.880000  19.600000 ;
      RECT  7.085000  19.530000 14.880000  19.600000 ;
      RECT  7.085000  19.600000 14.950000  19.670000 ;
      RECT  7.085000  19.600000 14.950000  19.670000 ;
      RECT  7.085000  19.670000 15.020000  19.740000 ;
      RECT  7.085000  19.670000 15.020000  19.740000 ;
      RECT  7.085000  19.740000 15.090000  19.755000 ;
      RECT  7.085000  19.740000 15.090000  19.755000 ;
      RECT  7.085000  19.755000 15.105000  31.430000 ;
      RECT  7.085000  31.430000 15.035000  31.500000 ;
      RECT  7.085000  31.430000 15.035000  31.500000 ;
      RECT  7.085000  31.500000 14.965000  31.570000 ;
      RECT  7.085000  31.500000 14.965000  31.570000 ;
      RECT  7.085000  31.570000 14.895000  31.640000 ;
      RECT  7.085000  31.570000 14.895000  31.640000 ;
      RECT  7.085000  31.640000 14.825000  31.710000 ;
      RECT  7.085000  31.640000 14.825000  31.710000 ;
      RECT  7.085000  31.710000 14.755000  31.780000 ;
      RECT  7.085000  31.710000 14.755000  31.780000 ;
      RECT  7.085000  31.780000 14.690000  31.845000 ;
      RECT  7.085000  31.780000 14.690000  31.845000 ;
      RECT  7.085000  31.845000 14.690000  37.185000 ;
      RECT  7.085000  37.185000 14.620000  37.255000 ;
      RECT  7.085000  37.185000 14.620000  37.255000 ;
      RECT  7.085000  37.255000 14.550000  37.325000 ;
      RECT  7.085000  37.255000 14.550000  37.325000 ;
      RECT  7.085000  37.325000 14.480000  37.395000 ;
      RECT  7.085000  37.325000 14.480000  37.395000 ;
      RECT  7.085000  37.395000 14.410000  37.465000 ;
      RECT  7.085000  37.395000 14.410000  37.465000 ;
      RECT  7.085000  37.465000 14.340000  37.535000 ;
      RECT  7.085000  37.465000 14.340000  37.535000 ;
      RECT  7.085000  37.535000 14.270000  37.605000 ;
      RECT  7.085000  37.535000 14.270000  37.605000 ;
      RECT  7.085000  37.605000 14.200000  37.675000 ;
      RECT  7.085000  37.605000 14.200000  37.675000 ;
      RECT  7.085000  37.675000 14.130000  37.745000 ;
      RECT  7.085000  37.675000 14.130000  37.745000 ;
      RECT  7.085000  37.745000 14.060000  37.815000 ;
      RECT  7.085000  37.745000 14.060000  37.815000 ;
      RECT  7.085000  37.815000 13.990000  37.885000 ;
      RECT  7.085000  37.815000 13.990000  37.885000 ;
      RECT  7.085000  37.885000 13.920000  37.955000 ;
      RECT  7.085000  37.885000 13.920000  37.955000 ;
      RECT  7.085000  37.955000 13.850000  38.025000 ;
      RECT  7.085000  37.955000 13.850000  38.025000 ;
      RECT  7.085000  38.025000 13.780000  38.095000 ;
      RECT  7.085000  38.025000 13.780000  38.095000 ;
      RECT  7.085000  38.095000 13.710000  38.165000 ;
      RECT  7.085000  38.095000 13.710000  38.165000 ;
      RECT  7.085000  38.165000 13.640000  38.235000 ;
      RECT  7.085000  38.165000 13.640000  38.235000 ;
      RECT  7.085000  38.235000 13.570000  38.305000 ;
      RECT  7.085000  38.235000 13.570000  38.305000 ;
      RECT  7.085000  38.305000 13.500000  38.375000 ;
      RECT  7.085000  38.305000 13.500000  38.375000 ;
      RECT  7.085000  38.375000 13.430000  38.445000 ;
      RECT  7.085000  38.375000 13.430000  38.445000 ;
      RECT  7.085000  38.445000 13.360000  38.515000 ;
      RECT  7.085000  38.445000 13.360000  38.515000 ;
      RECT  7.085000  38.515000 13.290000  38.585000 ;
      RECT  7.085000  38.515000 13.290000  38.585000 ;
      RECT  7.085000  38.585000 13.220000  38.655000 ;
      RECT  7.085000  38.585000 13.220000  38.655000 ;
      RECT  7.085000  38.655000 13.150000  38.725000 ;
      RECT  7.085000  38.655000 13.150000  38.725000 ;
      RECT  7.085000  38.725000 13.080000  38.795000 ;
      RECT  7.085000  38.725000 13.080000  38.795000 ;
      RECT  7.085000  38.795000 13.010000  38.865000 ;
      RECT  7.085000  38.795000 13.010000  38.865000 ;
      RECT  7.085000  38.865000 12.940000  38.935000 ;
      RECT  7.085000  38.865000 12.940000  38.935000 ;
      RECT  7.085000  38.935000 12.870000  39.005000 ;
      RECT  7.085000  38.935000 12.870000  39.005000 ;
      RECT  7.085000  39.005000 12.840000  39.035000 ;
      RECT  7.085000  39.005000 12.840000  39.035000 ;
      RECT  7.085000  39.035000 12.770000  39.105000 ;
      RECT  7.085000  39.035000 12.770000  39.105000 ;
      RECT  7.090000   1.675000 12.475000   1.745000 ;
      RECT  7.090000   1.675000 12.475000   1.745000 ;
      RECT  7.160000   1.745000 12.475000   1.815000 ;
      RECT  7.160000   1.745000 12.475000   1.815000 ;
      RECT  7.230000   1.815000 12.475000   1.885000 ;
      RECT  7.230000   1.815000 12.475000   1.885000 ;
      RECT  7.300000   1.885000 12.475000   1.955000 ;
      RECT  7.300000   1.885000 12.475000   1.955000 ;
      RECT  7.370000   1.955000 12.475000   2.025000 ;
      RECT  7.370000   1.955000 12.475000   2.025000 ;
      RECT  7.440000   2.025000 12.475000   2.095000 ;
      RECT  7.440000   2.025000 12.475000   2.095000 ;
      RECT  7.510000   2.095000 12.475000   2.165000 ;
      RECT  7.510000   2.095000 12.475000   2.165000 ;
      RECT  7.580000   2.165000 12.475000   2.235000 ;
      RECT  7.580000   2.165000 12.475000   2.235000 ;
      RECT  7.650000   2.235000 12.475000   2.305000 ;
      RECT  7.650000   2.235000 12.475000   2.305000 ;
      RECT  7.715000  56.630000 14.210000  57.835000 ;
      RECT  7.715000  57.835000 14.055000  57.990000 ;
      RECT  7.715000  57.990000 14.055000  58.450000 ;
      RECT  7.715000  58.450000 76.775000  73.555000 ;
      RECT  7.715000  73.555000 76.775000  74.045000 ;
      RECT  7.720000   2.305000 12.475000   2.375000 ;
      RECT  7.720000   2.305000 12.475000   2.375000 ;
      RECT  7.790000   2.375000 12.475000   2.445000 ;
      RECT  7.790000   2.375000 12.475000   2.445000 ;
      RECT  7.855000  56.685000 14.070000  57.780000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 14.000000  57.850000 ;
      RECT  7.855000  57.780000 14.000000  57.850000 ;
      RECT  7.855000  57.850000 13.930000  57.920000 ;
      RECT  7.855000  57.850000 13.930000  57.920000 ;
      RECT  7.855000  57.920000 13.915000  57.935000 ;
      RECT  7.855000  57.920000 13.915000  57.935000 ;
      RECT  7.855000  57.935000 13.915000  58.590000 ;
      RECT  7.855000  58.590000 76.635000  73.500000 ;
      RECT  7.860000   2.445000 12.475000   2.515000 ;
      RECT  7.860000   2.445000 12.475000   2.515000 ;
      RECT  7.885000  56.655000 14.070000  56.685000 ;
      RECT  7.885000  56.655000 14.070000  56.685000 ;
      RECT  7.925000  73.500000 76.635000  73.570000 ;
      RECT  7.925000  73.500000 76.635000  73.570000 ;
      RECT  7.930000   2.515000 12.475000   2.585000 ;
      RECT  7.930000   2.515000 12.475000   2.585000 ;
      RECT  7.955000  56.585000 14.070000  56.655000 ;
      RECT  7.955000  56.585000 14.070000  56.655000 ;
      RECT  7.995000  73.570000 76.635000  73.640000 ;
      RECT  7.995000  73.570000 76.635000  73.640000 ;
      RECT  8.000000   2.585000 12.475000   2.655000 ;
      RECT  8.000000   2.585000 12.475000   2.655000 ;
      RECT  8.025000  56.515000 14.070000  56.585000 ;
      RECT  8.025000  56.515000 14.070000  56.585000 ;
      RECT  8.065000  73.640000 76.635000  73.710000 ;
      RECT  8.065000  73.640000 76.635000  73.710000 ;
      RECT  8.070000   2.655000 12.475000   2.725000 ;
      RECT  8.070000   2.655000 12.475000   2.725000 ;
      RECT  8.095000  56.445000 14.070000  56.515000 ;
      RECT  8.095000  56.445000 14.070000  56.515000 ;
      RECT  8.135000  73.710000 76.635000  73.780000 ;
      RECT  8.135000  73.710000 76.635000  73.780000 ;
      RECT  8.140000   2.725000 12.475000   2.795000 ;
      RECT  8.140000   2.725000 12.475000   2.795000 ;
      RECT  8.165000  56.375000 14.070000  56.445000 ;
      RECT  8.165000  56.375000 14.070000  56.445000 ;
      RECT  8.205000  73.780000 76.635000  73.850000 ;
      RECT  8.205000  73.780000 76.635000  73.850000 ;
      RECT  8.205000  74.045000 76.775000  74.620000 ;
      RECT  8.205000  74.620000 76.775000  75.025000 ;
      RECT  8.210000   2.795000 12.475000   2.865000 ;
      RECT  8.210000   2.795000 12.475000   2.865000 ;
      RECT  8.235000  56.305000 14.070000  56.375000 ;
      RECT  8.235000  56.305000 14.070000  56.375000 ;
      RECT  8.275000  73.850000 76.635000  73.920000 ;
      RECT  8.275000  73.850000 76.635000  73.920000 ;
      RECT  8.280000   2.865000 12.475000   2.935000 ;
      RECT  8.280000   2.865000 12.475000   2.935000 ;
      RECT  8.305000  56.235000 14.070000  56.305000 ;
      RECT  8.305000  56.235000 14.070000  56.305000 ;
      RECT  8.345000  73.920000 76.635000  73.990000 ;
      RECT  8.345000  73.920000 76.635000  73.990000 ;
      RECT  8.345000  73.990000 76.635000  74.565000 ;
      RECT  8.350000   2.935000 12.475000   3.005000 ;
      RECT  8.350000   2.935000 12.475000   3.005000 ;
      RECT  8.375000  54.130000 14.210000  55.970000 ;
      RECT  8.375000  55.970000 14.210000  56.630000 ;
      RECT  8.375000  56.165000 14.070000  56.235000 ;
      RECT  8.375000  56.165000 14.070000  56.235000 ;
      RECT  8.415000  74.565000 76.635000  74.635000 ;
      RECT  8.415000  74.565000 76.635000  74.635000 ;
      RECT  8.420000   3.005000 12.475000   3.075000 ;
      RECT  8.420000   3.005000 12.475000   3.075000 ;
      RECT  8.445000  56.095000 14.070000  56.165000 ;
      RECT  8.445000  56.095000 14.070000  56.165000 ;
      RECT  8.485000  74.635000 76.635000  74.705000 ;
      RECT  8.485000  74.635000 76.635000  74.705000 ;
      RECT  8.490000   3.075000 12.475000   3.145000 ;
      RECT  8.490000   3.075000 12.475000   3.145000 ;
      RECT  8.515000  54.185000 14.070000  56.025000 ;
      RECT  8.515000  56.025000 14.070000  56.095000 ;
      RECT  8.515000  56.025000 14.070000  56.095000 ;
      RECT  8.525000  54.175000 14.070000  54.185000 ;
      RECT  8.525000  54.175000 14.070000  54.185000 ;
      RECT  8.555000  74.705000 76.635000  74.775000 ;
      RECT  8.555000  74.705000 76.635000  74.775000 ;
      RECT  8.560000   3.145000 12.475000   3.215000 ;
      RECT  8.560000   3.145000 12.475000   3.215000 ;
      RECT  8.595000  44.245000 11.110000  47.445000 ;
      RECT  8.595000  47.445000 11.880000  48.215000 ;
      RECT  8.595000  48.215000 14.210000  48.745000 ;
      RECT  8.595000  48.745000 14.210000  53.910000 ;
      RECT  8.595000  53.910000 14.210000  54.130000 ;
      RECT  8.595000  54.105000 14.070000  54.175000 ;
      RECT  8.595000  54.105000 14.070000  54.175000 ;
      RECT  8.610000  75.025000 76.775000  77.135000 ;
      RECT  8.610000  77.135000 76.775000  77.225000 ;
      RECT  8.625000  74.775000 76.635000  74.845000 ;
      RECT  8.625000  74.775000 76.635000  74.845000 ;
      RECT  8.630000   3.215000 12.475000   3.285000 ;
      RECT  8.630000   3.215000 12.475000   3.285000 ;
      RECT  8.665000  54.035000 14.070000  54.105000 ;
      RECT  8.665000  54.035000 14.070000  54.105000 ;
      RECT  8.695000  74.845000 76.635000  74.915000 ;
      RECT  8.695000  74.845000 76.635000  74.915000 ;
      RECT  8.700000   3.285000 12.475000   3.355000 ;
      RECT  8.700000   3.285000 12.475000   3.355000 ;
      RECT  8.700000  77.225000 76.775000  77.685000 ;
      RECT  8.735000  44.300000 10.970000  45.265000 ;
      RECT  8.735000  45.335000  8.805000  45.405000 ;
      RECT  8.735000  45.335000  8.805000  45.405000 ;
      RECT  8.735000  45.405000  8.875000  45.475000 ;
      RECT  8.735000  45.405000  8.875000  45.475000 ;
      RECT  8.735000  45.475000  8.945000  45.545000 ;
      RECT  8.735000  45.475000  8.945000  45.545000 ;
      RECT  8.735000  45.545000  9.015000  45.615000 ;
      RECT  8.735000  45.545000  9.015000  45.615000 ;
      RECT  8.735000  45.615000  9.085000  45.685000 ;
      RECT  8.735000  45.615000  9.085000  45.685000 ;
      RECT  8.735000  45.685000  9.155000  45.755000 ;
      RECT  8.735000  45.685000  9.155000  45.755000 ;
      RECT  8.735000  45.755000  9.225000  45.825000 ;
      RECT  8.735000  45.755000  9.225000  45.825000 ;
      RECT  8.735000  45.825000  9.295000  45.895000 ;
      RECT  8.735000  45.825000  9.295000  45.895000 ;
      RECT  8.735000  45.895000  9.365000  45.965000 ;
      RECT  8.735000  45.895000  9.365000  45.965000 ;
      RECT  8.735000  45.965000  9.435000  46.035000 ;
      RECT  8.735000  45.965000  9.435000  46.035000 ;
      RECT  8.735000  46.035000  9.505000  46.105000 ;
      RECT  8.735000  46.035000  9.505000  46.105000 ;
      RECT  8.735000  46.105000  9.575000  46.175000 ;
      RECT  8.735000  46.105000  9.575000  46.175000 ;
      RECT  8.735000  46.175000  9.645000  46.245000 ;
      RECT  8.735000  46.175000  9.645000  46.245000 ;
      RECT  8.735000  46.245000  9.715000  46.315000 ;
      RECT  8.735000  46.245000  9.715000  46.315000 ;
      RECT  8.735000  46.315000  9.785000  46.385000 ;
      RECT  8.735000  46.315000  9.785000  46.385000 ;
      RECT  8.735000  46.385000  9.855000  46.455000 ;
      RECT  8.735000  46.385000  9.855000  46.455000 ;
      RECT  8.735000  46.455000  9.925000  46.525000 ;
      RECT  8.735000  46.455000  9.925000  46.525000 ;
      RECT  8.735000  46.525000  9.995000  46.595000 ;
      RECT  8.735000  46.525000  9.995000  46.595000 ;
      RECT  8.735000  46.595000 10.065000  46.665000 ;
      RECT  8.735000  46.595000 10.065000  46.665000 ;
      RECT  8.735000  46.665000 10.135000  46.735000 ;
      RECT  8.735000  46.665000 10.135000  46.735000 ;
      RECT  8.735000  46.735000 10.205000  46.805000 ;
      RECT  8.735000  46.735000 10.205000  46.805000 ;
      RECT  8.735000  46.805000 10.275000  46.875000 ;
      RECT  8.735000  46.805000 10.275000  46.875000 ;
      RECT  8.735000  46.875000 10.345000  46.945000 ;
      RECT  8.735000  46.875000 10.345000  46.945000 ;
      RECT  8.735000  46.945000 10.415000  47.015000 ;
      RECT  8.735000  46.945000 10.415000  47.015000 ;
      RECT  8.735000  47.015000 10.485000  47.085000 ;
      RECT  8.735000  47.015000 10.485000  47.085000 ;
      RECT  8.735000  47.085000 10.555000  47.155000 ;
      RECT  8.735000  47.085000 10.555000  47.155000 ;
      RECT  8.735000  47.155000 10.625000  47.225000 ;
      RECT  8.735000  47.155000 10.625000  47.225000 ;
      RECT  8.735000  47.225000 10.695000  47.295000 ;
      RECT  8.735000  47.225000 10.695000  47.295000 ;
      RECT  8.735000  47.295000 10.765000  47.365000 ;
      RECT  8.735000  47.295000 10.765000  47.365000 ;
      RECT  8.735000  47.365000 10.835000  47.435000 ;
      RECT  8.735000  47.365000 10.835000  47.435000 ;
      RECT  8.735000  47.435000 10.905000  47.500000 ;
      RECT  8.735000  47.435000 10.905000  47.500000 ;
      RECT  8.735000  47.500000 10.970000  47.570000 ;
      RECT  8.735000  47.500000 10.970000  47.570000 ;
      RECT  8.735000  47.570000 11.040000  47.640000 ;
      RECT  8.735000  47.570000 11.040000  47.640000 ;
      RECT  8.735000  47.640000 11.110000  47.710000 ;
      RECT  8.735000  47.640000 11.110000  47.710000 ;
      RECT  8.735000  47.710000 11.180000  47.780000 ;
      RECT  8.735000  47.710000 11.180000  47.780000 ;
      RECT  8.735000  47.780000 11.250000  47.850000 ;
      RECT  8.735000  47.780000 11.250000  47.850000 ;
      RECT  8.735000  47.850000 11.320000  47.920000 ;
      RECT  8.735000  47.850000 11.320000  47.920000 ;
      RECT  8.735000  47.920000 11.390000  47.990000 ;
      RECT  8.735000  47.920000 11.390000  47.990000 ;
      RECT  8.735000  47.990000 11.460000  48.060000 ;
      RECT  8.735000  47.990000 11.460000  48.060000 ;
      RECT  8.735000  48.060000 11.530000  48.130000 ;
      RECT  8.735000  48.060000 11.530000  48.130000 ;
      RECT  8.735000  48.130000 11.600000  48.200000 ;
      RECT  8.735000  48.130000 11.600000  48.200000 ;
      RECT  8.735000  48.200000 11.670000  48.270000 ;
      RECT  8.735000  48.200000 11.670000  48.270000 ;
      RECT  8.735000  48.270000 11.740000  48.340000 ;
      RECT  8.735000  48.270000 11.740000  48.340000 ;
      RECT  8.735000  48.340000 11.810000  48.355000 ;
      RECT  8.735000  48.340000 11.810000  48.355000 ;
      RECT  8.735000  48.355000 13.625000  48.425000 ;
      RECT  8.735000  48.355000 13.625000  48.425000 ;
      RECT  8.735000  48.425000 13.695000  48.495000 ;
      RECT  8.735000  48.425000 13.695000  48.495000 ;
      RECT  8.735000  48.495000 13.765000  48.565000 ;
      RECT  8.735000  48.495000 13.765000  48.565000 ;
      RECT  8.735000  48.565000 13.835000  48.635000 ;
      RECT  8.735000  48.565000 13.835000  48.635000 ;
      RECT  8.735000  48.635000 13.905000  48.705000 ;
      RECT  8.735000  48.635000 13.905000  48.705000 ;
      RECT  8.735000  48.705000 13.975000  48.775000 ;
      RECT  8.735000  48.705000 13.975000  48.775000 ;
      RECT  8.735000  48.775000 14.045000  48.800000 ;
      RECT  8.735000  48.775000 14.045000  48.800000 ;
      RECT  8.735000  48.800000 14.070000  53.965000 ;
      RECT  8.735000  48.800000 14.070000  56.025000 ;
      RECT  8.735000  48.800000 14.070000  56.685000 ;
      RECT  8.735000  48.800000 14.070000  56.685000 ;
      RECT  8.735000  48.800000 14.070000  56.685000 ;
      RECT  8.735000  48.800000 14.070000  56.685000 ;
      RECT  8.735000  53.965000 14.070000  54.035000 ;
      RECT  8.735000  53.965000 14.070000  54.035000 ;
      RECT  8.750000  74.915000 76.635000  74.970000 ;
      RECT  8.750000  74.915000 76.635000  74.970000 ;
      RECT  8.750000  74.970000 76.635000  77.080000 ;
      RECT  8.755000  44.280000 10.970000  44.300000 ;
      RECT  8.770000   3.355000 12.475000   3.425000 ;
      RECT  8.770000   3.355000 12.475000   3.425000 ;
      RECT  8.795000  77.080000 76.635000  77.125000 ;
      RECT  8.795000  77.080000 76.635000  77.125000 ;
      RECT  8.825000  44.210000 10.970000  44.280000 ;
      RECT  8.840000   3.425000 12.475000   3.495000 ;
      RECT  8.840000   3.425000 12.475000   3.495000 ;
      RECT  8.840000  74.970000 76.635000  96.080000 ;
      RECT  8.840000  74.970000 76.635000  96.080000 ;
      RECT  8.840000  77.125000 76.635000  77.170000 ;
      RECT  8.840000  77.125000 76.635000  77.170000 ;
      RECT  8.845000   3.695000 12.615000   5.410000 ;
      RECT  8.845000   5.410000 13.830000   6.625000 ;
      RECT  8.845000   6.625000 13.830000   6.920000 ;
      RECT  8.895000  44.140000 10.970000  44.210000 ;
      RECT  8.910000   3.495000 12.475000   3.565000 ;
      RECT  8.910000   3.495000 12.475000   3.565000 ;
      RECT  8.965000  44.070000 10.970000  44.140000 ;
      RECT  8.980000   3.565000 12.475000   3.635000 ;
      RECT  8.980000   3.565000 12.475000   3.635000 ;
      RECT  8.985000   1.325000 12.475000   5.465000 ;
      RECT  8.985000   1.325000 12.475000   5.465000 ;
      RECT  8.985000   1.325000 12.475000   5.465000 ;
      RECT  8.985000   1.325000 12.475000   5.465000 ;
      RECT  8.985000   3.635000 12.475000   3.640000 ;
      RECT  8.985000   3.635000 12.475000   3.640000 ;
      RECT  8.985000   5.465000 12.475000   5.535000 ;
      RECT  8.985000   5.465000 12.475000   5.535000 ;
      RECT  8.985000   5.535000 12.545000   5.605000 ;
      RECT  8.985000   5.535000 12.545000   5.605000 ;
      RECT  8.985000   5.605000 12.615000   5.675000 ;
      RECT  8.985000   5.605000 12.615000   5.675000 ;
      RECT  8.985000   5.675000 12.685000   5.745000 ;
      RECT  8.985000   5.675000 12.685000   5.745000 ;
      RECT  8.985000   5.745000 12.755000   5.815000 ;
      RECT  8.985000   5.745000 12.755000   5.815000 ;
      RECT  8.985000   5.815000 12.825000   5.885000 ;
      RECT  8.985000   5.815000 12.825000   5.885000 ;
      RECT  8.985000   5.885000 12.895000   5.955000 ;
      RECT  8.985000   5.885000 12.895000   5.955000 ;
      RECT  8.985000   5.955000 12.965000   6.025000 ;
      RECT  8.985000   5.955000 12.965000   6.025000 ;
      RECT  8.985000   6.025000 13.035000   6.095000 ;
      RECT  8.985000   6.025000 13.035000   6.095000 ;
      RECT  8.985000   6.095000 13.105000   6.165000 ;
      RECT  8.985000   6.095000 13.105000   6.165000 ;
      RECT  8.985000   6.165000 13.175000   6.235000 ;
      RECT  8.985000   6.165000 13.175000   6.235000 ;
      RECT  8.985000   6.235000 13.245000   6.305000 ;
      RECT  8.985000   6.235000 13.245000   6.305000 ;
      RECT  8.985000   6.305000 13.315000   6.375000 ;
      RECT  8.985000   6.305000 13.315000   6.375000 ;
      RECT  8.985000   6.375000 13.385000   6.445000 ;
      RECT  8.985000   6.375000 13.385000   6.445000 ;
      RECT  8.985000   6.445000 13.455000   6.515000 ;
      RECT  8.985000   6.445000 13.455000   6.515000 ;
      RECT  8.985000   6.515000 13.525000   6.585000 ;
      RECT  8.985000   6.515000 13.525000   6.585000 ;
      RECT  8.985000   6.585000 13.595000   6.655000 ;
      RECT  8.985000   6.585000 13.595000   6.655000 ;
      RECT  8.985000   6.655000 13.665000   6.680000 ;
      RECT  8.985000   6.655000 13.665000   6.680000 ;
      RECT  8.985000   6.680000 13.690000   7.060000 ;
      RECT  9.035000  44.000000 10.970000  44.070000 ;
      RECT  9.060000  43.775000 11.110000  44.245000 ;
      RECT  9.105000  43.930000 10.970000  44.000000 ;
      RECT  9.175000  43.860000 10.970000  43.930000 ;
      RECT  9.245000  43.790000 10.970000  43.860000 ;
      RECT  9.315000  43.720000 10.970000  43.790000 ;
      RECT  9.375000  43.660000 10.970000  43.720000 ;
      RECT  9.445000  43.590000 11.030000  43.660000 ;
      RECT  9.515000  43.520000 11.100000  43.590000 ;
      RECT  9.585000  43.450000 11.170000  43.520000 ;
      RECT  9.655000  43.380000 11.240000  43.450000 ;
      RECT  9.725000  43.310000 11.310000  43.380000 ;
      RECT  9.795000  43.240000 11.380000  43.310000 ;
      RECT  9.865000  43.170000 11.450000  43.240000 ;
      RECT  9.935000  43.100000 11.520000  43.170000 ;
      RECT 10.005000  43.030000 11.590000  43.100000 ;
      RECT 10.075000  42.960000 11.660000  43.030000 ;
      RECT 10.145000  42.890000 11.730000  42.960000 ;
      RECT 10.215000  42.820000 11.800000  42.890000 ;
      RECT 10.285000  42.750000 11.870000  42.820000 ;
      RECT 10.355000  42.680000 11.940000  42.750000 ;
      RECT 10.425000  42.610000 12.010000  42.680000 ;
      RECT 10.495000  42.540000 12.080000  42.610000 ;
      RECT 10.565000  42.470000 12.150000  42.540000 ;
      RECT 10.635000  42.400000 12.220000  42.470000 ;
      RECT 10.705000  42.330000 12.290000  42.400000 ;
      RECT 10.775000  42.260000 12.360000  42.330000 ;
      RECT 10.845000  42.190000 12.430000  42.260000 ;
      RECT 10.915000  42.120000 12.500000  42.190000 ;
      RECT 10.985000  42.050000 12.570000  42.120000 ;
      RECT 11.055000  41.980000 12.640000  42.050000 ;
      RECT 11.125000  41.910000 12.710000  41.980000 ;
      RECT 11.195000  41.840000 12.780000  41.910000 ;
      RECT 11.265000  41.770000 12.850000  41.840000 ;
      RECT 11.335000  41.700000 12.920000  41.770000 ;
      RECT 11.405000  41.630000 12.990000  41.700000 ;
      RECT 11.475000  41.560000 13.060000  41.630000 ;
      RECT 11.545000  41.490000 13.130000  41.560000 ;
      RECT 11.615000  41.420000 13.200000  41.490000 ;
      RECT 11.650000  44.005000 29.985000  47.215000 ;
      RECT 11.650000  47.215000 29.985000  47.675000 ;
      RECT 11.685000  41.350000 13.270000  41.420000 ;
      RECT 11.740000  41.295000 13.340000  41.350000 ;
      RECT 11.790000  44.060000 29.845000  47.160000 ;
      RECT 11.810000  41.225000 13.340000  41.295000 ;
      RECT 11.850000  44.000000 29.845000  44.060000 ;
      RECT 11.850000  44.000000 29.845000  44.060000 ;
      RECT 11.860000  47.160000 29.845000  47.230000 ;
      RECT 11.860000  47.160000 29.845000  47.230000 ;
      RECT 11.880000  41.155000 13.340000  41.225000 ;
      RECT 11.920000  43.930000 29.845000  44.000000 ;
      RECT 11.920000  43.930000 29.845000  44.000000 ;
      RECT 11.930000  47.230000 29.845000  47.300000 ;
      RECT 11.930000  47.230000 29.845000  47.300000 ;
      RECT 11.950000  41.085000 13.340000  41.155000 ;
      RECT 11.990000  43.860000 29.845000  43.930000 ;
      RECT 11.990000  43.860000 29.845000  43.930000 ;
      RECT 12.000000  47.300000 29.845000  47.370000 ;
      RECT 12.000000  47.300000 29.845000  47.370000 ;
      RECT 12.020000  41.015000 13.340000  41.085000 ;
      RECT 12.060000  43.790000 29.845000  43.860000 ;
      RECT 12.060000  43.790000 29.845000  43.860000 ;
      RECT 12.070000  47.370000 29.845000  47.440000 ;
      RECT 12.070000  47.370000 29.845000  47.440000 ;
      RECT 12.090000  40.945000 13.340000  41.015000 ;
      RECT 12.130000  43.720000 29.845000  43.790000 ;
      RECT 12.130000  43.720000 29.845000  43.790000 ;
      RECT 12.140000  47.440000 29.845000  47.510000 ;
      RECT 12.140000  47.440000 29.845000  47.510000 ;
      RECT 12.160000  40.875000 13.340000  40.945000 ;
      RECT 12.165000  47.510000 29.845000  47.535000 ;
      RECT 12.165000  47.510000 29.845000  47.535000 ;
      RECT 12.200000  43.650000 29.845000  43.720000 ;
      RECT 12.200000  43.650000 29.845000  43.720000 ;
      RECT 12.230000  40.805000 13.340000  40.875000 ;
      RECT 12.270000  43.580000 29.845000  43.650000 ;
      RECT 12.270000  43.580000 29.845000  43.650000 ;
      RECT 12.300000  40.735000 13.340000  40.805000 ;
      RECT 12.340000  43.510000 29.845000  43.580000 ;
      RECT 12.340000  43.510000 29.845000  43.580000 ;
      RECT 12.370000  40.665000 13.340000  40.735000 ;
      RECT 12.410000  43.440000 29.845000  43.510000 ;
      RECT 12.410000  43.440000 29.845000  43.510000 ;
      RECT 12.440000  40.595000 13.340000  40.665000 ;
      RECT 12.465000  40.370000 13.480000  41.405000 ;
      RECT 12.480000  43.370000 29.845000  43.440000 ;
      RECT 12.480000  43.370000 29.845000  43.440000 ;
      RECT 12.510000  40.525000 13.340000  40.595000 ;
      RECT 12.550000  43.300000 29.845000  43.370000 ;
      RECT 12.550000  43.300000 29.845000  43.370000 ;
      RECT 12.580000  40.455000 13.340000  40.525000 ;
      RECT 12.620000  43.230000 29.845000  43.300000 ;
      RECT 12.620000  43.230000 29.845000  43.300000 ;
      RECT 12.650000  40.385000 13.340000  40.455000 ;
      RECT 12.690000  43.160000 29.845000  43.230000 ;
      RECT 12.690000  43.160000 29.845000  43.230000 ;
      RECT 12.720000  40.315000 13.340000  40.385000 ;
      RECT 12.745000  40.290000 13.340000  40.315000 ;
      RECT 12.760000  43.090000 29.845000  43.160000 ;
      RECT 12.760000  43.090000 29.845000  43.160000 ;
      RECT 12.815000  40.220000 13.365000  40.290000 ;
      RECT 12.830000  43.020000 29.845000  43.090000 ;
      RECT 12.830000  43.020000 29.845000  43.090000 ;
      RECT 12.885000  40.150000 13.435000  40.220000 ;
      RECT 12.900000  42.950000 29.845000  43.020000 ;
      RECT 12.900000  42.950000 29.845000  43.020000 ;
      RECT 12.955000  40.080000 13.505000  40.150000 ;
      RECT 12.970000  42.880000 29.845000  42.950000 ;
      RECT 12.970000  42.880000 29.845000  42.950000 ;
      RECT 13.025000  40.010000 13.575000  40.080000 ;
      RECT 13.040000  42.810000 29.845000  42.880000 ;
      RECT 13.040000  42.810000 29.845000  42.880000 ;
      RECT 13.095000  39.940000 13.645000  40.010000 ;
      RECT 13.110000  42.740000 29.845000  42.810000 ;
      RECT 13.110000  42.740000 29.845000  42.810000 ;
      RECT 13.155000   0.000000 16.170000   2.380000 ;
      RECT 13.155000   2.380000 16.955000   3.160000 ;
      RECT 13.155000   3.160000 16.955000   5.180000 ;
      RECT 13.155000   5.180000 16.955000   6.395000 ;
      RECT 13.165000  39.870000 13.715000  39.940000 ;
      RECT 13.180000  42.670000 29.845000  42.740000 ;
      RECT 13.180000  42.670000 29.845000  42.740000 ;
      RECT 13.235000  39.800000 13.785000  39.870000 ;
      RECT 13.250000  42.600000 29.845000  42.670000 ;
      RECT 13.250000  42.600000 29.845000  42.670000 ;
      RECT 13.295000   0.000000 13.595000   0.070000 ;
      RECT 13.295000   0.000000 13.595000   0.070000 ;
      RECT 13.295000   0.070000 13.665000   0.140000 ;
      RECT 13.295000   0.070000 13.665000   0.140000 ;
      RECT 13.295000   0.140000 13.735000   0.210000 ;
      RECT 13.295000   0.140000 13.735000   0.210000 ;
      RECT 13.295000   0.210000 13.805000   0.280000 ;
      RECT 13.295000   0.210000 13.805000   0.280000 ;
      RECT 13.295000   0.280000 13.875000   0.350000 ;
      RECT 13.295000   0.280000 13.875000   0.350000 ;
      RECT 13.295000   0.350000 13.945000   0.420000 ;
      RECT 13.295000   0.350000 13.945000   0.420000 ;
      RECT 13.295000   0.420000 14.015000   0.490000 ;
      RECT 13.295000   0.420000 14.015000   0.490000 ;
      RECT 13.295000   0.490000 14.085000   0.560000 ;
      RECT 13.295000   0.490000 14.085000   0.560000 ;
      RECT 13.295000   0.560000 14.155000   0.630000 ;
      RECT 13.295000   0.560000 14.155000   0.630000 ;
      RECT 13.295000   0.630000 14.225000   0.700000 ;
      RECT 13.295000   0.630000 14.225000   0.700000 ;
      RECT 13.295000   0.700000 14.295000   0.770000 ;
      RECT 13.295000   0.700000 14.295000   0.770000 ;
      RECT 13.295000   0.770000 14.365000   0.840000 ;
      RECT 13.295000   0.770000 14.365000   0.840000 ;
      RECT 13.295000   0.840000 14.435000   0.910000 ;
      RECT 13.295000   0.840000 14.435000   0.910000 ;
      RECT 13.295000   0.910000 14.505000   0.980000 ;
      RECT 13.295000   0.910000 14.505000   0.980000 ;
      RECT 13.295000   0.980000 14.575000   1.050000 ;
      RECT 13.295000   0.980000 14.575000   1.050000 ;
      RECT 13.295000   1.050000 14.645000   1.120000 ;
      RECT 13.295000   1.050000 14.645000   1.120000 ;
      RECT 13.295000   1.120000 14.715000   1.190000 ;
      RECT 13.295000   1.120000 14.715000   1.190000 ;
      RECT 13.295000   1.190000 14.785000   1.260000 ;
      RECT 13.295000   1.190000 14.785000   1.260000 ;
      RECT 13.295000   1.260000 14.855000   1.330000 ;
      RECT 13.295000   1.260000 14.855000   1.330000 ;
      RECT 13.295000   1.330000 14.925000   1.400000 ;
      RECT 13.295000   1.330000 14.925000   1.400000 ;
      RECT 13.295000   1.400000 14.995000   1.470000 ;
      RECT 13.295000   1.400000 14.995000   1.470000 ;
      RECT 13.295000   1.470000 15.065000   1.540000 ;
      RECT 13.295000   1.470000 15.065000   1.540000 ;
      RECT 13.295000   1.540000 15.135000   1.610000 ;
      RECT 13.295000   1.540000 15.135000   1.610000 ;
      RECT 13.295000   1.610000 15.205000   1.680000 ;
      RECT 13.295000   1.610000 15.205000   1.680000 ;
      RECT 13.295000   1.680000 15.275000   1.750000 ;
      RECT 13.295000   1.680000 15.275000   1.750000 ;
      RECT 13.295000   1.750000 15.345000   1.820000 ;
      RECT 13.295000   1.750000 15.345000   1.820000 ;
      RECT 13.295000   1.820000 15.415000   1.890000 ;
      RECT 13.295000   1.820000 15.415000   1.890000 ;
      RECT 13.295000   1.890000 15.485000   1.960000 ;
      RECT 13.295000   1.890000 15.485000   1.960000 ;
      RECT 13.295000   1.960000 15.555000   2.030000 ;
      RECT 13.295000   1.960000 15.555000   2.030000 ;
      RECT 13.295000   2.030000 15.625000   2.100000 ;
      RECT 13.295000   2.030000 15.625000   2.100000 ;
      RECT 13.295000   2.100000 15.695000   2.170000 ;
      RECT 13.295000   2.100000 15.695000   2.170000 ;
      RECT 13.295000   2.170000 15.765000   2.240000 ;
      RECT 13.295000   2.170000 15.765000   2.240000 ;
      RECT 13.295000   2.240000 15.835000   2.310000 ;
      RECT 13.295000   2.240000 15.835000   2.310000 ;
      RECT 13.295000   2.310000 15.905000   2.380000 ;
      RECT 13.295000   2.310000 15.905000   2.380000 ;
      RECT 13.295000   2.380000 15.975000   2.435000 ;
      RECT 13.295000   2.380000 15.975000   2.435000 ;
      RECT 13.295000   2.435000 16.030000   2.505000 ;
      RECT 13.295000   2.435000 16.030000   2.505000 ;
      RECT 13.295000   2.505000 16.100000   2.575000 ;
      RECT 13.295000   2.505000 16.100000   2.575000 ;
      RECT 13.295000   2.575000 16.170000   2.645000 ;
      RECT 13.295000   2.575000 16.170000   2.645000 ;
      RECT 13.295000   2.645000 16.240000   2.715000 ;
      RECT 13.295000   2.645000 16.240000   2.715000 ;
      RECT 13.295000   2.715000 16.310000   2.785000 ;
      RECT 13.295000   2.715000 16.310000   2.785000 ;
      RECT 13.295000   2.785000 16.380000   2.855000 ;
      RECT 13.295000   2.785000 16.380000   2.855000 ;
      RECT 13.295000   2.855000 16.450000   2.925000 ;
      RECT 13.295000   2.855000 16.450000   2.925000 ;
      RECT 13.295000   2.925000 16.520000   2.995000 ;
      RECT 13.295000   2.925000 16.520000   2.995000 ;
      RECT 13.295000   2.995000 16.590000   3.065000 ;
      RECT 13.295000   2.995000 16.590000   3.065000 ;
      RECT 13.295000   3.065000 16.660000   3.135000 ;
      RECT 13.295000   3.065000 16.660000   3.135000 ;
      RECT 13.295000   3.135000 16.730000   3.205000 ;
      RECT 13.295000   3.135000 16.730000   3.205000 ;
      RECT 13.295000   3.205000 16.800000   3.220000 ;
      RECT 13.295000   3.205000 16.800000   3.220000 ;
      RECT 13.295000   3.220000 16.815000   5.125000 ;
      RECT 13.305000  39.730000 13.855000  39.800000 ;
      RECT 13.320000  39.520000 13.480000  40.370000 ;
      RECT 13.320000  42.530000 29.845000  42.600000 ;
      RECT 13.320000  42.530000 29.845000  42.600000 ;
      RECT 13.365000   5.125000 16.815000   5.195000 ;
      RECT 13.365000   5.125000 16.815000   5.195000 ;
      RECT 13.375000  39.660000 13.925000  39.730000 ;
      RECT 13.390000  42.460000 29.845000  42.530000 ;
      RECT 13.390000  42.460000 29.845000  42.530000 ;
      RECT 13.435000   5.195000 16.815000   5.265000 ;
      RECT 13.435000   5.195000 16.815000   5.265000 ;
      RECT 13.445000  39.590000 13.995000  39.660000 ;
      RECT 13.460000  42.390000 29.845000  42.460000 ;
      RECT 13.460000  42.390000 29.845000  42.460000 ;
      RECT 13.505000   5.265000 16.815000   5.335000 ;
      RECT 13.505000   5.265000 16.815000   5.335000 ;
      RECT 13.515000  39.520000 14.065000  39.590000 ;
      RECT 13.530000  42.320000 29.845000  42.390000 ;
      RECT 13.530000  42.320000 29.845000  42.390000 ;
      RECT 13.575000   5.335000 16.815000   5.405000 ;
      RECT 13.575000   5.335000 16.815000   5.405000 ;
      RECT 13.585000  39.450000 14.135000  39.520000 ;
      RECT 13.600000  42.250000 29.845000  42.320000 ;
      RECT 13.600000  42.250000 29.845000  42.320000 ;
      RECT 13.645000   5.405000 16.815000   5.475000 ;
      RECT 13.645000   5.405000 16.815000   5.475000 ;
      RECT 13.655000  39.380000 14.205000  39.450000 ;
      RECT 13.670000  42.180000 29.845000  42.250000 ;
      RECT 13.670000  42.180000 29.845000  42.250000 ;
      RECT 13.690000  39.345000 15.195000  39.380000 ;
      RECT 13.715000   5.475000 16.815000   5.545000 ;
      RECT 13.715000   5.475000 16.815000   5.545000 ;
      RECT 13.740000  42.110000 29.845000  42.180000 ;
      RECT 13.740000  42.110000 29.845000  42.180000 ;
      RECT 13.760000  39.275000 15.230000  39.345000 ;
      RECT 13.785000   5.545000 16.815000   5.615000 ;
      RECT 13.785000   5.545000 16.815000   5.615000 ;
      RECT 13.810000  42.040000 29.845000  42.110000 ;
      RECT 13.810000  42.040000 29.845000  42.110000 ;
      RECT 13.830000  39.205000 15.300000  39.275000 ;
      RECT 13.855000   5.615000 16.815000   5.685000 ;
      RECT 13.855000   5.615000 16.815000   5.685000 ;
      RECT 13.880000  41.970000 29.845000  42.040000 ;
      RECT 13.880000  41.970000 29.845000  42.040000 ;
      RECT 13.900000  39.135000 15.370000  39.205000 ;
      RECT 13.910000  47.675000 29.985000  48.515000 ;
      RECT 13.925000   5.685000 16.815000   5.755000 ;
      RECT 13.925000   5.685000 16.815000   5.755000 ;
      RECT 13.950000  41.900000 29.845000  41.970000 ;
      RECT 13.950000  41.900000 29.845000  41.970000 ;
      RECT 13.970000  39.065000 15.440000  39.135000 ;
      RECT 13.995000   5.755000 16.815000   5.825000 ;
      RECT 13.995000   5.755000 16.815000   5.825000 ;
      RECT 14.020000  40.600000 29.985000  41.635000 ;
      RECT 14.020000  41.635000 29.985000  44.005000 ;
      RECT 14.020000  41.830000 29.845000  41.900000 ;
      RECT 14.020000  41.830000 29.845000  41.900000 ;
      RECT 14.035000  47.535000 29.845000  47.605000 ;
      RECT 14.035000  47.535000 29.845000  47.605000 ;
      RECT 14.040000  38.995000 15.510000  39.065000 ;
      RECT 14.065000   5.825000 16.815000   5.895000 ;
      RECT 14.065000   5.825000 16.815000   5.895000 ;
      RECT 14.090000  41.760000 29.845000  41.830000 ;
      RECT 14.090000  41.760000 29.845000  41.830000 ;
      RECT 14.105000  47.605000 29.845000  47.675000 ;
      RECT 14.105000  47.605000 29.845000  47.675000 ;
      RECT 14.110000  38.925000 15.580000  38.995000 ;
      RECT 14.135000   5.895000 16.815000   5.965000 ;
      RECT 14.135000   5.895000 16.815000   5.965000 ;
      RECT 14.160000  40.655000 29.845000  41.690000 ;
      RECT 14.160000  41.690000 29.845000  41.760000 ;
      RECT 14.160000  41.690000 29.845000  41.760000 ;
      RECT 14.175000  47.675000 29.845000  47.745000 ;
      RECT 14.175000  47.675000 29.845000  47.745000 ;
      RECT 14.180000  38.855000 15.650000  38.925000 ;
      RECT 14.195000  40.620000 29.845000  40.655000 ;
      RECT 14.195000  40.620000 29.845000  40.655000 ;
      RECT 14.205000   5.965000 16.815000   6.035000 ;
      RECT 14.205000   5.965000 16.815000   6.035000 ;
      RECT 14.245000  47.745000 29.845000  47.815000 ;
      RECT 14.245000  47.745000 29.845000  47.815000 ;
      RECT 14.250000  38.785000 15.720000  38.855000 ;
      RECT 14.265000  40.550000 29.845000  40.620000 ;
      RECT 14.265000  40.550000 29.845000  40.620000 ;
      RECT 14.275000   6.035000 16.815000   6.105000 ;
      RECT 14.275000   6.035000 16.815000   6.105000 ;
      RECT 14.315000  47.815000 29.845000  47.885000 ;
      RECT 14.315000  47.815000 29.845000  47.885000 ;
      RECT 14.320000  38.715000 15.790000  38.785000 ;
      RECT 14.335000  40.480000 29.845000  40.550000 ;
      RECT 14.335000  40.480000 29.845000  40.550000 ;
      RECT 14.345000   6.105000 16.815000   6.175000 ;
      RECT 14.345000   6.105000 16.815000   6.175000 ;
      RECT 14.370000   6.395000 16.955000   6.615000 ;
      RECT 14.370000   6.615000 16.470000   7.100000 ;
      RECT 14.370000   7.100000 16.470000  11.600000 ;
      RECT 14.370000  11.600000 16.565000  11.695000 ;
      RECT 14.370000  11.695000 16.565000  12.320000 ;
      RECT 14.370000  12.320000 16.470000  12.415000 ;
      RECT 14.370000  12.415000 16.470000  18.055000 ;
      RECT 14.370000  18.055000 16.470000  19.470000 ;
      RECT 14.385000  47.885000 29.845000  47.955000 ;
      RECT 14.385000  47.885000 29.845000  47.955000 ;
      RECT 14.390000  38.645000 15.860000  38.715000 ;
      RECT 14.405000  40.410000 29.845000  40.480000 ;
      RECT 14.405000  40.410000 29.845000  40.480000 ;
      RECT 14.415000   6.175000 16.815000   6.245000 ;
      RECT 14.415000   6.175000 16.815000   6.245000 ;
      RECT 14.455000  47.955000 29.845000  48.025000 ;
      RECT 14.455000  47.955000 29.845000  48.025000 ;
      RECT 14.460000  38.575000 15.930000  38.645000 ;
      RECT 14.475000  40.340000 29.845000  40.410000 ;
      RECT 14.475000  40.340000 29.845000  40.410000 ;
      RECT 14.485000   6.245000 16.815000   6.315000 ;
      RECT 14.485000   6.245000 16.815000   6.315000 ;
      RECT 14.510000   6.315000 16.815000   6.340000 ;
      RECT 14.510000   6.315000 16.815000   6.340000 ;
      RECT 14.510000   6.560000 16.745000   6.630000 ;
      RECT 14.510000   6.630000 16.675000   6.700000 ;
      RECT 14.510000   6.700000 16.605000   6.770000 ;
      RECT 14.510000   6.770000 16.535000   6.840000 ;
      RECT 14.510000   6.840000 16.465000   6.910000 ;
      RECT 14.510000   6.910000 16.395000   6.980000 ;
      RECT 14.510000   6.980000 16.330000   7.045000 ;
      RECT 14.510000   7.045000 16.330000  11.655000 ;
      RECT 14.510000  11.655000 16.330000  11.705000 ;
      RECT 14.510000  11.705000 16.380000  11.750000 ;
      RECT 14.510000  11.750000 16.425000  12.265000 ;
      RECT 14.510000  12.265000 16.380000  12.310000 ;
      RECT 14.510000  12.310000 16.335000  12.355000 ;
      RECT 14.510000  12.355000 16.330000  12.360000 ;
      RECT 14.510000  12.360000 16.330000  18.000000 ;
      RECT 14.525000  48.025000 29.845000  48.095000 ;
      RECT 14.525000  48.025000 29.845000  48.095000 ;
      RECT 14.530000  38.505000 16.000000  38.575000 ;
      RECT 14.545000  40.270000 29.845000  40.340000 ;
      RECT 14.545000  40.270000 29.845000  40.340000 ;
      RECT 14.560000  40.060000 29.985000  40.600000 ;
      RECT 14.580000   6.340000 16.815000   6.410000 ;
      RECT 14.580000   6.340000 16.815000   6.410000 ;
      RECT 14.580000  18.000000 16.330000  18.070000 ;
      RECT 14.595000  48.095000 29.845000  48.165000 ;
      RECT 14.595000  48.095000 29.845000  48.165000 ;
      RECT 14.600000  38.435000 16.070000  38.505000 ;
      RECT 14.615000  40.200000 29.845000  40.270000 ;
      RECT 14.615000  40.200000 29.845000  40.270000 ;
      RECT 14.650000   6.410000 16.815000   6.480000 ;
      RECT 14.650000   6.410000 16.815000   6.480000 ;
      RECT 14.650000  18.070000 16.330000  18.140000 ;
      RECT 14.665000  48.165000 29.845000  48.235000 ;
      RECT 14.665000  48.165000 29.845000  48.235000 ;
      RECT 14.670000  38.365000 16.140000  38.435000 ;
      RECT 14.720000   6.480000 16.815000   6.550000 ;
      RECT 14.720000   6.480000 16.815000   6.550000 ;
      RECT 14.720000  18.140000 16.330000  18.210000 ;
      RECT 14.730000   6.550000 16.815000   6.560000 ;
      RECT 14.730000   6.550000 16.815000   6.560000 ;
      RECT 14.735000  48.235000 29.845000  48.305000 ;
      RECT 14.735000  48.235000 29.845000  48.305000 ;
      RECT 14.740000  38.295000 16.210000  38.365000 ;
      RECT 14.750000  48.515000 29.985000  51.370000 ;
      RECT 14.750000  51.370000 29.565000  51.790000 ;
      RECT 14.750000  51.790000 24.535000  53.195000 ;
      RECT 14.750000  53.195000 24.535000  56.895000 ;
      RECT 14.750000  56.895000 24.210000  57.220000 ;
      RECT 14.750000  57.220000 22.940000  57.765000 ;
      RECT 14.750000  57.765000 22.940000  57.780000 ;
      RECT 14.765000  57.780000 76.775000  57.990000 ;
      RECT 14.790000  18.210000 16.330000  18.280000 ;
      RECT 14.800000   6.560000 16.745000   6.630000 ;
      RECT 14.800000   6.560000 16.745000   6.630000 ;
      RECT 14.805000  48.305000 29.845000  48.375000 ;
      RECT 14.805000  48.305000 29.845000  48.375000 ;
      RECT 14.810000  38.225000 16.280000  38.295000 ;
      RECT 14.860000  18.280000 16.330000  18.350000 ;
      RECT 14.870000   6.630000 16.675000   6.700000 ;
      RECT 14.870000   6.630000 16.675000   6.700000 ;
      RECT 14.875000  48.375000 29.845000  48.445000 ;
      RECT 14.875000  48.375000 29.845000  48.445000 ;
      RECT 14.880000  38.155000 16.350000  38.225000 ;
      RECT 14.890000  48.445000 29.845000  48.460000 ;
      RECT 14.890000  48.445000 29.845000  48.460000 ;
      RECT 14.890000  48.460000 29.845000  51.315000 ;
      RECT 14.890000  51.315000 29.775000  51.385000 ;
      RECT 14.890000  51.315000 29.775000  51.385000 ;
      RECT 14.890000  51.385000 29.705000  51.455000 ;
      RECT 14.890000  51.385000 29.705000  51.455000 ;
      RECT 14.890000  51.455000 29.635000  51.525000 ;
      RECT 14.890000  51.455000 29.635000  51.525000 ;
      RECT 14.890000  51.525000 29.565000  51.595000 ;
      RECT 14.890000  51.525000 29.565000  51.595000 ;
      RECT 14.890000  51.595000 29.510000  51.650000 ;
      RECT 14.890000  51.595000 29.510000  51.650000 ;
      RECT 14.890000  51.650000 24.395000  56.840000 ;
      RECT 14.890000  51.650000 25.815000  51.720000 ;
      RECT 14.890000  51.650000 25.815000  51.720000 ;
      RECT 14.890000  51.720000 25.745000  51.790000 ;
      RECT 14.890000  51.720000 25.745000  51.790000 ;
      RECT 14.890000  51.790000 25.675000  51.860000 ;
      RECT 14.890000  51.790000 25.675000  51.860000 ;
      RECT 14.890000  51.860000 25.605000  51.930000 ;
      RECT 14.890000  51.860000 25.605000  51.930000 ;
      RECT 14.890000  51.930000 25.535000  52.000000 ;
      RECT 14.890000  51.930000 25.535000  52.000000 ;
      RECT 14.890000  52.000000 25.465000  52.070000 ;
      RECT 14.890000  52.000000 25.465000  52.070000 ;
      RECT 14.890000  52.070000 25.395000  52.140000 ;
      RECT 14.890000  52.070000 25.395000  52.140000 ;
      RECT 14.890000  52.140000 25.325000  52.210000 ;
      RECT 14.890000  52.140000 25.325000  52.210000 ;
      RECT 14.890000  52.210000 25.255000  52.280000 ;
      RECT 14.890000  52.210000 25.255000  52.280000 ;
      RECT 14.890000  52.280000 25.185000  52.350000 ;
      RECT 14.890000  52.280000 25.185000  52.350000 ;
      RECT 14.890000  52.350000 25.115000  52.420000 ;
      RECT 14.890000  52.350000 25.115000  52.420000 ;
      RECT 14.890000  52.420000 25.045000  52.490000 ;
      RECT 14.890000  52.420000 25.045000  52.490000 ;
      RECT 14.890000  52.490000 24.975000  52.560000 ;
      RECT 14.890000  52.490000 24.975000  52.560000 ;
      RECT 14.890000  52.560000 24.905000  52.630000 ;
      RECT 14.890000  52.560000 24.905000  52.630000 ;
      RECT 14.890000  52.630000 24.835000  52.700000 ;
      RECT 14.890000  52.630000 24.835000  52.700000 ;
      RECT 14.890000  52.700000 24.765000  52.770000 ;
      RECT 14.890000  52.700000 24.765000  52.770000 ;
      RECT 14.890000  52.770000 24.695000  52.840000 ;
      RECT 14.890000  52.770000 24.695000  52.840000 ;
      RECT 14.890000  52.840000 24.625000  52.910000 ;
      RECT 14.890000  52.840000 24.625000  52.910000 ;
      RECT 14.890000  52.910000 24.555000  52.980000 ;
      RECT 14.890000  52.910000 24.555000  52.980000 ;
      RECT 14.890000  52.980000 24.485000  53.050000 ;
      RECT 14.890000  52.980000 24.485000  53.050000 ;
      RECT 14.890000  53.050000 24.415000  53.120000 ;
      RECT 14.890000  53.050000 24.415000  53.120000 ;
      RECT 14.890000  53.120000 24.395000  53.140000 ;
      RECT 14.890000  53.120000 24.395000  53.140000 ;
      RECT 14.890000  53.140000 24.395000  56.840000 ;
      RECT 14.890000  56.840000 24.325000  56.910000 ;
      RECT 14.890000  56.840000 24.325000  56.910000 ;
      RECT 14.890000  56.910000 24.255000  56.980000 ;
      RECT 14.890000  56.910000 24.255000  56.980000 ;
      RECT 14.890000  56.980000 24.185000  57.050000 ;
      RECT 14.890000  56.980000 24.185000  57.050000 ;
      RECT 14.890000  57.050000 24.155000  57.080000 ;
      RECT 14.890000  57.050000 24.155000  57.080000 ;
      RECT 14.890000  57.080000 22.800000  57.710000 ;
      RECT 14.930000  18.350000 16.330000  18.420000 ;
      RECT 14.940000   6.700000 16.605000   6.770000 ;
      RECT 14.940000   6.700000 16.605000   6.770000 ;
      RECT 14.950000  38.085000 16.420000  38.155000 ;
      RECT 14.960000  57.710000 22.800000  57.780000 ;
      RECT 14.960000  57.710000 22.800000  57.780000 ;
      RECT 14.975000  57.990000 76.775000  58.450000 ;
      RECT 15.000000  18.420000 16.330000  18.490000 ;
      RECT 15.010000   6.770000 16.535000   6.840000 ;
      RECT 15.010000   6.770000 16.535000   6.840000 ;
      RECT 15.020000  38.015000 16.490000  38.085000 ;
      RECT 15.030000  57.780000 22.800000  57.850000 ;
      RECT 15.030000  57.780000 22.800000  57.850000 ;
      RECT 15.070000  18.490000 16.330000  18.560000 ;
      RECT 15.080000   6.840000 16.465000   6.910000 ;
      RECT 15.080000   6.840000 16.465000   6.910000 ;
      RECT 15.090000  37.945000 16.560000  38.015000 ;
      RECT 15.100000  57.850000 22.800000  57.920000 ;
      RECT 15.100000  57.850000 22.800000  57.920000 ;
      RECT 15.105000  57.920000 76.635000  57.925000 ;
      RECT 15.105000  57.920000 76.635000  57.925000 ;
      RECT 15.110000  57.925000 76.635000  57.930000 ;
      RECT 15.110000  57.925000 76.635000  57.930000 ;
      RECT 15.115000  57.920000 76.635000  73.500000 ;
      RECT 15.115000  57.920000 76.635000  73.500000 ;
      RECT 15.115000  57.920000 76.635000  73.500000 ;
      RECT 15.115000  57.920000 76.635000  73.500000 ;
      RECT 15.115000  57.930000 76.635000  57.935000 ;
      RECT 15.115000  57.930000 76.635000  57.935000 ;
      RECT 15.115000  57.935000 76.635000  58.590000 ;
      RECT 15.140000  18.560000 16.330000  18.630000 ;
      RECT 15.150000   6.910000 16.395000   6.980000 ;
      RECT 15.150000   6.910000 16.395000   6.980000 ;
      RECT 15.160000  37.875000 16.630000  37.945000 ;
      RECT 15.210000  18.630000 16.330000  18.700000 ;
      RECT 15.215000   6.980000 16.330000   7.045000 ;
      RECT 15.215000   6.980000 16.330000   7.045000 ;
      RECT 15.230000  37.805000 16.700000  37.875000 ;
      RECT 15.280000  18.700000 16.330000  18.770000 ;
      RECT 15.300000  37.735000 16.770000  37.805000 ;
      RECT 15.350000  18.770000 16.330000  18.840000 ;
      RECT 15.370000  32.130000 16.225000  34.380000 ;
      RECT 15.370000  34.380000 17.435000  35.590000 ;
      RECT 15.370000  35.590000 17.435000  37.335000 ;
      RECT 15.370000  37.335000 17.305000  37.470000 ;
      RECT 15.370000  37.665000 16.840000  37.735000 ;
      RECT 15.420000  18.840000 16.330000  18.910000 ;
      RECT 15.440000  37.595000 16.910000  37.665000 ;
      RECT 15.490000  18.910000 16.330000  18.980000 ;
      RECT 15.510000  32.185000 16.085000  34.435000 ;
      RECT 15.510000  34.435000 16.085000  34.505000 ;
      RECT 15.510000  34.505000 16.155000  34.575000 ;
      RECT 15.510000  34.575000 16.225000  34.645000 ;
      RECT 15.510000  34.645000 16.295000  34.715000 ;
      RECT 15.510000  34.715000 16.365000  34.785000 ;
      RECT 15.510000  34.785000 16.435000  34.855000 ;
      RECT 15.510000  34.855000 16.505000  34.925000 ;
      RECT 15.510000  34.925000 16.575000  34.995000 ;
      RECT 15.510000  34.995000 16.645000  35.065000 ;
      RECT 15.510000  35.065000 16.715000  35.135000 ;
      RECT 15.510000  35.135000 16.785000  35.205000 ;
      RECT 15.510000  35.205000 16.855000  35.275000 ;
      RECT 15.510000  35.275000 16.925000  35.345000 ;
      RECT 15.510000  35.345000 16.995000  35.415000 ;
      RECT 15.510000  35.415000 17.065000  35.485000 ;
      RECT 15.510000  35.485000 17.135000  35.555000 ;
      RECT 15.510000  35.555000 17.205000  35.625000 ;
      RECT 15.510000  35.625000 17.275000  35.645000 ;
      RECT 15.510000  35.645000 17.295000  37.280000 ;
      RECT 15.510000  37.280000 17.225000  37.350000 ;
      RECT 15.510000  37.350000 17.155000  37.420000 ;
      RECT 15.510000  37.420000 17.085000  37.490000 ;
      RECT 15.510000  37.490000 17.050000  37.525000 ;
      RECT 15.510000  37.525000 16.980000  37.595000 ;
      RECT 15.560000  18.980000 16.330000  19.050000 ;
      RECT 15.575000  32.120000 16.085000  32.185000 ;
      RECT 15.590000  40.145000 29.845000  40.200000 ;
      RECT 15.590000  40.145000 29.845000  40.200000 ;
      RECT 15.630000  19.050000 16.330000  19.120000 ;
      RECT 15.645000  32.050000 16.085000  32.120000 ;
      RECT 15.660000  40.075000 29.845000  40.145000 ;
      RECT 15.660000  40.075000 29.845000  40.145000 ;
      RECT 15.700000  19.120000 16.330000  19.190000 ;
      RECT 15.715000  31.980000 16.085000  32.050000 ;
      RECT 15.730000  40.005000 29.845000  40.075000 ;
      RECT 15.730000  40.005000 29.845000  40.075000 ;
      RECT 15.770000  19.190000 16.330000  19.260000 ;
      RECT 15.785000  19.470000 16.470000  31.255000 ;
      RECT 15.785000  31.255000 16.225000  31.500000 ;
      RECT 15.785000  31.500000 16.225000  31.715000 ;
      RECT 15.785000  31.715000 16.225000  32.130000 ;
      RECT 15.785000  31.910000 16.085000  31.980000 ;
      RECT 15.800000  39.935000 29.845000  40.005000 ;
      RECT 15.800000  39.935000 29.845000  40.005000 ;
      RECT 15.840000  19.260000 16.330000  19.330000 ;
      RECT 15.855000  31.840000 16.085000  31.910000 ;
      RECT 15.870000  39.865000 29.845000  39.935000 ;
      RECT 15.870000  39.865000 29.845000  39.935000 ;
      RECT 15.910000  19.330000 16.330000  19.400000 ;
      RECT 15.925000  19.400000 16.330000  19.415000 ;
      RECT 15.925000  19.415000 16.330000  31.200000 ;
      RECT 15.925000  31.200000 16.260000  31.270000 ;
      RECT 15.925000  31.270000 16.190000  31.340000 ;
      RECT 15.925000  31.340000 16.120000  31.410000 ;
      RECT 15.925000  31.410000 16.085000  31.445000 ;
      RECT 15.925000  31.445000 16.085000  31.770000 ;
      RECT 15.925000  31.770000 16.085000  31.840000 ;
      RECT 15.940000  39.795000 29.845000  39.865000 ;
      RECT 15.940000  39.795000 29.845000  39.865000 ;
      RECT 16.010000  39.725000 29.845000  39.795000 ;
      RECT 16.010000  39.725000 29.845000  39.795000 ;
      RECT 16.080000  39.655000 29.845000  39.725000 ;
      RECT 16.080000  39.655000 29.845000  39.725000 ;
      RECT 16.150000  39.585000 29.845000  39.655000 ;
      RECT 16.150000  39.585000 29.845000  39.655000 ;
      RECT 16.220000  39.515000 29.845000  39.585000 ;
      RECT 16.220000  39.515000 29.845000  39.585000 ;
      RECT 16.290000  39.445000 29.845000  39.515000 ;
      RECT 16.290000  39.445000 29.845000  39.515000 ;
      RECT 16.360000  39.375000 29.845000  39.445000 ;
      RECT 16.360000  39.375000 29.845000  39.445000 ;
      RECT 16.430000  39.305000 29.845000  39.375000 ;
      RECT 16.430000  39.305000 29.845000  39.375000 ;
      RECT 16.445000  39.095000 29.985000  40.060000 ;
      RECT 16.500000  39.235000 29.845000  39.305000 ;
      RECT 16.500000  39.235000 29.845000  39.305000 ;
      RECT 16.550000  39.185000 22.815000  39.235000 ;
      RECT 16.550000  39.185000 22.815000  39.235000 ;
      RECT 16.620000  39.115000 22.815000  39.185000 ;
      RECT 16.620000  39.115000 22.815000  39.185000 ;
      RECT 16.690000  39.045000 22.815000  39.115000 ;
      RECT 16.690000  39.045000 22.815000  39.115000 ;
      RECT 16.710000   0.000000 22.215000   2.150000 ;
      RECT 16.710000   2.150000 22.215000   2.935000 ;
      RECT 16.760000  38.975000 22.815000  39.045000 ;
      RECT 16.760000  38.975000 22.815000  39.045000 ;
      RECT 16.765000  31.730000 23.335000  34.150000 ;
      RECT 16.765000  34.150000 23.335000  35.360000 ;
      RECT 16.830000  38.905000 22.815000  38.975000 ;
      RECT 16.830000  38.905000 22.815000  38.975000 ;
      RECT 16.850000   0.000000 22.075000   2.095000 ;
      RECT 16.900000  38.835000 22.815000  38.905000 ;
      RECT 16.900000  38.835000 22.815000  38.905000 ;
      RECT 16.905000  31.785000 23.195000  34.095000 ;
      RECT 16.920000   2.095000 22.075000   2.165000 ;
      RECT 16.920000   2.095000 22.075000   2.165000 ;
      RECT 16.940000  31.750000 23.195000  31.785000 ;
      RECT 16.940000  31.750000 23.195000  31.785000 ;
      RECT 16.970000  38.765000 22.815000  38.835000 ;
      RECT 16.970000  38.765000 22.815000  38.835000 ;
      RECT 16.975000  34.095000 23.195000  34.165000 ;
      RECT 16.975000  34.095000 23.195000  34.165000 ;
      RECT 16.985000  38.555000 22.955000  39.095000 ;
      RECT 16.990000   2.165000 22.075000   2.235000 ;
      RECT 16.990000   2.165000 22.075000   2.235000 ;
      RECT 17.010000   7.330000 22.625000  14.545000 ;
      RECT 17.010000  14.545000 23.515000  15.435000 ;
      RECT 17.010000  15.435000 23.515000  24.940000 ;
      RECT 17.010000  24.940000 23.335000  25.120000 ;
      RECT 17.010000  25.120000 23.335000  31.485000 ;
      RECT 17.010000  31.485000 23.335000  31.730000 ;
      RECT 17.010000  31.680000 23.195000  31.750000 ;
      RECT 17.010000  31.680000 23.195000  31.750000 ;
      RECT 17.040000  38.695000 22.815000  38.765000 ;
      RECT 17.040000  38.695000 22.815000  38.765000 ;
      RECT 17.045000  34.165000 23.195000  34.235000 ;
      RECT 17.045000  34.165000 23.195000  34.235000 ;
      RECT 17.060000   2.235000 22.075000   2.305000 ;
      RECT 17.060000   2.235000 22.075000   2.305000 ;
      RECT 17.080000  31.610000 23.195000  31.680000 ;
      RECT 17.080000  31.610000 23.195000  31.680000 ;
      RECT 17.110000  38.625000 22.815000  38.695000 ;
      RECT 17.110000  38.625000 22.815000  38.695000 ;
      RECT 17.115000  34.235000 23.195000  34.305000 ;
      RECT 17.115000  34.235000 23.195000  34.305000 ;
      RECT 17.130000   2.305000 22.075000   2.375000 ;
      RECT 17.130000   2.305000 22.075000   2.375000 ;
      RECT 17.150000   7.385000 22.485000  14.600000 ;
      RECT 17.150000   7.385000 22.485000  15.490000 ;
      RECT 17.150000  14.600000 22.485000  14.670000 ;
      RECT 17.150000  14.600000 22.485000  14.670000 ;
      RECT 17.150000  14.670000 22.555000  14.740000 ;
      RECT 17.150000  14.670000 22.555000  14.740000 ;
      RECT 17.150000  14.740000 22.625000  14.810000 ;
      RECT 17.150000  14.740000 22.625000  14.810000 ;
      RECT 17.150000  14.810000 22.695000  14.880000 ;
      RECT 17.150000  14.810000 22.695000  14.880000 ;
      RECT 17.150000  14.880000 22.765000  14.950000 ;
      RECT 17.150000  14.880000 22.765000  14.950000 ;
      RECT 17.150000  14.950000 22.835000  15.020000 ;
      RECT 17.150000  14.950000 22.835000  15.020000 ;
      RECT 17.150000  15.020000 22.905000  15.090000 ;
      RECT 17.150000  15.020000 22.905000  15.090000 ;
      RECT 17.150000  15.090000 22.975000  15.160000 ;
      RECT 17.150000  15.090000 22.975000  15.160000 ;
      RECT 17.150000  15.160000 23.045000  15.230000 ;
      RECT 17.150000  15.160000 23.045000  15.230000 ;
      RECT 17.150000  15.230000 23.115000  15.300000 ;
      RECT 17.150000  15.230000 23.115000  15.300000 ;
      RECT 17.150000  15.300000 23.185000  15.370000 ;
      RECT 17.150000  15.300000 23.185000  15.370000 ;
      RECT 17.150000  15.370000 23.255000  15.440000 ;
      RECT 17.150000  15.370000 23.255000  15.440000 ;
      RECT 17.150000  15.440000 23.325000  15.490000 ;
      RECT 17.150000  15.440000 23.325000  15.490000 ;
      RECT 17.150000  15.490000 23.375000  24.885000 ;
      RECT 17.150000  24.885000 23.305000  24.955000 ;
      RECT 17.150000  24.885000 23.305000  24.955000 ;
      RECT 17.150000  24.955000 23.235000  25.025000 ;
      RECT 17.150000  24.955000 23.235000  25.025000 ;
      RECT 17.150000  25.025000 23.195000  25.065000 ;
      RECT 17.150000  25.025000 23.195000  25.065000 ;
      RECT 17.150000  25.065000 23.195000  31.540000 ;
      RECT 17.150000  31.540000 23.195000  31.610000 ;
      RECT 17.150000  31.540000 23.195000  31.610000 ;
      RECT 17.165000   7.370000 22.485000   7.385000 ;
      RECT 17.165000   7.370000 22.485000   7.385000 ;
      RECT 17.180000  38.355000 23.135000  38.555000 ;
      RECT 17.180000  38.555000 22.815000  38.625000 ;
      RECT 17.180000  38.555000 22.815000  38.625000 ;
      RECT 17.185000  34.305000 23.195000  34.375000 ;
      RECT 17.185000  34.305000 23.195000  34.375000 ;
      RECT 17.200000   2.375000 22.075000   2.445000 ;
      RECT 17.200000   2.375000 22.075000   2.445000 ;
      RECT 17.235000   7.300000 22.485000   7.370000 ;
      RECT 17.235000   7.300000 22.485000   7.370000 ;
      RECT 17.250000  38.485000 22.815000  38.555000 ;
      RECT 17.250000  38.485000 22.815000  38.555000 ;
      RECT 17.255000  34.375000 23.195000  34.445000 ;
      RECT 17.255000  34.375000 23.195000  34.445000 ;
      RECT 17.270000   2.445000 22.075000   2.515000 ;
      RECT 17.270000   2.445000 22.075000   2.515000 ;
      RECT 17.305000   7.230000 22.485000   7.300000 ;
      RECT 17.305000   7.230000 22.485000   7.300000 ;
      RECT 17.320000  38.415000 22.815000  38.485000 ;
      RECT 17.320000  38.415000 22.815000  38.485000 ;
      RECT 17.325000  34.445000 23.195000  34.515000 ;
      RECT 17.325000  34.445000 23.195000  34.515000 ;
      RECT 17.340000   2.515000 22.075000   2.585000 ;
      RECT 17.340000   2.515000 22.075000   2.585000 ;
      RECT 17.375000   7.160000 22.485000   7.230000 ;
      RECT 17.375000   7.160000 22.485000   7.230000 ;
      RECT 17.380000  38.355000 23.080000  38.415000 ;
      RECT 17.380000  38.355000 23.080000  38.415000 ;
      RECT 17.395000  34.515000 23.195000  34.585000 ;
      RECT 17.395000  34.515000 23.195000  34.585000 ;
      RECT 17.410000   2.585000 22.075000   2.655000 ;
      RECT 17.410000   2.585000 22.075000   2.655000 ;
      RECT 17.435000  38.300000 23.140000  38.355000 ;
      RECT 17.435000  38.300000 23.140000  38.355000 ;
      RECT 17.445000   6.895000 22.625000   7.330000 ;
      RECT 17.445000   7.090000 22.485000   7.160000 ;
      RECT 17.445000   7.090000 22.485000   7.160000 ;
      RECT 17.465000  34.585000 23.195000  34.655000 ;
      RECT 17.465000  34.585000 23.195000  34.655000 ;
      RECT 17.480000   2.655000 22.075000   2.725000 ;
      RECT 17.480000   2.655000 22.075000   2.725000 ;
      RECT 17.485000  38.250000 23.195000  38.300000 ;
      RECT 17.485000  38.250000 23.195000  38.300000 ;
      RECT 17.495000   2.935000 22.215000   6.480000 ;
      RECT 17.495000   6.480000 22.575000   6.845000 ;
      RECT 17.495000   6.845000 22.625000   6.895000 ;
      RECT 17.515000   7.020000 22.485000   7.090000 ;
      RECT 17.515000   7.020000 22.485000   7.090000 ;
      RECT 17.535000  34.655000 23.195000  34.725000 ;
      RECT 17.535000  34.655000 23.195000  34.725000 ;
      RECT 17.550000   2.725000 22.075000   2.795000 ;
      RECT 17.550000   2.725000 22.075000   2.795000 ;
      RECT 17.555000  38.180000 23.195000  38.250000 ;
      RECT 17.555000  38.180000 23.195000  38.250000 ;
      RECT 17.585000   6.950000 22.485000   7.020000 ;
      RECT 17.585000   6.950000 22.485000   7.020000 ;
      RECT 17.605000  34.725000 23.195000  34.795000 ;
      RECT 17.605000  34.725000 23.195000  34.795000 ;
      RECT 17.610000   6.925000 22.460000   6.950000 ;
      RECT 17.610000   6.925000 22.460000   6.950000 ;
      RECT 17.620000   2.795000 22.075000   2.865000 ;
      RECT 17.620000   2.795000 22.075000   2.865000 ;
      RECT 17.625000  38.110000 23.195000  38.180000 ;
      RECT 17.625000  38.110000 23.195000  38.180000 ;
      RECT 17.635000   0.000000 22.075000   6.540000 ;
      RECT 17.635000   0.000000 22.075000   6.540000 ;
      RECT 17.635000   2.865000 22.075000   2.880000 ;
      RECT 17.635000   2.865000 22.075000   2.880000 ;
      RECT 17.635000   2.880000 22.075000   6.540000 ;
      RECT 17.635000   2.880000 22.075000   6.900000 ;
      RECT 17.635000   2.880000 22.075000   6.900000 ;
      RECT 17.635000   2.880000 22.075000   6.900000 ;
      RECT 17.635000   2.880000 22.075000   6.900000 ;
      RECT 17.635000   6.540000 22.075000   6.610000 ;
      RECT 17.635000   6.540000 22.075000   6.610000 ;
      RECT 17.635000   6.610000 22.145000   6.680000 ;
      RECT 17.635000   6.610000 22.145000   6.680000 ;
      RECT 17.635000   6.680000 22.215000   6.750000 ;
      RECT 17.635000   6.680000 22.215000   6.750000 ;
      RECT 17.635000   6.750000 22.285000   6.820000 ;
      RECT 17.635000   6.750000 22.285000   6.820000 ;
      RECT 17.635000   6.820000 22.355000   6.890000 ;
      RECT 17.635000   6.820000 22.355000   6.890000 ;
      RECT 17.635000   6.890000 22.425000   6.900000 ;
      RECT 17.635000   6.890000 22.425000   6.900000 ;
      RECT 17.635000   6.900000 22.435000   6.925000 ;
      RECT 17.635000   6.900000 22.435000   6.925000 ;
      RECT 17.675000  34.795000 23.195000  34.865000 ;
      RECT 17.675000  34.795000 23.195000  34.865000 ;
      RECT 17.695000  38.040000 23.195000  38.110000 ;
      RECT 17.695000  38.040000 23.195000  38.110000 ;
      RECT 17.745000  34.865000 23.195000  34.935000 ;
      RECT 17.745000  34.865000 23.195000  34.935000 ;
      RECT 17.765000  37.970000 23.195000  38.040000 ;
      RECT 17.765000  37.970000 23.195000  38.040000 ;
      RECT 17.815000  34.935000 23.195000  35.005000 ;
      RECT 17.815000  34.935000 23.195000  35.005000 ;
      RECT 17.835000  37.900000 23.195000  37.970000 ;
      RECT 17.835000  37.900000 23.195000  37.970000 ;
      RECT 17.885000  35.005000 23.195000  35.075000 ;
      RECT 17.885000  35.005000 23.195000  35.075000 ;
      RECT 17.905000  37.830000 23.195000  37.900000 ;
      RECT 17.905000  37.830000 23.195000  37.900000 ;
      RECT 17.955000  35.075000 23.195000  35.145000 ;
      RECT 17.955000  35.075000 23.195000  35.145000 ;
      RECT 17.975000  35.360000 23.335000  37.565000 ;
      RECT 17.975000  37.565000 23.335000  38.355000 ;
      RECT 17.975000  37.760000 23.195000  37.830000 ;
      RECT 17.975000  37.760000 23.195000  37.830000 ;
      RECT 18.025000  35.145000 23.195000  35.215000 ;
      RECT 18.025000  35.145000 23.195000  35.215000 ;
      RECT 18.045000  37.690000 23.195000  37.760000 ;
      RECT 18.045000  37.690000 23.195000  37.760000 ;
      RECT 18.095000  35.215000 23.195000  35.285000 ;
      RECT 18.095000  35.215000 23.195000  35.285000 ;
      RECT 18.115000  31.540000 23.195000  37.620000 ;
      RECT 18.115000  35.285000 23.195000  35.305000 ;
      RECT 18.115000  35.285000 23.195000  35.305000 ;
      RECT 18.115000  35.305000 23.195000  37.620000 ;
      RECT 18.115000  37.620000 23.195000  37.690000 ;
      RECT 18.115000  37.620000 23.195000  37.690000 ;
      RECT 22.755000   0.000000 26.460000   1.835000 ;
      RECT 22.755000   1.835000 28.350000   4.130000 ;
      RECT 22.755000   4.130000 29.070000   4.850000 ;
      RECT 22.755000   4.850000 29.070000   6.255000 ;
      RECT 22.755000   6.255000 29.070000   6.665000 ;
      RECT 22.895000   0.000000 26.320000   1.975000 ;
      RECT 22.895000   0.000000 26.320000   4.185000 ;
      RECT 22.895000   0.000000 26.320000   6.200000 ;
      RECT 22.895000   0.000000 26.320000   6.200000 ;
      RECT 22.895000   0.000000 26.320000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   4.185000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   4.185000 28.210000   4.255000 ;
      RECT 22.895000   4.185000 28.210000   4.255000 ;
      RECT 22.895000   4.255000 28.280000   4.325000 ;
      RECT 22.895000   4.255000 28.280000   4.325000 ;
      RECT 22.895000   4.325000 28.350000   4.395000 ;
      RECT 22.895000   4.325000 28.350000   4.395000 ;
      RECT 22.895000   4.395000 28.420000   4.465000 ;
      RECT 22.895000   4.395000 28.420000   4.465000 ;
      RECT 22.895000   4.465000 28.490000   4.535000 ;
      RECT 22.895000   4.465000 28.490000   4.535000 ;
      RECT 22.895000   4.535000 28.560000   4.605000 ;
      RECT 22.895000   4.535000 28.560000   4.605000 ;
      RECT 22.895000   4.605000 28.630000   4.675000 ;
      RECT 22.895000   4.605000 28.630000   4.675000 ;
      RECT 22.895000   4.675000 28.700000   4.745000 ;
      RECT 22.895000   4.675000 28.700000   4.745000 ;
      RECT 22.895000   4.745000 28.770000   4.815000 ;
      RECT 22.895000   4.745000 28.770000   4.815000 ;
      RECT 22.895000   4.815000 28.840000   4.885000 ;
      RECT 22.895000   4.815000 28.840000   4.885000 ;
      RECT 22.895000   4.885000 28.910000   4.905000 ;
      RECT 22.895000   4.885000 28.910000   4.905000 ;
      RECT 22.895000   4.905000 28.930000   6.200000 ;
      RECT 22.965000   6.200000 28.930000   6.270000 ;
      RECT 22.965000   6.200000 28.930000   6.270000 ;
      RECT 23.035000   6.270000 28.930000   6.340000 ;
      RECT 23.035000   6.270000 28.930000   6.340000 ;
      RECT 23.105000   6.340000 28.930000   6.410000 ;
      RECT 23.105000   6.340000 28.930000   6.410000 ;
      RECT 23.165000   6.665000 29.070000   6.920000 ;
      RECT 23.165000   6.920000 31.550000  14.315000 ;
      RECT 23.165000  14.315000 31.550000  15.205000 ;
      RECT 23.175000   6.410000 28.930000   6.480000 ;
      RECT 23.175000   6.410000 28.930000   6.480000 ;
      RECT 23.245000   6.480000 28.930000   6.550000 ;
      RECT 23.245000   6.480000 28.930000   6.550000 ;
      RECT 23.305000   6.550000 28.930000   6.610000 ;
      RECT 23.305000   6.550000 28.930000   6.610000 ;
      RECT 23.305000   6.610000 28.930000   7.060000 ;
      RECT 23.305000   7.060000 31.410000  14.260000 ;
      RECT 23.375000  14.260000 31.410000  14.330000 ;
      RECT 23.375000  14.260000 31.410000  14.330000 ;
      RECT 23.445000  14.330000 31.410000  14.400000 ;
      RECT 23.445000  14.330000 31.410000  14.400000 ;
      RECT 23.515000  14.400000 31.410000  14.470000 ;
      RECT 23.515000  14.400000 31.410000  14.470000 ;
      RECT 23.585000  14.470000 31.410000  14.540000 ;
      RECT 23.585000  14.470000 31.410000  14.540000 ;
      RECT 23.655000  14.540000 31.410000  14.610000 ;
      RECT 23.655000  14.540000 31.410000  14.610000 ;
      RECT 23.725000  14.610000 31.410000  14.680000 ;
      RECT 23.725000  14.610000 31.410000  14.680000 ;
      RECT 23.795000  14.680000 31.410000  14.750000 ;
      RECT 23.795000  14.680000 31.410000  14.750000 ;
      RECT 23.865000  14.750000 31.410000  14.820000 ;
      RECT 23.865000  14.750000 31.410000  14.820000 ;
      RECT 23.875000  25.345000 29.985000  36.515000 ;
      RECT 23.875000  36.515000 30.250000  36.780000 ;
      RECT 23.875000  36.780000 30.250000  37.685000 ;
      RECT 23.875000  37.685000 29.985000  37.950000 ;
      RECT 23.875000  37.950000 29.985000  39.095000 ;
      RECT 23.935000  14.820000 31.410000  14.890000 ;
      RECT 23.935000  14.820000 31.410000  14.890000 ;
      RECT 24.005000  14.890000 31.410000  14.960000 ;
      RECT 24.005000  14.890000 31.410000  14.960000 ;
      RECT 24.015000  25.405000 29.845000  37.630000 ;
      RECT 24.015000  36.570000 29.845000  36.640000 ;
      RECT 24.015000  36.570000 29.845000  36.640000 ;
      RECT 24.015000  36.640000 29.915000  36.710000 ;
      RECT 24.015000  36.640000 29.915000  36.710000 ;
      RECT 24.015000  36.710000 29.985000  36.780000 ;
      RECT 24.015000  36.710000 29.985000  36.780000 ;
      RECT 24.015000  36.780000 30.055000  36.835000 ;
      RECT 24.015000  36.780000 30.055000  36.835000 ;
      RECT 24.015000  36.835000 30.110000  37.245000 ;
      RECT 24.015000  37.245000 30.110000  37.630000 ;
      RECT 24.015000  37.630000 30.040000  37.700000 ;
      RECT 24.015000  37.630000 30.040000  37.700000 ;
      RECT 24.015000  37.700000 29.970000  37.770000 ;
      RECT 24.015000  37.700000 29.970000  37.770000 ;
      RECT 24.015000  37.770000 29.900000  37.840000 ;
      RECT 24.015000  37.770000 29.900000  37.840000 ;
      RECT 24.015000  37.840000 29.845000  37.895000 ;
      RECT 24.015000  37.840000 29.845000  37.895000 ;
      RECT 24.015000  37.895000 29.845000  39.235000 ;
      RECT 24.055000  15.205000 31.550000  16.005000 ;
      RECT 24.055000  16.005000 29.985000  17.570000 ;
      RECT 24.055000  17.570000 29.985000  25.165000 ;
      RECT 24.055000  25.165000 29.985000  25.345000 ;
      RECT 24.055000  25.365000 29.845000  25.405000 ;
      RECT 24.055000  25.365000 29.845000  25.405000 ;
      RECT 24.075000  14.960000 31.410000  15.030000 ;
      RECT 24.075000  14.960000 31.410000  15.030000 ;
      RECT 24.125000  25.295000 29.845000  25.365000 ;
      RECT 24.125000  25.295000 29.845000  25.365000 ;
      RECT 24.145000  15.030000 31.410000  15.100000 ;
      RECT 24.145000  15.030000 31.410000  15.100000 ;
      RECT 24.195000  15.100000 31.410000  15.150000 ;
      RECT 24.195000  15.100000 31.410000  15.150000 ;
      RECT 24.195000  15.150000 31.410000  15.950000 ;
      RECT 24.195000  15.950000 29.845000  25.225000 ;
      RECT 24.195000  15.950000 31.340000  16.020000 ;
      RECT 24.195000  15.950000 31.340000  16.020000 ;
      RECT 24.195000  16.020000 31.270000  16.090000 ;
      RECT 24.195000  16.020000 31.270000  16.090000 ;
      RECT 24.195000  16.090000 31.200000  16.160000 ;
      RECT 24.195000  16.090000 31.200000  16.160000 ;
      RECT 24.195000  16.160000 31.130000  16.230000 ;
      RECT 24.195000  16.160000 31.130000  16.230000 ;
      RECT 24.195000  16.230000 31.060000  16.300000 ;
      RECT 24.195000  16.230000 31.060000  16.300000 ;
      RECT 24.195000  16.300000 30.990000  16.370000 ;
      RECT 24.195000  16.300000 30.990000  16.370000 ;
      RECT 24.195000  16.370000 30.920000  16.440000 ;
      RECT 24.195000  16.370000 30.920000  16.440000 ;
      RECT 24.195000  16.440000 30.850000  16.510000 ;
      RECT 24.195000  16.440000 30.850000  16.510000 ;
      RECT 24.195000  16.510000 30.780000  16.580000 ;
      RECT 24.195000  16.510000 30.780000  16.580000 ;
      RECT 24.195000  16.580000 30.710000  16.650000 ;
      RECT 24.195000  16.580000 30.710000  16.650000 ;
      RECT 24.195000  16.650000 30.640000  16.720000 ;
      RECT 24.195000  16.650000 30.640000  16.720000 ;
      RECT 24.195000  16.720000 30.570000  16.790000 ;
      RECT 24.195000  16.720000 30.570000  16.790000 ;
      RECT 24.195000  16.790000 30.500000  16.860000 ;
      RECT 24.195000  16.790000 30.500000  16.860000 ;
      RECT 24.195000  16.860000 30.430000  16.930000 ;
      RECT 24.195000  16.860000 30.430000  16.930000 ;
      RECT 24.195000  16.930000 30.360000  17.000000 ;
      RECT 24.195000  16.930000 30.360000  17.000000 ;
      RECT 24.195000  17.000000 30.290000  17.070000 ;
      RECT 24.195000  17.000000 30.290000  17.070000 ;
      RECT 24.195000  17.070000 30.220000  17.140000 ;
      RECT 24.195000  17.070000 30.220000  17.140000 ;
      RECT 24.195000  17.140000 30.150000  17.210000 ;
      RECT 24.195000  17.140000 30.150000  17.210000 ;
      RECT 24.195000  17.210000 30.080000  17.280000 ;
      RECT 24.195000  17.210000 30.080000  17.280000 ;
      RECT 24.195000  17.280000 30.010000  17.350000 ;
      RECT 24.195000  17.280000 30.010000  17.350000 ;
      RECT 24.195000  17.350000 29.940000  17.420000 ;
      RECT 24.195000  17.350000 29.940000  17.420000 ;
      RECT 24.195000  17.420000 29.870000  17.490000 ;
      RECT 24.195000  17.420000 29.870000  17.490000 ;
      RECT 24.195000  17.490000 29.845000  17.515000 ;
      RECT 24.195000  17.490000 29.845000  17.515000 ;
      RECT 24.195000  17.515000 29.845000  25.225000 ;
      RECT 24.195000  25.225000 29.845000  25.295000 ;
      RECT 24.195000  25.225000 29.845000  25.295000 ;
      RECT 24.535000  57.880000 76.635000  57.920000 ;
      RECT 24.535000  57.880000 76.635000  57.920000 ;
      RECT 24.605000  57.810000 76.635000  57.880000 ;
      RECT 24.605000  57.810000 76.635000  57.880000 ;
      RECT 24.675000  57.740000 76.635000  57.810000 ;
      RECT 24.675000  57.740000 76.635000  57.810000 ;
      RECT 24.745000  57.670000 76.635000  57.740000 ;
      RECT 24.745000  57.670000 76.635000  57.740000 ;
      RECT 24.815000  57.600000 76.635000  57.670000 ;
      RECT 24.815000  57.600000 76.635000  57.670000 ;
      RECT 24.885000  57.530000 76.635000  57.600000 ;
      RECT 24.885000  57.530000 76.635000  57.600000 ;
      RECT 24.955000  57.460000 76.635000  57.530000 ;
      RECT 24.955000  57.460000 76.635000  57.530000 ;
      RECT 25.025000  57.390000 76.635000  57.460000 ;
      RECT 25.025000  57.390000 76.635000  57.460000 ;
      RECT 25.095000  53.425000 76.775000  57.125000 ;
      RECT 25.095000  57.125000 76.775000  57.780000 ;
      RECT 25.095000  57.320000 76.635000  57.390000 ;
      RECT 25.095000  57.320000 76.635000  57.390000 ;
      RECT 25.165000  57.250000 76.635000  57.320000 ;
      RECT 25.165000  57.250000 76.635000  57.320000 ;
      RECT 25.235000  53.480000 76.635000  57.180000 ;
      RECT 25.235000  53.480000 76.635000  57.920000 ;
      RECT 25.235000  53.480000 76.635000  73.500000 ;
      RECT 25.235000  57.180000 76.635000  57.250000 ;
      RECT 25.235000  57.180000 76.635000  57.250000 ;
      RECT 25.260000  53.260000 76.775000  53.425000 ;
      RECT 25.260000  53.455000 76.635000  53.480000 ;
      RECT 25.260000  53.455000 76.635000  53.480000 ;
      RECT 25.330000  53.385000 76.635000  53.455000 ;
      RECT 25.330000  53.385000 76.635000  53.455000 ;
      RECT 25.400000  53.315000 76.635000  53.385000 ;
      RECT 25.400000  53.315000 76.635000  53.385000 ;
      RECT 25.455000  53.260000 76.580000  53.315000 ;
      RECT 25.455000  53.260000 76.580000  53.315000 ;
      RECT 25.525000  53.190000 76.510000  53.260000 ;
      RECT 25.525000  53.190000 76.510000  53.260000 ;
      RECT 25.595000  53.120000 76.440000  53.190000 ;
      RECT 25.595000  53.120000 76.440000  53.190000 ;
      RECT 25.665000  53.050000 76.370000  53.120000 ;
      RECT 25.665000  53.050000 76.370000  53.120000 ;
      RECT 25.735000  52.980000 76.300000  53.050000 ;
      RECT 25.735000  52.980000 76.300000  53.050000 ;
      RECT 25.805000  52.910000 76.230000  52.980000 ;
      RECT 25.805000  52.910000 76.230000  52.980000 ;
      RECT 25.875000  52.840000 76.160000  52.910000 ;
      RECT 25.875000  52.840000 76.160000  52.910000 ;
      RECT 25.945000  52.575000 76.775000  53.260000 ;
      RECT 25.945000  52.770000 76.090000  52.840000 ;
      RECT 25.945000  52.770000 76.090000  52.840000 ;
      RECT 26.015000  52.700000 76.020000  52.770000 ;
      RECT 26.015000  52.700000 76.020000  52.770000 ;
      RECT 26.085000  52.630000 75.950000  52.700000 ;
      RECT 26.085000  52.630000 75.950000  52.700000 ;
      RECT 26.155000  52.560000 75.950000  52.630000 ;
      RECT 26.155000  52.560000 75.950000  52.630000 ;
      RECT 26.165000  52.350000 76.090000  52.575000 ;
      RECT 26.225000  52.490000 75.950000  52.560000 ;
      RECT 26.225000  52.490000 75.950000  52.560000 ;
      RECT 27.000000   0.000000 28.350000   1.835000 ;
      RECT 27.140000   0.000000 28.210000   1.975000 ;
      RECT 28.890000   0.000000 30.610000   2.320000 ;
      RECT 28.890000   2.320000 31.165000   2.880000 ;
      RECT 28.890000   2.880000 31.165000   3.900000 ;
      RECT 28.890000   3.900000 31.165000   4.505000 ;
      RECT 29.030000   0.000000 30.470000   2.380000 ;
      RECT 29.030000   2.380000 30.470000   2.450000 ;
      RECT 29.030000   2.450000 30.540000   2.520000 ;
      RECT 29.030000   2.520000 30.610000   2.590000 ;
      RECT 29.030000   2.590000 30.680000   2.660000 ;
      RECT 29.030000   2.660000 30.750000   2.730000 ;
      RECT 29.030000   2.730000 30.820000   2.800000 ;
      RECT 29.030000   2.800000 30.890000   2.870000 ;
      RECT 29.030000   2.870000 30.960000   2.935000 ;
      RECT 29.030000   2.935000 31.025000   3.845000 ;
      RECT 29.100000   3.845000 31.025000   3.915000 ;
      RECT 29.170000   3.915000 31.025000   3.985000 ;
      RECT 29.240000   3.985000 31.025000   4.055000 ;
      RECT 29.310000   4.055000 31.025000   4.125000 ;
      RECT 29.380000   4.125000 31.025000   4.195000 ;
      RECT 29.450000   4.195000 31.025000   4.265000 ;
      RECT 29.490000   4.505000 31.285000   4.620000 ;
      RECT 29.520000   4.265000 31.025000   4.335000 ;
      RECT 29.590000   4.335000 31.025000   4.405000 ;
      RECT 29.610000   4.620000 31.550000   4.890000 ;
      RECT 29.610000   4.890000 31.550000   6.920000 ;
      RECT 29.660000   4.405000 31.025000   4.475000 ;
      RECT 29.730000   4.475000 31.025000   4.545000 ;
      RECT 29.745000   4.545000 31.025000   4.560000 ;
      RECT 29.750000   4.560000 31.025000   4.565000 ;
      RECT 29.750000   4.565000 31.025000   4.635000 ;
      RECT 29.750000   4.635000 31.100000   4.705000 ;
      RECT 29.750000   4.705000 31.170000   4.775000 ;
      RECT 29.750000   4.775000 31.240000   4.845000 ;
      RECT 29.750000   4.845000 31.310000   4.915000 ;
      RECT 29.750000   4.915000 31.380000   4.945000 ;
      RECT 29.750000   4.945000 31.410000   7.060000 ;
      RECT 29.895000  52.445000 75.950000  52.490000 ;
      RECT 29.895000  52.445000 75.950000  52.490000 ;
      RECT 29.965000  52.375000 75.950000  52.445000 ;
      RECT 29.965000  52.375000 75.950000  52.445000 ;
      RECT 30.035000  52.305000 75.950000  52.375000 ;
      RECT 30.035000  52.305000 75.950000  52.375000 ;
      RECT 30.105000  52.235000 75.950000  52.305000 ;
      RECT 30.105000  52.235000 75.950000  52.305000 ;
      RECT 30.175000  52.165000 75.950000  52.235000 ;
      RECT 30.175000  52.165000 75.950000  52.235000 ;
      RECT 30.245000  52.095000 75.950000  52.165000 ;
      RECT 30.245000  52.095000 75.950000  52.165000 ;
      RECT 30.315000  52.025000 75.950000  52.095000 ;
      RECT 30.315000  52.025000 75.950000  52.095000 ;
      RECT 30.385000  51.955000 75.950000  52.025000 ;
      RECT 30.385000  51.955000 75.950000  52.025000 ;
      RECT 30.455000  51.885000 75.950000  51.955000 ;
      RECT 30.455000  51.885000 75.950000  51.955000 ;
      RECT 30.525000  17.795000 79.180000  36.285000 ;
      RECT 30.525000  36.285000 79.180000  36.550000 ;
      RECT 30.525000  38.180000 79.180000  47.610000 ;
      RECT 30.525000  47.610000 76.090000  50.700000 ;
      RECT 30.525000  50.700000 76.090000  51.620000 ;
      RECT 30.525000  51.620000 76.090000  52.350000 ;
      RECT 30.525000  51.815000 75.950000  51.885000 ;
      RECT 30.525000  51.815000 75.950000  51.885000 ;
      RECT 30.595000  51.745000 75.950000  51.815000 ;
      RECT 30.595000  51.745000 75.950000  51.815000 ;
      RECT 30.665000  17.855000 79.175000  36.230000 ;
      RECT 30.665000  38.235000 79.175000  42.955000 ;
      RECT 30.665000  42.955000 75.950000  52.490000 ;
      RECT 30.665000  42.955000 79.040000  47.555000 ;
      RECT 30.665000  47.555000 75.950000  52.490000 ;
      RECT 30.665000  47.555000 78.970000  47.625000 ;
      RECT 30.665000  47.555000 78.970000  47.625000 ;
      RECT 30.665000  47.625000 78.900000  47.695000 ;
      RECT 30.665000  47.625000 78.900000  47.695000 ;
      RECT 30.665000  47.695000 78.830000  47.765000 ;
      RECT 30.665000  47.695000 78.830000  47.765000 ;
      RECT 30.665000  47.765000 78.760000  47.835000 ;
      RECT 30.665000  47.765000 78.760000  47.835000 ;
      RECT 30.665000  47.835000 78.690000  47.905000 ;
      RECT 30.665000  47.835000 78.690000  47.905000 ;
      RECT 30.665000  47.905000 78.620000  47.975000 ;
      RECT 30.665000  47.905000 78.620000  47.975000 ;
      RECT 30.665000  47.975000 78.550000  48.045000 ;
      RECT 30.665000  47.975000 78.550000  48.045000 ;
      RECT 30.665000  48.045000 78.480000  48.115000 ;
      RECT 30.665000  48.045000 78.480000  48.115000 ;
      RECT 30.665000  48.115000 78.410000  48.185000 ;
      RECT 30.665000  48.115000 78.410000  48.185000 ;
      RECT 30.665000  48.185000 78.340000  48.255000 ;
      RECT 30.665000  48.185000 78.340000  48.255000 ;
      RECT 30.665000  48.255000 78.270000  48.325000 ;
      RECT 30.665000  48.255000 78.270000  48.325000 ;
      RECT 30.665000  48.325000 78.200000  48.395000 ;
      RECT 30.665000  48.325000 78.200000  48.395000 ;
      RECT 30.665000  48.395000 78.130000  48.465000 ;
      RECT 30.665000  48.395000 78.130000  48.465000 ;
      RECT 30.665000  48.465000 78.060000  48.535000 ;
      RECT 30.665000  48.465000 78.060000  48.535000 ;
      RECT 30.665000  48.535000 77.990000  48.605000 ;
      RECT 30.665000  48.535000 77.990000  48.605000 ;
      RECT 30.665000  48.605000 77.920000  48.675000 ;
      RECT 30.665000  48.605000 77.920000  48.675000 ;
      RECT 30.665000  48.675000 77.850000  48.745000 ;
      RECT 30.665000  48.675000 77.850000  48.745000 ;
      RECT 30.665000  48.745000 77.780000  48.815000 ;
      RECT 30.665000  48.745000 77.780000  48.815000 ;
      RECT 30.665000  48.815000 77.710000  48.885000 ;
      RECT 30.665000  48.815000 77.710000  48.885000 ;
      RECT 30.665000  48.885000 77.640000  48.955000 ;
      RECT 30.665000  48.885000 77.640000  48.955000 ;
      RECT 30.665000  48.955000 77.570000  49.025000 ;
      RECT 30.665000  48.955000 77.570000  49.025000 ;
      RECT 30.665000  49.025000 77.500000  49.095000 ;
      RECT 30.665000  49.025000 77.500000  49.095000 ;
      RECT 30.665000  49.095000 77.430000  49.165000 ;
      RECT 30.665000  49.095000 77.430000  49.165000 ;
      RECT 30.665000  49.165000 77.360000  49.235000 ;
      RECT 30.665000  49.165000 77.360000  49.235000 ;
      RECT 30.665000  49.235000 77.290000  49.305000 ;
      RECT 30.665000  49.235000 77.290000  49.305000 ;
      RECT 30.665000  49.305000 77.220000  49.375000 ;
      RECT 30.665000  49.305000 77.220000  49.375000 ;
      RECT 30.665000  49.375000 77.150000  49.445000 ;
      RECT 30.665000  49.375000 77.150000  49.445000 ;
      RECT 30.665000  49.445000 77.080000  49.515000 ;
      RECT 30.665000  49.445000 77.080000  49.515000 ;
      RECT 30.665000  49.515000 77.010000  49.585000 ;
      RECT 30.665000  49.515000 77.010000  49.585000 ;
      RECT 30.665000  49.585000 76.940000  49.655000 ;
      RECT 30.665000  49.585000 76.940000  49.655000 ;
      RECT 30.665000  49.655000 76.870000  49.725000 ;
      RECT 30.665000  49.655000 76.870000  49.725000 ;
      RECT 30.665000  49.725000 76.800000  49.795000 ;
      RECT 30.665000  49.725000 76.800000  49.795000 ;
      RECT 30.665000  49.795000 76.730000  49.865000 ;
      RECT 30.665000  49.795000 76.730000  49.865000 ;
      RECT 30.665000  49.865000 76.660000  49.935000 ;
      RECT 30.665000  49.865000 76.660000  49.935000 ;
      RECT 30.665000  49.935000 76.590000  50.005000 ;
      RECT 30.665000  49.935000 76.590000  50.005000 ;
      RECT 30.665000  50.005000 76.520000  50.075000 ;
      RECT 30.665000  50.005000 76.520000  50.075000 ;
      RECT 30.665000  50.075000 76.450000  50.145000 ;
      RECT 30.665000  50.075000 76.450000  50.145000 ;
      RECT 30.665000  50.145000 76.380000  50.215000 ;
      RECT 30.665000  50.145000 76.380000  50.215000 ;
      RECT 30.665000  50.215000 76.310000  50.285000 ;
      RECT 30.665000  50.215000 76.310000  50.285000 ;
      RECT 30.665000  50.285000 76.240000  50.355000 ;
      RECT 30.665000  50.285000 76.240000  50.355000 ;
      RECT 30.665000  50.355000 76.170000  50.425000 ;
      RECT 30.665000  50.355000 76.170000  50.425000 ;
      RECT 30.665000  50.425000 76.100000  50.495000 ;
      RECT 30.665000  50.425000 76.100000  50.495000 ;
      RECT 30.665000  50.495000 76.030000  50.565000 ;
      RECT 30.665000  50.495000 76.030000  50.565000 ;
      RECT 30.665000  50.565000 75.960000  50.635000 ;
      RECT 30.665000  50.565000 75.960000  50.635000 ;
      RECT 30.665000  50.635000 75.950000  50.645000 ;
      RECT 30.665000  50.635000 75.950000  50.645000 ;
      RECT 30.665000  50.645000 75.950000  51.675000 ;
      RECT 30.665000  51.675000 75.950000  51.745000 ;
      RECT 30.665000  51.675000 75.950000  51.745000 ;
      RECT 30.715000  17.805000 79.175000  17.855000 ;
      RECT 30.715000  17.805000 79.175000  17.855000 ;
      RECT 30.720000  38.180000 79.175000  38.235000 ;
      RECT 30.720000  38.180000 79.175000  38.235000 ;
      RECT 30.735000  36.230000 79.175000  36.300000 ;
      RECT 30.735000  36.230000 79.175000  36.300000 ;
      RECT 30.785000  17.735000 79.175000  17.805000 ;
      RECT 30.785000  17.735000 79.175000  17.805000 ;
      RECT 30.790000  36.550000 79.180000  37.915000 ;
      RECT 30.790000  37.915000 79.180000  38.180000 ;
      RECT 30.790000  38.110000 79.175000  38.180000 ;
      RECT 30.790000  38.110000 79.175000  38.180000 ;
      RECT 30.805000  36.300000 79.175000  36.370000 ;
      RECT 30.805000  36.300000 79.175000  36.370000 ;
      RECT 30.855000  17.665000 79.175000  17.735000 ;
      RECT 30.855000  17.665000 79.175000  17.735000 ;
      RECT 30.860000  38.040000 79.175000  38.110000 ;
      RECT 30.860000  38.040000 79.175000  38.110000 ;
      RECT 30.875000  36.370000 79.175000  36.440000 ;
      RECT 30.875000  36.370000 79.175000  36.440000 ;
      RECT 30.925000  17.595000 79.175000  17.665000 ;
      RECT 30.925000  17.595000 79.175000  17.665000 ;
      RECT 30.930000  17.855000 79.175000  42.955000 ;
      RECT 30.930000  36.440000 79.175000  36.495000 ;
      RECT 30.930000  36.440000 79.175000  36.495000 ;
      RECT 30.930000  37.970000 79.175000  38.040000 ;
      RECT 30.930000  37.970000 79.175000  38.040000 ;
      RECT 30.995000  17.525000 79.175000  17.595000 ;
      RECT 30.995000  17.525000 79.175000  17.595000 ;
      RECT 31.065000  17.455000 79.175000  17.525000 ;
      RECT 31.065000  17.455000 79.175000  17.525000 ;
      RECT 31.135000  17.385000 79.175000  17.455000 ;
      RECT 31.135000  17.385000 79.175000  17.455000 ;
      RECT 31.150000   0.000000 31.675000   2.095000 ;
      RECT 31.150000   2.095000 31.675000   2.620000 ;
      RECT 31.205000  17.315000 79.175000  17.385000 ;
      RECT 31.205000  17.315000 79.175000  17.385000 ;
      RECT 31.210000  17.310000 79.170000  17.315000 ;
      RECT 31.210000  17.310000 79.170000  17.315000 ;
      RECT 31.235000  17.090000 79.180000  17.795000 ;
      RECT 31.275000  17.245000 79.105000  17.310000 ;
      RECT 31.275000  17.245000 79.105000  17.310000 ;
      RECT 31.290000   0.000000 31.535000   2.040000 ;
      RECT 31.340000  17.180000 79.040000  17.245000 ;
      RECT 31.340000  17.180000 79.040000  17.245000 ;
      RECT 31.355000  17.165000 79.040000  17.180000 ;
      RECT 31.355000  17.165000 79.040000  17.180000 ;
      RECT 31.360000   2.040000 31.535000   2.110000 ;
      RECT 31.375000  17.145000 79.040000  17.165000 ;
      RECT 31.375000  17.145000 79.040000  17.165000 ;
      RECT 31.430000   2.110000 31.535000   2.180000 ;
      RECT 31.435000  17.085000 78.980000  17.145000 ;
      RECT 31.435000  17.085000 78.980000  17.145000 ;
      RECT 31.500000   2.180000 31.535000   2.250000 ;
      RECT 31.505000  17.015000 78.910000  17.085000 ;
      RECT 31.505000  17.015000 78.910000  17.085000 ;
      RECT 31.575000  16.945000 78.840000  17.015000 ;
      RECT 31.575000  16.945000 78.840000  17.015000 ;
      RECT 31.645000  16.875000 78.770000  16.945000 ;
      RECT 31.645000  16.875000 78.770000  16.945000 ;
      RECT 31.705000   4.105000 45.105000   4.275000 ;
      RECT 31.705000   4.275000 45.105000   4.660000 ;
      RECT 31.715000  16.805000 78.700000  16.875000 ;
      RECT 31.715000  16.805000 78.700000  16.875000 ;
      RECT 31.785000  16.735000 78.630000  16.805000 ;
      RECT 31.785000  16.735000 78.630000  16.805000 ;
      RECT 31.855000  16.665000 78.560000  16.735000 ;
      RECT 31.855000  16.665000 78.560000  16.735000 ;
      RECT 31.925000  16.595000 78.490000  16.665000 ;
      RECT 31.925000  16.595000 78.490000  16.665000 ;
      RECT 31.940000   4.245000 44.965000   4.315000 ;
      RECT 31.940000  16.380000 79.180000  17.090000 ;
      RECT 31.995000  16.525000 78.420000  16.595000 ;
      RECT 31.995000  16.525000 78.420000  16.595000 ;
      RECT 32.010000   4.315000 44.965000   4.385000 ;
      RECT 32.020000  16.500000 78.420000  16.525000 ;
      RECT 32.020000  16.500000 78.420000  16.525000 ;
      RECT 32.080000   4.385000 44.965000   4.455000 ;
      RECT 32.090000   4.660000 45.105000   5.145000 ;
      RECT 32.090000   5.145000 45.715000   5.760000 ;
      RECT 32.090000   5.760000 45.715000   6.920000 ;
      RECT 32.090000   6.920000 78.570000  10.110000 ;
      RECT 32.090000  10.110000 78.475000  10.205000 ;
      RECT 32.090000  10.205000 78.475000  16.235000 ;
      RECT 32.090000  16.235000 78.475000  16.380000 ;
      RECT 32.090000  16.430000 78.420000  16.500000 ;
      RECT 32.090000  16.430000 78.420000  16.500000 ;
      RECT 32.150000   4.455000 44.965000   4.525000 ;
      RECT 32.160000  16.360000 78.420000  16.430000 ;
      RECT 32.160000  16.360000 78.420000  16.430000 ;
      RECT 32.215000   0.000000 35.320000   1.840000 ;
      RECT 32.215000   1.840000 34.995000   2.165000 ;
      RECT 32.215000   2.165000 34.995000   4.025000 ;
      RECT 32.215000   4.025000 45.105000   4.105000 ;
      RECT 32.220000   4.525000 44.965000   4.595000 ;
      RECT 32.230000   4.245000 44.965000   4.605000 ;
      RECT 32.230000   4.595000 44.965000   4.605000 ;
      RECT 32.230000   4.605000 44.965000   5.205000 ;
      RECT 32.230000   5.205000 44.965000   5.275000 ;
      RECT 32.230000   5.205000 44.965000   5.275000 ;
      RECT 32.230000   5.275000 45.035000   5.345000 ;
      RECT 32.230000   5.275000 45.035000   5.345000 ;
      RECT 32.230000   5.345000 45.105000   5.415000 ;
      RECT 32.230000   5.345000 45.105000   5.415000 ;
      RECT 32.230000   5.415000 45.175000   5.485000 ;
      RECT 32.230000   5.415000 45.175000   5.485000 ;
      RECT 32.230000   5.485000 45.245000   5.555000 ;
      RECT 32.230000   5.485000 45.245000   5.555000 ;
      RECT 32.230000   5.555000 45.315000   5.625000 ;
      RECT 32.230000   5.555000 45.315000   5.625000 ;
      RECT 32.230000   5.625000 45.385000   5.695000 ;
      RECT 32.230000   5.625000 45.385000   5.695000 ;
      RECT 32.230000   5.695000 45.455000   5.765000 ;
      RECT 32.230000   5.695000 45.455000   5.765000 ;
      RECT 32.230000   5.765000 45.525000   5.815000 ;
      RECT 32.230000   5.765000 45.525000   5.815000 ;
      RECT 32.230000   5.815000 45.575000   7.060000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.430000   8.230000 ;
      RECT 32.230000   8.230000 78.430000   8.295000 ;
      RECT 32.230000   8.230000 78.430000   8.295000 ;
      RECT 32.230000   8.295000 78.495000   8.360000 ;
      RECT 32.230000   8.295000 78.495000   8.360000 ;
      RECT 32.230000   8.360000 78.560000   8.365000 ;
      RECT 32.230000   8.360000 78.560000   8.365000 ;
      RECT 32.230000   8.365000 78.565000   9.910000 ;
      RECT 32.230000   9.910000 78.500000   9.975000 ;
      RECT 32.230000   9.910000 78.500000   9.975000 ;
      RECT 32.230000   9.975000 78.435000  10.040000 ;
      RECT 32.230000   9.975000 78.435000  10.040000 ;
      RECT 32.230000  10.040000 78.430000  10.045000 ;
      RECT 32.230000  10.040000 78.430000  10.045000 ;
      RECT 32.230000  10.045000 78.430000  10.055000 ;
      RECT 32.230000  10.055000 78.425000  10.060000 ;
      RECT 32.230000  10.055000 78.425000  10.060000 ;
      RECT 32.230000  10.060000 78.420000  10.065000 ;
      RECT 32.230000  10.060000 78.420000  10.065000 ;
      RECT 32.230000  10.065000 78.420000  16.290000 ;
      RECT 32.230000  10.065000 78.420000  17.855000 ;
      RECT 32.230000  16.290000 78.420000  16.360000 ;
      RECT 32.230000  16.290000 78.420000  16.360000 ;
      RECT 32.355000   0.000000 35.180000   1.785000 ;
      RECT 32.355000   1.785000 35.110000   1.855000 ;
      RECT 32.355000   1.855000 35.040000   1.925000 ;
      RECT 32.355000   1.925000 34.970000   1.995000 ;
      RECT 32.355000   1.995000 34.900000   2.065000 ;
      RECT 32.355000   2.065000 34.855000   2.110000 ;
      RECT 32.355000   2.110000 34.855000   4.165000 ;
      RECT 32.355000   4.165000 44.965000   4.245000 ;
      RECT 35.535000   2.390000 38.250000   3.855000 ;
      RECT 35.535000   3.855000 45.105000   4.025000 ;
      RECT 35.675000   2.450000 38.110000   3.995000 ;
      RECT 35.675000   3.995000 44.965000   4.165000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.720000   2.405000 38.110000   2.450000 ;
      RECT 35.790000   2.335000 38.110000   2.405000 ;
      RECT 35.860000   0.000000 38.250000   2.070000 ;
      RECT 35.860000   2.070000 38.250000   2.390000 ;
      RECT 35.860000   2.265000 38.110000   2.335000 ;
      RECT 35.930000   2.195000 38.110000   2.265000 ;
      RECT 36.000000   0.000000 38.110000   2.125000 ;
      RECT 36.000000   2.125000 38.110000   2.195000 ;
      RECT 38.790000   0.000000 45.105000   3.855000 ;
      RECT 38.930000   0.000000 44.965000   3.995000 ;
      RECT 38.930000   0.000000 44.965000   4.605000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 45.645000   0.000000 49.715000   0.220000 ;
      RECT 45.645000   0.220000 49.450000   0.485000 ;
      RECT 45.645000   0.485000 49.450000   0.965000 ;
      RECT 45.645000   0.965000 66.400000   1.135000 ;
      RECT 45.645000   1.135000 66.400000   1.615000 ;
      RECT 45.645000   1.615000 68.135000   4.100000 ;
      RECT 45.645000   4.100000 77.010000   4.920000 ;
      RECT 45.645000   4.920000 77.010000   5.375000 ;
      RECT 45.785000   0.000000 49.310000   0.165000 ;
      RECT 45.785000   0.165000 49.310000   0.430000 ;
      RECT 45.785000   0.165000 49.505000   0.235000 ;
      RECT 45.785000   0.235000 49.435000   0.305000 ;
      RECT 45.785000   0.305000 49.365000   0.375000 ;
      RECT 45.785000   0.375000 49.310000   0.430000 ;
      RECT 45.785000   0.430000 49.310000   1.105000 ;
      RECT 45.785000   1.105000 66.260000   4.865000 ;
      RECT 45.785000   1.105000 66.260000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.240000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   4.240000 76.870000   4.865000 ;
      RECT 45.855000   4.865000 76.870000   4.935000 ;
      RECT 45.855000   4.865000 76.870000   4.935000 ;
      RECT 45.925000   4.935000 76.870000   5.005000 ;
      RECT 45.925000   4.935000 76.870000   5.005000 ;
      RECT 45.995000   5.005000 76.870000   5.075000 ;
      RECT 45.995000   5.005000 76.870000   5.075000 ;
      RECT 46.065000   5.075000 76.870000   5.145000 ;
      RECT 46.065000   5.075000 76.870000   5.145000 ;
      RECT 46.100000   5.375000 78.570000   5.530000 ;
      RECT 46.135000   5.145000 76.870000   5.215000 ;
      RECT 46.135000   5.145000 76.870000   5.215000 ;
      RECT 46.205000   5.215000 76.870000   5.285000 ;
      RECT 46.205000   5.215000 76.870000   5.285000 ;
      RECT 46.255000   5.530000 78.570000   6.920000 ;
      RECT 46.275000   5.285000 76.870000   5.355000 ;
      RECT 46.275000   5.285000 76.870000   5.355000 ;
      RECT 46.345000   5.355000 76.870000   5.425000 ;
      RECT 46.345000   5.355000 76.870000   5.425000 ;
      RECT 46.395000   5.425000 76.870000   5.475000 ;
      RECT 46.395000   5.425000 76.870000   5.475000 ;
      RECT 46.395000   5.475000 76.870000   5.515000 ;
      RECT 46.395000   5.515000 78.430000   7.060000 ;
      RECT 49.310000   0.000000 49.575000   0.165000 ;
      RECT 50.255000   0.000000 66.695000   0.240000 ;
      RECT 50.255000   0.240000 66.695000   0.485000 ;
      RECT 50.395000   0.000000 50.640000   0.185000 ;
      RECT 50.465000   0.185000 66.555000   0.255000 ;
      RECT 50.500000   0.485000 66.695000   0.840000 ;
      RECT 50.500000   0.840000 66.570000   0.965000 ;
      RECT 50.535000   0.255000 66.555000   0.325000 ;
      RECT 50.605000   0.325000 66.555000   0.395000 ;
      RECT 50.640000   0.000000 66.260000   4.865000 ;
      RECT 50.640000   0.395000 66.555000   0.430000 ;
      RECT 50.640000   0.785000 66.485000   0.855000 ;
      RECT 50.640000   0.855000 66.415000   0.925000 ;
      RECT 50.640000   0.925000 66.345000   0.995000 ;
      RECT 50.640000   0.995000 66.275000   1.065000 ;
      RECT 50.640000   1.065000 66.260000   1.080000 ;
      RECT 66.260000   0.000000 66.555000   0.185000 ;
      RECT 66.260000   0.430000 66.555000   0.785000 ;
      RECT 67.235000   0.000000 68.135000   0.870000 ;
      RECT 67.235000   0.870000 68.135000   1.135000 ;
      RECT 67.375000   0.000000 67.995000   0.815000 ;
      RECT 67.445000   0.815000 67.995000   0.885000 ;
      RECT 67.500000   1.135000 68.135000   1.615000 ;
      RECT 67.515000   0.885000 67.995000   0.955000 ;
      RECT 67.585000   0.955000 67.995000   1.025000 ;
      RECT 67.640000   1.025000 67.995000   1.080000 ;
      RECT 67.640000   1.080000 67.995000   1.755000 ;
      RECT 69.065000   0.000000 76.140000   2.110000 ;
      RECT 69.065000   2.110000 77.010000   2.985000 ;
      RECT 69.065000   2.985000 77.010000   4.100000 ;
      RECT 69.205000   0.000000 76.000000   3.005000 ;
      RECT 69.205000   2.170000 76.000000   2.240000 ;
      RECT 69.205000   2.170000 76.000000   2.240000 ;
      RECT 69.205000   2.240000 76.070000   2.310000 ;
      RECT 69.205000   2.240000 76.070000   2.310000 ;
      RECT 69.205000   2.310000 76.140000   2.380000 ;
      RECT 69.205000   2.310000 76.140000   2.380000 ;
      RECT 69.205000   2.380000 76.210000   2.450000 ;
      RECT 69.205000   2.380000 76.210000   2.450000 ;
      RECT 69.205000   2.450000 76.280000   2.520000 ;
      RECT 69.205000   2.450000 76.280000   2.520000 ;
      RECT 69.205000   2.520000 76.350000   2.590000 ;
      RECT 69.205000   2.520000 76.350000   2.590000 ;
      RECT 69.205000   2.590000 76.420000   2.660000 ;
      RECT 69.205000   2.590000 76.420000   2.660000 ;
      RECT 69.205000   2.660000 76.490000   2.730000 ;
      RECT 69.205000   2.660000 76.490000   2.730000 ;
      RECT 69.205000   2.730000 76.560000   2.800000 ;
      RECT 69.205000   2.730000 76.560000   2.800000 ;
      RECT 69.205000   2.800000 76.630000   2.870000 ;
      RECT 69.205000   2.800000 76.630000   2.870000 ;
      RECT 69.205000   2.870000 76.700000   2.940000 ;
      RECT 69.205000   2.870000 76.700000   2.940000 ;
      RECT 69.205000   2.940000 76.770000   3.010000 ;
      RECT 69.205000   2.940000 76.770000   3.010000 ;
      RECT 69.205000   3.010000 76.840000   3.040000 ;
      RECT 69.205000   3.010000 76.840000   3.040000 ;
      RECT 69.205000   3.040000 76.870000   4.240000 ;
      RECT 76.570000  50.910000 79.435000  52.365000 ;
      RECT 76.570000  52.365000 79.435000  53.050000 ;
      RECT 76.710000  50.965000 79.435000  52.310000 ;
      RECT 76.775000  50.900000 79.435000  50.965000 ;
      RECT 76.780000  52.310000 79.435000  52.380000 ;
      RECT 76.845000  50.830000 79.435000  50.900000 ;
      RECT 76.850000  52.380000 79.435000  52.450000 ;
      RECT 76.915000  50.760000 79.435000  50.830000 ;
      RECT 76.920000  52.450000 79.435000  52.520000 ;
      RECT 76.985000  50.690000 79.435000  50.760000 ;
      RECT 76.990000  52.520000 79.435000  52.590000 ;
      RECT 77.055000  50.620000 79.435000  50.690000 ;
      RECT 77.060000   0.000000 77.470000   0.925000 ;
      RECT 77.060000   0.925000 77.350000   1.045000 ;
      RECT 77.060000   1.045000 77.250000   1.565000 ;
      RECT 77.060000   1.565000 77.250000   1.605000 ;
      RECT 77.060000  52.590000 79.435000  52.660000 ;
      RECT 77.100000   1.605000 78.570000   2.535000 ;
      RECT 77.125000  50.550000 79.435000  50.620000 ;
      RECT 77.130000  52.660000 79.435000  52.730000 ;
      RECT 77.195000  50.480000 79.435000  50.550000 ;
      RECT 77.200000  52.730000 79.435000  52.800000 ;
      RECT 77.255000  53.050000 79.435000  96.135000 ;
      RECT 77.255000  96.135000 79.435000  96.280000 ;
      RECT 77.265000  50.410000 79.435000  50.480000 ;
      RECT 77.270000  52.800000 79.435000  52.870000 ;
      RECT 77.335000  50.340000 79.435000  50.410000 ;
      RECT 77.340000  52.870000 79.435000  52.940000 ;
      RECT 77.395000  52.940000 79.435000  52.995000 ;
      RECT 77.395000  52.995000 79.435000  96.080000 ;
      RECT 77.395000  96.280000 80.000000  96.365000 ;
      RECT 77.405000  50.270000 79.435000  50.340000 ;
      RECT 77.465000  96.080000 79.435000  96.150000 ;
      RECT 77.475000  50.200000 79.435000  50.270000 ;
      RECT 77.505000   1.745000 78.430000   1.815000 ;
      RECT 77.535000  96.150000 79.435000  96.220000 ;
      RECT 77.545000  50.130000 79.435000  50.200000 ;
      RECT 77.575000   1.815000 78.430000   1.885000 ;
      RECT 77.595000  96.220000 79.435000  96.280000 ;
      RECT 77.615000  50.060000 79.435000  50.130000 ;
      RECT 77.645000   1.885000 78.430000   1.955000 ;
      RECT 77.665000  96.280000 80.000000  96.350000 ;
      RECT 77.685000  49.990000 79.435000  50.060000 ;
      RECT 77.715000   1.955000 78.430000   2.025000 ;
      RECT 77.735000  96.350000 80.000000  96.420000 ;
      RECT 77.755000  49.920000 79.435000  49.990000 ;
      RECT 77.785000   2.025000 78.430000   2.095000 ;
      RECT 77.805000  96.420000 80.000000  96.490000 ;
      RECT 77.820000  96.490000 80.000000  96.505000 ;
      RECT 77.825000  49.850000 79.435000  49.920000 ;
      RECT 77.855000   2.095000 78.430000   2.165000 ;
      RECT 77.895000  49.780000 79.435000  49.850000 ;
      RECT 77.925000   2.165000 78.430000   2.235000 ;
      RECT 77.965000  49.710000 79.435000  49.780000 ;
      RECT 77.995000   2.235000 78.430000   2.305000 ;
      RECT 78.010000   0.000000 78.565000   0.815000 ;
      RECT 78.010000   0.815000 78.565000   1.045000 ;
      RECT 78.030000   2.535000 78.570000   5.375000 ;
      RECT 78.035000  49.640000 79.435000  49.710000 ;
      RECT 78.065000   2.305000 78.430000   2.375000 ;
      RECT 78.105000  49.570000 79.435000  49.640000 ;
      RECT 78.135000   2.375000 78.430000   2.445000 ;
      RECT 78.150000   0.000000 78.425000   0.760000 ;
      RECT 78.170000   2.445000 78.430000   2.480000 ;
      RECT 78.170000   2.480000 78.430000   5.515000 ;
      RECT 78.175000  49.500000 79.435000  49.570000 ;
      RECT 78.220000   0.760000 78.425000   0.830000 ;
      RECT 78.245000  49.430000 79.435000  49.500000 ;
      RECT 78.290000   0.830000 78.425000   0.900000 ;
      RECT 78.295000   0.900000 78.425000   0.905000 ;
      RECT 78.315000  49.360000 79.435000  49.430000 ;
      RECT 78.350000   1.045000 78.565000   1.275000 ;
      RECT 78.350000   1.275000 78.570000   1.280000 ;
      RECT 78.350000   1.280000 78.570000   1.605000 ;
      RECT 78.385000  49.290000 79.435000  49.360000 ;
      RECT 78.455000  49.220000 79.435000  49.290000 ;
      RECT 78.525000  49.150000 79.435000  49.220000 ;
      RECT 78.595000  49.080000 79.435000  49.150000 ;
      RECT 78.665000  49.010000 79.435000  49.080000 ;
      RECT 78.735000  48.940000 79.435000  49.010000 ;
      RECT 78.805000  48.870000 79.435000  48.940000 ;
      RECT 78.875000  48.800000 79.435000  48.870000 ;
      RECT 78.945000  10.505000 79.435000  16.185000 ;
      RECT 78.945000  16.185000 79.435000  16.675000 ;
      RECT 78.945000  48.730000 79.435000  48.800000 ;
      RECT 79.015000  48.660000 79.435000  48.730000 ;
      RECT 79.045000   0.000000 79.435000   1.065000 ;
      RECT 79.045000   1.065000 79.435000   1.070000 ;
      RECT 79.050000   1.070000 79.435000  10.400000 ;
      RECT 79.050000  10.400000 79.435000  10.505000 ;
      RECT 79.085000  10.560000 79.435000  16.130000 ;
      RECT 79.085000  48.590000 79.435000  48.660000 ;
      RECT 79.135000  10.510000 79.435000  10.560000 ;
      RECT 79.155000  16.130000 79.435000  16.200000 ;
      RECT 79.155000  48.520000 79.435000  48.590000 ;
      RECT 79.185000   0.000000 79.435000   1.010000 ;
      RECT 79.190000   1.010000 79.435000   1.015000 ;
      RECT 79.190000   1.015000 79.435000  10.455000 ;
      RECT 79.190000  10.455000 79.435000  10.510000 ;
      RECT 79.225000  16.200000 79.435000  16.270000 ;
      RECT 79.225000  48.450000 79.435000  48.520000 ;
      RECT 79.295000  16.270000 79.435000  16.340000 ;
      RECT 79.295000  48.380000 79.435000  48.450000 ;
      RECT 79.365000  16.340000 79.435000  16.410000 ;
      RECT 79.365000  48.310000 79.435000  48.380000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.100000 106.585000 ;
      RECT  0.000000 118.955000  0.100000 178.610000 ;
      RECT  0.000000 178.610000  2.960000 181.470000 ;
      RECT  0.000000 178.800000  0.150000 178.950000 ;
      RECT  0.000000 178.950000  0.300000 179.100000 ;
      RECT  0.000000 179.100000  0.450000 179.250000 ;
      RECT  0.000000 179.250000  0.600000 179.400000 ;
      RECT  0.000000 179.400000  0.750000 179.550000 ;
      RECT  0.000000 179.550000  0.900000 179.700000 ;
      RECT  0.000000 179.700000  1.050000 179.850000 ;
      RECT  0.000000 179.850000  1.200000 180.000000 ;
      RECT  0.000000 180.000000  1.350000 180.150000 ;
      RECT  0.000000 180.150000  1.500000 180.300000 ;
      RECT  0.000000 180.300000  1.650000 180.450000 ;
      RECT  0.000000 180.450000  1.800000 180.600000 ;
      RECT  0.000000 180.600000  1.950000 180.750000 ;
      RECT  0.000000 180.750000  2.100000 180.900000 ;
      RECT  0.000000 180.900000  2.250000 181.050000 ;
      RECT  0.000000 181.050000  2.400000 181.200000 ;
      RECT  0.000000 181.200000  2.550000 181.350000 ;
      RECT  0.000000 181.350000  2.700000 181.500000 ;
      RECT  0.000000 181.470000 80.000000 200.000000 ;
      RECT  0.000000 181.500000  2.850000 181.570000 ;
      RECT  0.000000 181.570000  7.970000 184.570000 ;
      RECT  0.000000 184.570000  7.965000 184.575000 ;
      RECT  0.000000 184.575000  3.005000 196.995000 ;
      RECT  0.000000 196.995000 80.000000 200.000000 ;
      RECT  1.320000   0.000000 45.565000  36.930000 ;
      RECT  1.320000  36.930000 46.275000  37.640000 ;
      RECT  1.320000  37.640000 60.310000  47.660000 ;
      RECT  1.320000  47.660000 61.410000  74.310000 ;
      RECT  1.320000  74.310000 62.735000  75.635000 ;
      RECT  1.320000  75.635000 68.390000  76.345000 ;
      RECT  1.320000  76.345000 68.390000 102.210000 ;
      RECT  1.320000 102.210000 78.280000 106.585000 ;
      RECT  1.320000 118.955000 78.280000 176.780000 ;
      RECT  1.320000 176.780000 80.000000 178.110000 ;
      RECT  1.320000 178.110000 80.000000 180.140000 ;
      RECT  1.415000   0.945000 45.465000   1.675000 ;
      RECT  1.420000   0.000000 45.465000   0.945000 ;
      RECT  1.420000   1.675000 45.465000   3.950000 ;
      RECT  1.420000   3.950000  4.425000  36.970000 ;
      RECT  1.420000  36.970000 45.465000  37.120000 ;
      RECT  1.420000  37.120000 45.615000  37.270000 ;
      RECT  1.420000  37.270000 45.765000  37.420000 ;
      RECT  1.420000  37.420000 45.915000  37.570000 ;
      RECT  1.420000  37.570000 46.065000  37.720000 ;
      RECT  1.420000  37.720000 46.215000  37.740000 ;
      RECT  1.420000  37.740000  4.425000  74.350000 ;
      RECT  1.420000  74.350000 61.310000  74.500000 ;
      RECT  1.420000  74.500000 61.460000  74.650000 ;
      RECT  1.420000  74.650000 61.610000  74.800000 ;
      RECT  1.420000  74.800000 61.760000  74.950000 ;
      RECT  1.420000  74.950000 61.910000  75.100000 ;
      RECT  1.420000  75.100000 62.060000  75.250000 ;
      RECT  1.420000  75.250000 62.210000  75.400000 ;
      RECT  1.420000  75.400000 62.360000  75.550000 ;
      RECT  1.420000  75.550000 62.510000  75.700000 ;
      RECT  1.420000  75.700000 62.660000  75.735000 ;
      RECT  1.420000  75.735000 67.640000  75.885000 ;
      RECT  1.420000  75.885000 67.790000  76.035000 ;
      RECT  1.420000  76.035000 67.940000  76.185000 ;
      RECT  1.420000  76.185000 68.090000  76.335000 ;
      RECT  1.420000  76.335000 68.240000  76.385000 ;
      RECT  1.420000  76.385000 68.290000 106.585000 ;
      RECT  1.420000 118.955000  4.460000 121.960000 ;
      RECT  1.420000 121.960000  4.425000 173.875000 ;
      RECT  1.420000 173.875000  4.475000 176.880000 ;
      RECT  1.420000 176.880000  4.475000 176.960000 ;
      RECT  1.420000 176.960000  4.555000 177.040000 ;
      RECT  1.420000 177.040000  7.970000 178.070000 ;
      RECT  1.440000 178.070000 80.000000 178.090000 ;
      RECT  1.460000 102.310000 78.180000 118.955000 ;
      RECT  1.460000 102.310000 78.180000 118.955000 ;
      RECT  1.460000 178.090000 80.000000 178.110000 ;
      RECT  1.460000 178.110000  7.970000 178.145000 ;
      RECT  1.645000 178.145000 80.000000 178.295000 ;
      RECT  1.795000 178.295000 80.000000 178.445000 ;
      RECT  1.945000 178.445000 80.000000 178.595000 ;
      RECT  2.000000 106.585000 78.280000 118.955000 ;
      RECT  2.095000 178.595000 80.000000 178.745000 ;
      RECT  2.245000 178.745000 80.000000 178.895000 ;
      RECT  2.395000 178.895000 80.000000 179.045000 ;
      RECT  2.545000 179.045000 80.000000 179.195000 ;
      RECT  2.695000 179.195000 80.000000 179.345000 ;
      RECT  2.845000 179.345000 80.000000 179.495000 ;
      RECT  2.995000 179.495000 80.000000 179.645000 ;
      RECT  3.000000 184.570000 77.000000 197.000000 ;
      RECT  3.145000 179.645000 80.000000 179.795000 ;
      RECT  3.295000 179.795000 80.000000 179.945000 ;
      RECT  3.390000 179.945000 80.000000 180.040000 ;
      RECT  4.420000   3.000000 42.465000  38.215000 ;
      RECT  4.420000  38.215000 42.465000  38.365000 ;
      RECT  4.420000  38.215000 42.465000  38.365000 ;
      RECT  4.420000  38.365000 42.615000  38.515000 ;
      RECT  4.420000  38.365000 42.615000  38.515000 ;
      RECT  4.420000  38.515000 42.765000  38.665000 ;
      RECT  4.420000  38.515000 42.765000  38.665000 ;
      RECT  4.420000  38.665000 42.915000  38.815000 ;
      RECT  4.420000  38.665000 42.915000  38.815000 ;
      RECT  4.420000  38.815000 43.065000  38.965000 ;
      RECT  4.420000  38.815000 43.065000  38.965000 ;
      RECT  4.420000  38.965000 43.215000  39.115000 ;
      RECT  4.420000  38.965000 43.215000  39.115000 ;
      RECT  4.420000  39.115000 43.365000  39.265000 ;
      RECT  4.420000  39.115000 43.365000  39.265000 ;
      RECT  4.420000  39.265000 43.515000  39.415000 ;
      RECT  4.420000  39.265000 43.515000  39.415000 ;
      RECT  4.420000  39.415000 43.665000  39.565000 ;
      RECT  4.420000  39.415000 43.665000  39.565000 ;
      RECT  4.420000  39.565000 43.815000  39.715000 ;
      RECT  4.420000  39.565000 43.815000  39.715000 ;
      RECT  4.420000  39.715000 43.965000  39.865000 ;
      RECT  4.420000  39.715000 43.965000  39.865000 ;
      RECT  4.420000  39.865000 44.115000  40.015000 ;
      RECT  4.420000  39.865000 44.115000  40.015000 ;
      RECT  4.420000  40.015000 44.265000  40.165000 ;
      RECT  4.420000  40.015000 44.265000  40.165000 ;
      RECT  4.420000  40.165000 44.415000  40.315000 ;
      RECT  4.420000  40.165000 44.415000  40.315000 ;
      RECT  4.420000  40.315000 44.565000  40.465000 ;
      RECT  4.420000  40.315000 44.565000  40.465000 ;
      RECT  4.420000  40.465000 44.715000  40.615000 ;
      RECT  4.420000  40.465000 44.715000  40.615000 ;
      RECT  4.420000  40.615000 44.865000  40.740000 ;
      RECT  4.420000  40.615000 44.865000  40.740000 ;
      RECT  4.420000  40.740000 57.210000  50.760000 ;
      RECT  4.420000  50.760000 58.310000  75.595000 ;
      RECT  4.420000  75.595000 58.310000  75.745000 ;
      RECT  4.420000  75.595000 58.310000  75.745000 ;
      RECT  4.420000  75.745000 58.460000  75.895000 ;
      RECT  4.420000  75.745000 58.460000  75.895000 ;
      RECT  4.420000  75.895000 58.610000  76.045000 ;
      RECT  4.420000  75.895000 58.610000  76.045000 ;
      RECT  4.420000  76.045000 58.760000  76.195000 ;
      RECT  4.420000  76.045000 58.760000  76.195000 ;
      RECT  4.420000  76.195000 58.910000  76.345000 ;
      RECT  4.420000  76.195000 58.910000  76.345000 ;
      RECT  4.420000  76.345000 59.060000  76.495000 ;
      RECT  4.420000  76.345000 59.060000  76.495000 ;
      RECT  4.420000  76.495000 59.210000  76.645000 ;
      RECT  4.420000  76.495000 59.210000  76.645000 ;
      RECT  4.420000  76.645000 59.360000  76.795000 ;
      RECT  4.420000  76.645000 59.360000  76.795000 ;
      RECT  4.420000  76.795000 59.510000  76.945000 ;
      RECT  4.420000  76.795000 59.510000  76.945000 ;
      RECT  4.420000  76.945000 59.660000  77.095000 ;
      RECT  4.420000  76.945000 59.660000  77.095000 ;
      RECT  4.420000  77.095000 59.810000  77.245000 ;
      RECT  4.420000  77.095000 59.810000  77.245000 ;
      RECT  4.420000  77.245000 59.960000  77.395000 ;
      RECT  4.420000  77.245000 59.960000  77.395000 ;
      RECT  4.420000  77.395000 60.110000  77.545000 ;
      RECT  4.420000  77.395000 60.110000  77.545000 ;
      RECT  4.420000  77.545000 60.260000  77.695000 ;
      RECT  4.420000  77.545000 60.260000  77.695000 ;
      RECT  4.420000  77.695000 60.410000  77.845000 ;
      RECT  4.420000  77.695000 60.410000  77.845000 ;
      RECT  4.420000  77.845000 60.560000  77.995000 ;
      RECT  4.420000  77.845000 60.560000  77.995000 ;
      RECT  4.420000  77.995000 60.710000  78.145000 ;
      RECT  4.420000  77.995000 60.710000  78.145000 ;
      RECT  4.420000  78.145000 60.860000  78.295000 ;
      RECT  4.420000  78.145000 60.860000  78.295000 ;
      RECT  4.420000  78.295000 61.010000  78.445000 ;
      RECT  4.420000  78.295000 61.010000  78.445000 ;
      RECT  4.420000  78.445000 61.160000  78.595000 ;
      RECT  4.420000  78.445000 61.160000  78.595000 ;
      RECT  4.420000  78.595000 61.310000  78.735000 ;
      RECT  4.420000  78.595000 61.310000  78.735000 ;
      RECT  4.420000  78.735000 65.285000 103.585000 ;
      RECT  4.420000 121.955000 75.175000 176.825000 ;
      RECT  4.460000 103.585000 65.285000 105.310000 ;
      RECT  4.460000 105.310000 75.175000 121.955000 ;
      RECT  4.525000 176.825000 75.175000 176.930000 ;
      RECT  4.525000 176.825000 75.175000 176.930000 ;
      RECT  4.630000 176.930000 75.175000 177.035000 ;
      RECT  4.630000 176.930000 75.175000 177.035000 ;
      RECT  4.635000 177.035000 75.175000 177.040000 ;
      RECT  4.635000 177.035000 75.175000 177.040000 ;
      RECT  4.865000 180.140000 80.000000 181.470000 ;
      RECT  4.965000 178.070000  7.970000 178.110000 ;
      RECT  4.965000 178.145000  7.970000 181.570000 ;
      RECT  7.965000 177.040000 75.175000 179.880000 ;
      RECT  7.965000 179.880000 77.000000 184.570000 ;
      RECT 42.460000   3.950000 45.465000  36.970000 ;
      RECT 42.465000  37.740000 52.000000  40.745000 ;
      RECT 46.495000   0.000000 62.520000   5.430000 ;
      RECT 46.495000   5.430000 61.960000   5.990000 ;
      RECT 46.495000   5.990000 59.300000   7.300000 ;
      RECT 46.495000   7.300000 59.300000  11.060000 ;
      RECT 46.495000  11.060000 61.170000  12.930000 ;
      RECT 46.495000  12.930000 61.170000  18.080000 ;
      RECT 46.495000  18.080000 60.310000  18.940000 ;
      RECT 46.495000  18.940000 60.310000  35.570000 ;
      RECT 46.495000  35.570000 47.660000  36.315000 ;
      RECT 46.495000  36.315000 47.880000  36.535000 ;
      RECT 46.495000  36.535000 47.880000  36.540000 ;
      RECT 46.495000  36.540000 47.880000  36.610000 ;
      RECT 46.565000  36.610000 47.780000  36.710000 ;
      RECT 46.595000   0.000000 62.420000   3.005000 ;
      RECT 46.595000   3.005000 49.600000   5.390000 ;
      RECT 46.595000   5.390000 62.270000   5.540000 ;
      RECT 46.595000   5.540000 62.120000   5.690000 ;
      RECT 46.595000   5.690000 61.970000   5.840000 ;
      RECT 46.595000   5.840000 61.920000   5.890000 ;
      RECT 46.595000   5.890000 60.420000   6.040000 ;
      RECT 46.595000   6.040000 60.270000   6.190000 ;
      RECT 46.595000   6.190000 60.120000   6.340000 ;
      RECT 46.595000   6.340000 59.970000   6.490000 ;
      RECT 46.595000   6.490000 59.820000   6.640000 ;
      RECT 46.595000   6.640000 59.670000   6.790000 ;
      RECT 46.595000   6.790000 59.520000   6.940000 ;
      RECT 46.595000   6.940000 59.370000   7.090000 ;
      RECT 46.595000   7.090000 59.220000   7.240000 ;
      RECT 46.595000   7.240000 59.200000   7.260000 ;
      RECT 46.595000   7.260000 59.200000  35.470000 ;
      RECT 46.595000  11.100000 59.200000  11.250000 ;
      RECT 46.595000  11.250000 59.350000  11.400000 ;
      RECT 46.595000  11.400000 59.500000  11.550000 ;
      RECT 46.595000  11.550000 59.650000  11.700000 ;
      RECT 46.595000  11.700000 59.800000  11.850000 ;
      RECT 46.595000  11.850000 59.950000  12.000000 ;
      RECT 46.595000  12.000000 60.100000  12.150000 ;
      RECT 46.595000  12.150000 60.250000  12.300000 ;
      RECT 46.595000  12.300000 60.400000  12.450000 ;
      RECT 46.595000  12.450000 60.550000  12.600000 ;
      RECT 46.595000  12.600000 60.700000  12.750000 ;
      RECT 46.595000  12.750000 60.850000  12.900000 ;
      RECT 46.595000  12.900000 61.000000  12.970000 ;
      RECT 46.595000  18.040000 60.920000  18.190000 ;
      RECT 46.595000  18.190000 60.770000  18.340000 ;
      RECT 46.595000  18.340000 60.620000  18.490000 ;
      RECT 46.595000  18.490000 60.470000  18.640000 ;
      RECT 46.595000  18.640000 60.320000  18.790000 ;
      RECT 46.595000  18.790000 60.210000  18.900000 ;
      RECT 46.595000  35.470000 47.560000  36.355000 ;
      RECT 46.595000  36.355000 47.560000  36.425000 ;
      RECT 46.595000  36.425000 47.630000  36.495000 ;
      RECT 46.595000  36.495000 47.700000  36.500000 ;
      RECT 46.650000  36.500000 47.705000  36.555000 ;
      RECT 46.705000  36.555000 47.760000  36.610000 ;
      RECT 48.310000  37.640000 60.210000  37.740000 ;
      RECT 48.460000  37.490000 60.210000  37.640000 ;
      RECT 48.610000  37.340000 60.210000  37.490000 ;
      RECT 48.760000  37.190000 60.210000  37.340000 ;
      RECT 48.810000  36.545000 60.310000  37.000000 ;
      RECT 48.810000  37.000000 60.310000  37.640000 ;
      RECT 48.910000  36.585000 52.145000  37.040000 ;
      RECT 48.910000  37.040000 60.210000  37.190000 ;
      RECT 49.025000  36.470000 60.210000  36.585000 ;
      RECT 49.040000  35.570000 60.310000  36.315000 ;
      RECT 49.040000  36.315000 60.310000  36.545000 ;
      RECT 49.140000  35.470000 52.145000  36.585000 ;
      RECT 49.140000  36.355000 60.210000  36.470000 ;
      RECT 49.510000  40.685000 57.210000  40.740000 ;
      RECT 49.510000  40.685000 57.210000  40.740000 ;
      RECT 49.595000   3.000000 59.065000   3.150000 ;
      RECT 49.595000   3.000000 59.065000   3.150000 ;
      RECT 49.595000   3.150000 58.915000   3.300000 ;
      RECT 49.595000   3.150000 58.915000   3.300000 ;
      RECT 49.595000   3.300000 58.765000   3.450000 ;
      RECT 49.595000   3.300000 58.765000   3.450000 ;
      RECT 49.595000   3.450000 58.615000   3.600000 ;
      RECT 49.595000   3.450000 58.615000   3.600000 ;
      RECT 49.595000   3.600000 58.465000   3.750000 ;
      RECT 49.595000   3.600000 58.465000   3.750000 ;
      RECT 49.595000   3.750000 58.315000   3.900000 ;
      RECT 49.595000   3.750000 58.315000   3.900000 ;
      RECT 49.595000   3.900000 58.165000   4.050000 ;
      RECT 49.595000   3.900000 58.165000   4.050000 ;
      RECT 49.595000   4.050000 58.015000   4.200000 ;
      RECT 49.595000   4.050000 58.015000   4.200000 ;
      RECT 49.595000   4.200000 57.865000   4.350000 ;
      RECT 49.595000   4.200000 57.865000   4.350000 ;
      RECT 49.595000   4.350000 57.715000   4.500000 ;
      RECT 49.595000   4.350000 57.715000   4.500000 ;
      RECT 49.595000   4.500000 57.565000   4.650000 ;
      RECT 49.595000   4.500000 57.565000   4.650000 ;
      RECT 49.595000   4.650000 57.415000   4.800000 ;
      RECT 49.595000   4.650000 57.415000   4.800000 ;
      RECT 49.595000   4.800000 57.265000   4.950000 ;
      RECT 49.595000   4.800000 57.265000   4.950000 ;
      RECT 49.595000   4.950000 57.115000   5.100000 ;
      RECT 49.595000   4.950000 57.115000   5.100000 ;
      RECT 49.595000   5.100000 56.965000   5.250000 ;
      RECT 49.595000   5.100000 56.965000   5.250000 ;
      RECT 49.595000   5.250000 56.815000   5.400000 ;
      RECT 49.595000   5.250000 56.815000   5.400000 ;
      RECT 49.595000   5.400000 56.665000   5.550000 ;
      RECT 49.595000   5.400000 56.665000   5.550000 ;
      RECT 49.595000   5.550000 56.515000   5.700000 ;
      RECT 49.595000   5.550000 56.515000   5.700000 ;
      RECT 49.595000   5.700000 56.365000   5.850000 ;
      RECT 49.595000   5.700000 56.365000   5.850000 ;
      RECT 49.595000   5.850000 56.215000   6.000000 ;
      RECT 49.595000   5.850000 56.215000   6.000000 ;
      RECT 49.595000   6.000000 56.200000   6.015000 ;
      RECT 49.595000   6.000000 56.200000   6.015000 ;
      RECT 49.595000   6.015000 56.200000  12.345000 ;
      RECT 49.595000  12.345000 56.200000  12.495000 ;
      RECT 49.595000  12.345000 56.200000  12.495000 ;
      RECT 49.595000  12.495000 56.350000  12.645000 ;
      RECT 49.595000  12.495000 56.350000  12.645000 ;
      RECT 49.595000  12.645000 56.500000  12.795000 ;
      RECT 49.595000  12.645000 56.500000  12.795000 ;
      RECT 49.595000  12.795000 56.650000  12.945000 ;
      RECT 49.595000  12.795000 56.650000  12.945000 ;
      RECT 49.595000  12.945000 56.800000  13.095000 ;
      RECT 49.595000  12.945000 56.800000  13.095000 ;
      RECT 49.595000  13.095000 56.950000  13.245000 ;
      RECT 49.595000  13.095000 56.950000  13.245000 ;
      RECT 49.595000  13.245000 57.100000  13.395000 ;
      RECT 49.595000  13.245000 57.100000  13.395000 ;
      RECT 49.595000  13.395000 57.250000  13.545000 ;
      RECT 49.595000  13.395000 57.250000  13.545000 ;
      RECT 49.595000  13.545000 57.400000  13.695000 ;
      RECT 49.595000  13.545000 57.400000  13.695000 ;
      RECT 49.595000  13.695000 57.550000  13.845000 ;
      RECT 49.595000  13.695000 57.550000  13.845000 ;
      RECT 49.595000  13.845000 57.700000  13.995000 ;
      RECT 49.595000  13.845000 57.700000  13.995000 ;
      RECT 49.595000  13.995000 57.850000  14.145000 ;
      RECT 49.595000  13.995000 57.850000  14.145000 ;
      RECT 49.595000  14.145000 58.000000  14.215000 ;
      RECT 49.595000  14.145000 58.000000  14.215000 ;
      RECT 49.595000  14.215000 58.070000  16.795000 ;
      RECT 49.595000  16.795000 57.920000  16.945000 ;
      RECT 49.595000  16.795000 57.920000  16.945000 ;
      RECT 49.595000  16.945000 57.770000  17.095000 ;
      RECT 49.595000  16.945000 57.770000  17.095000 ;
      RECT 49.595000  17.095000 57.620000  17.245000 ;
      RECT 49.595000  17.095000 57.620000  17.245000 ;
      RECT 49.595000  17.245000 57.470000  17.395000 ;
      RECT 49.595000  17.245000 57.470000  17.395000 ;
      RECT 49.595000  17.395000 57.320000  17.545000 ;
      RECT 49.595000  17.395000 57.320000  17.545000 ;
      RECT 49.595000  17.545000 57.210000  17.655000 ;
      RECT 49.595000  17.545000 57.210000  17.655000 ;
      RECT 49.595000  17.655000 57.210000  32.470000 ;
      RECT 49.660000  40.535000 57.210000  40.685000 ;
      RECT 49.660000  40.535000 57.210000  40.685000 ;
      RECT 49.810000  40.385000 57.210000  40.535000 ;
      RECT 49.810000  40.385000 57.210000  40.535000 ;
      RECT 49.960000  40.235000 57.210000  40.385000 ;
      RECT 49.960000  40.235000 57.210000  40.385000 ;
      RECT 50.110000  40.085000 57.210000  40.235000 ;
      RECT 50.110000  40.085000 57.210000  40.235000 ;
      RECT 50.260000  39.935000 57.210000  40.085000 ;
      RECT 50.260000  39.935000 57.210000  40.085000 ;
      RECT 50.410000  39.785000 57.210000  39.935000 ;
      RECT 50.410000  39.785000 57.210000  39.935000 ;
      RECT 50.560000  39.635000 57.210000  39.785000 ;
      RECT 50.560000  39.635000 57.210000  39.785000 ;
      RECT 50.710000  39.485000 57.210000  39.635000 ;
      RECT 50.710000  39.485000 57.210000  39.635000 ;
      RECT 50.860000  39.335000 57.210000  39.485000 ;
      RECT 50.860000  39.335000 57.210000  39.485000 ;
      RECT 51.010000  39.185000 57.210000  39.335000 ;
      RECT 51.010000  39.185000 57.210000  39.335000 ;
      RECT 51.160000  39.035000 57.210000  39.185000 ;
      RECT 51.160000  39.035000 57.210000  39.185000 ;
      RECT 51.310000  38.885000 57.210000  39.035000 ;
      RECT 51.310000  38.885000 57.210000  39.035000 ;
      RECT 51.460000  38.735000 57.210000  38.885000 ;
      RECT 51.460000  38.735000 57.210000  38.885000 ;
      RECT 51.610000  38.585000 57.210000  38.735000 ;
      RECT 51.610000  38.585000 57.210000  38.735000 ;
      RECT 51.760000  38.435000 57.210000  38.585000 ;
      RECT 51.760000  38.435000 57.210000  38.585000 ;
      RECT 51.910000  37.830000 57.210000  38.285000 ;
      RECT 51.910000  38.285000 57.210000  38.435000 ;
      RECT 51.910000  38.285000 57.210000  38.435000 ;
      RECT 52.025000  37.715000 57.210000  37.830000 ;
      RECT 52.025000  37.715000 57.210000  37.830000 ;
      RECT 52.140000  32.470000 57.210000  37.600000 ;
      RECT 52.140000  37.600000 57.210000  37.715000 ;
      RECT 52.140000  37.600000 57.210000  37.715000 ;
      RECT 56.825000   3.005000 62.420000   5.390000 ;
      RECT 57.205000  18.900000 60.210000  37.040000 ;
      RECT 57.205000  37.740000 60.210000  47.760000 ;
      RECT 57.210000  47.760000 61.310000  50.765000 ;
      RECT 58.065000  12.970000 61.070000  18.040000 ;
      RECT 58.305000  50.765000 61.310000  74.350000 ;
      RECT 60.685000   7.875000 62.520000   7.930000 ;
      RECT 60.685000   7.930000 62.520000  10.485000 ;
      RECT 60.685000  10.485000 62.520000  12.320000 ;
      RECT 60.785000   7.915000 62.365000   7.945000 ;
      RECT 60.785000   7.945000 62.395000   7.970000 ;
      RECT 60.785000   7.970000 62.420000  10.445000 ;
      RECT 60.930000   7.770000 62.220000   7.915000 ;
      RECT 60.935000  10.445000 62.420000  10.595000 ;
      RECT 61.080000   7.620000 62.070000   7.770000 ;
      RECT 61.085000  10.595000 62.420000  10.745000 ;
      RECT 61.190000   7.370000 62.465000   7.875000 ;
      RECT 61.230000   7.470000 61.920000   7.620000 ;
      RECT 61.235000  10.745000 62.420000  10.895000 ;
      RECT 61.385000  10.895000 62.420000  11.045000 ;
      RECT 61.535000  11.045000 62.420000  11.195000 ;
      RECT 61.685000  11.195000 62.420000  11.345000 ;
      RECT 61.695000  19.515000 62.325000  34.720000 ;
      RECT 61.795000  19.555000 62.225000  34.680000 ;
      RECT 61.795000  34.680000 62.075000  34.830000 ;
      RECT 61.795000  34.830000 61.925000  34.980000 ;
      RECT 61.835000  11.345000 62.420000  11.495000 ;
      RECT 61.925000  19.425000 62.225000  19.555000 ;
      RECT 61.985000  11.495000 62.420000  11.645000 ;
      RECT 62.075000  19.275000 62.225000  19.425000 ;
      RECT 62.135000  11.645000 62.420000  11.795000 ;
      RECT 62.285000  11.795000 62.420000  11.945000 ;
      RECT 63.080000  36.325000 78.280000  72.880000 ;
      RECT 63.080000  72.880000 78.280000  73.965000 ;
      RECT 63.180000  36.365000 67.095000  39.370000 ;
      RECT 63.180000  39.370000 66.185000  69.835000 ;
      RECT 63.180000  69.835000 71.940000  72.840000 ;
      RECT 63.195000  36.350000 78.180000  36.365000 ;
      RECT 63.330000  72.840000 78.180000  72.990000 ;
      RECT 63.345000  36.200000 78.180000  36.350000 ;
      RECT 63.480000  72.990000 78.180000  73.140000 ;
      RECT 63.495000  36.050000 78.180000  36.200000 ;
      RECT 63.630000  73.140000 78.180000  73.290000 ;
      RECT 63.645000  35.900000 78.180000  36.050000 ;
      RECT 63.780000  73.290000 78.180000  73.440000 ;
      RECT 63.795000  35.750000 78.180000  35.900000 ;
      RECT 63.930000  73.440000 78.180000  73.590000 ;
      RECT 63.945000  35.600000 78.180000  35.750000 ;
      RECT 63.995000  18.390000 78.280000  35.410000 ;
      RECT 63.995000  35.410000 78.280000  36.325000 ;
      RECT 64.080000  73.590000 78.180000  73.740000 ;
      RECT 64.095000  18.430000 67.290000  21.435000 ;
      RECT 64.095000  21.435000 67.100000  35.450000 ;
      RECT 64.095000  35.450000 78.180000  35.600000 ;
      RECT 64.190000   0.000000 78.280000  18.195000 ;
      RECT 64.190000  18.195000 78.280000  18.390000 ;
      RECT 64.190000  18.335000 78.180000  18.430000 ;
      RECT 64.205000  73.740000 78.180000  73.865000 ;
      RECT 64.290000   0.000000 78.180000   7.455000 ;
      RECT 64.290000   2.690000 78.180000   2.735000 ;
      RECT 64.290000   2.735000 78.225000   2.780000 ;
      RECT 64.290000   2.780000 78.270000   2.785000 ;
      RECT 64.290000   2.785000 78.180000  18.235000 ;
      RECT 64.290000  18.235000 78.180000  18.335000 ;
      RECT 66.180000  37.610000 75.175000  70.865000 ;
      RECT 66.195000  37.595000 75.175000  37.610000 ;
      RECT 66.195000  37.595000 75.175000  37.610000 ;
      RECT 66.345000  37.445000 75.175000  37.595000 ;
      RECT 66.345000  37.445000 75.175000  37.595000 ;
      RECT 66.495000  37.295000 75.175000  37.445000 ;
      RECT 66.495000  37.295000 75.175000  37.445000 ;
      RECT 66.645000  37.145000 75.175000  37.295000 ;
      RECT 66.645000  37.145000 75.175000  37.295000 ;
      RECT 66.795000  36.995000 75.175000  37.145000 ;
      RECT 66.795000  36.995000 75.175000  37.145000 ;
      RECT 66.945000  36.845000 75.175000  36.995000 ;
      RECT 66.945000  36.845000 75.175000  36.995000 ;
      RECT 67.095000  19.675000 75.175000  36.695000 ;
      RECT 67.095000  36.695000 75.175000  36.845000 ;
      RECT 67.095000  36.695000 75.175000  36.845000 ;
      RECT 67.100000  19.670000 75.175000  19.675000 ;
      RECT 67.100000  19.670000 75.175000  19.675000 ;
      RECT 67.195000  19.575000 75.175000  19.670000 ;
      RECT 67.195000  19.575000 75.175000  19.670000 ;
      RECT 67.290000   3.000000 75.175000   3.935000 ;
      RECT 67.290000   3.935000 75.175000   3.980000 ;
      RECT 67.290000   3.935000 75.175000   3.980000 ;
      RECT 67.290000   3.980000 75.225000   4.025000 ;
      RECT 67.290000   3.980000 75.225000   4.025000 ;
      RECT 67.290000   4.025000 75.270000   4.030000 ;
      RECT 67.290000   4.025000 75.270000   4.030000 ;
      RECT 67.290000   4.030000 75.270000   4.455000 ;
      RECT 67.290000   4.455000 75.175000  19.480000 ;
      RECT 67.290000  19.480000 75.175000  19.575000 ;
      RECT 67.290000  19.480000 75.175000  19.575000 ;
      RECT 68.680000  73.965000 78.280000  75.345000 ;
      RECT 68.870000  73.865000 78.180000  74.015000 ;
      RECT 69.020000  74.015000 78.180000  74.165000 ;
      RECT 69.170000  74.165000 78.180000  74.315000 ;
      RECT 69.320000  74.315000 78.180000  74.465000 ;
      RECT 69.470000  74.465000 78.180000  74.615000 ;
      RECT 69.620000  74.615000 78.180000  74.765000 ;
      RECT 69.770000  74.765000 78.180000  74.915000 ;
      RECT 69.920000  74.915000 78.180000  75.065000 ;
      RECT 70.060000  75.345000 78.280000 102.210000 ;
      RECT 70.070000  75.065000 78.180000  75.215000 ;
      RECT 70.110000  70.865000 75.175000  71.010000 ;
      RECT 70.110000  70.865000 75.175000  71.010000 ;
      RECT 70.160000  73.865000 78.180000 118.955000 ;
      RECT 70.160000  75.215000 78.180000  75.305000 ;
      RECT 70.260000  71.010000 75.175000  71.160000 ;
      RECT 70.260000  71.010000 75.175000  71.160000 ;
      RECT 70.410000  71.160000 75.175000  71.310000 ;
      RECT 70.410000  71.160000 75.175000  71.310000 ;
      RECT 70.560000  71.310000 75.175000  71.460000 ;
      RECT 70.560000  71.310000 75.175000  71.460000 ;
      RECT 70.710000  71.460000 75.175000  71.610000 ;
      RECT 70.710000  71.460000 75.175000  71.610000 ;
      RECT 70.860000  71.610000 75.175000  71.760000 ;
      RECT 70.860000  71.610000 75.175000  71.760000 ;
      RECT 71.010000  71.760000 75.175000  71.910000 ;
      RECT 71.010000  71.760000 75.175000  71.910000 ;
      RECT 71.160000  71.910000 75.175000  72.060000 ;
      RECT 71.160000  71.910000 75.175000  72.060000 ;
      RECT 71.310000  72.060000 75.175000  72.210000 ;
      RECT 71.310000  72.060000 75.175000  72.210000 ;
      RECT 71.460000  72.210000 75.175000  72.360000 ;
      RECT 71.460000  72.210000 75.175000  72.360000 ;
      RECT 71.610000  72.360000 75.175000  72.510000 ;
      RECT 71.610000  72.360000 75.175000  72.510000 ;
      RECT 71.760000  72.510000 75.175000  72.660000 ;
      RECT 71.760000  72.510000 75.175000  72.660000 ;
      RECT 71.910000  72.660000 75.175000  72.810000 ;
      RECT 71.910000  72.660000 75.175000  72.810000 ;
      RECT 72.060000  72.810000 75.175000  72.960000 ;
      RECT 72.060000  72.810000 75.175000  72.960000 ;
      RECT 72.210000  72.960000 75.175000  73.110000 ;
      RECT 72.210000  72.960000 75.175000  73.110000 ;
      RECT 72.360000  73.110000 75.175000  73.260000 ;
      RECT 72.360000  73.110000 75.175000  73.260000 ;
      RECT 72.510000  73.260000 75.175000  73.410000 ;
      RECT 72.510000  73.260000 75.175000  73.410000 ;
      RECT 72.660000  73.410000 75.175000  73.560000 ;
      RECT 72.660000  73.410000 75.175000  73.560000 ;
      RECT 72.810000  73.560000 75.175000  73.710000 ;
      RECT 72.810000  73.560000 75.175000  73.710000 ;
      RECT 72.960000  73.710000 75.175000  73.860000 ;
      RECT 72.960000  73.710000 75.175000  73.860000 ;
      RECT 73.110000  73.860000 75.175000  74.010000 ;
      RECT 73.110000  73.860000 75.175000  74.010000 ;
      RECT 73.160000  74.010000 75.175000  74.060000 ;
      RECT 73.160000  74.010000 75.175000  74.060000 ;
      RECT 73.160000  74.060000 75.175000 105.310000 ;
      RECT 75.175000  18.430000 78.180000  35.450000 ;
      RECT 75.175000  36.365000 78.180000  72.840000 ;
      RECT 75.175000 118.955000 78.180000 176.880000 ;
      RECT 75.175000 176.880000 80.000000 179.885000 ;
      RECT 75.270000   2.785000 78.275000   7.455000 ;
      RECT 76.995000 179.885000 80.000000 196.995000 ;
      RECT 78.180000   1.160000 78.190000   1.490000 ;
      RECT 79.870000   0.000000 80.000000 176.780000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000 80.000000   1.635000 ;
      RECT  0.000000   7.885000  4.675000   8.485000 ;
      RECT  0.000000   7.885000 80.000000   8.485000 ;
      RECT  0.000000  13.935000  4.675000  14.535000 ;
      RECT  0.000000  13.935000 80.000000  14.535000 ;
      RECT  0.000000  18.785000  4.675000  19.385000 ;
      RECT  0.000000  18.785000 80.000000  19.385000 ;
      RECT  0.000000  24.835000  4.675000  25.435000 ;
      RECT  0.000000  24.835000 80.000000  25.435000 ;
      RECT  0.000000  30.885000  4.675000  31.485000 ;
      RECT  0.000000  30.885000 80.000000  31.485000 ;
      RECT  0.000000  35.735000  4.675000  36.335000 ;
      RECT  0.000000  35.735000 80.000000  36.335000 ;
      RECT  0.000000  40.585000  4.675000  41.185000 ;
      RECT  0.000000  40.585000 80.000000  41.185000 ;
      RECT  0.000000  46.635000  4.675000  47.335000 ;
      RECT  0.000000  46.635000 80.000000  47.435000 ;
      RECT  0.000000  57.035000 80.000000  57.835000 ;
      RECT  0.000000  57.135000  4.675000  57.835000 ;
      RECT  0.000000  63.085000  4.675000  63.685000 ;
      RECT  0.000000  63.085000 80.000000  63.685000 ;
      RECT  0.000000  68.935000  4.675000  69.635000 ;
      RECT  0.000000  68.935000 80.000000  69.635000 ;
      RECT  0.000000  95.400000  3.005000 104.215000 ;
      RECT  0.000000  95.400000 80.000000 104.315000 ;
      RECT  0.000000 104.215000  9.485000 104.365000 ;
      RECT  0.000000 104.315000  7.705000 106.285000 ;
      RECT  0.000000 104.365000  9.335000 104.515000 ;
      RECT  0.000000 104.515000  9.185000 104.665000 ;
      RECT  0.000000 104.665000  9.035000 104.815000 ;
      RECT  0.000000 104.815000  8.885000 104.965000 ;
      RECT  0.000000 104.965000  8.735000 105.115000 ;
      RECT  0.000000 105.115000  8.585000 105.265000 ;
      RECT  0.000000 105.265000  8.435000 105.415000 ;
      RECT  0.000000 105.415000  8.285000 105.565000 ;
      RECT  0.000000 105.565000  8.135000 105.715000 ;
      RECT  0.000000 105.715000  7.985000 105.865000 ;
      RECT  0.000000 105.865000  7.835000 106.015000 ;
      RECT  0.000000 106.015000  7.685000 106.165000 ;
      RECT  0.000000 106.165000  7.665000 106.185000 ;
      RECT  0.000000 106.185000  1.600000 106.585000 ;
      RECT  0.000000 106.285000  1.700000 106.585000 ;
      RECT  0.000000 118.955000  1.600000 119.355000 ;
      RECT  0.000000 118.955000  1.700000 119.255000 ;
      RECT  0.000000 119.255000  9.685000 121.550000 ;
      RECT  0.000000 119.355000  7.350000 119.505000 ;
      RECT  0.000000 119.505000  7.500000 119.655000 ;
      RECT  0.000000 119.655000  7.650000 119.805000 ;
      RECT  0.000000 119.805000  7.800000 119.955000 ;
      RECT  0.000000 119.955000  7.950000 120.105000 ;
      RECT  0.000000 120.105000  8.100000 120.255000 ;
      RECT  0.000000 120.255000  8.250000 120.405000 ;
      RECT  0.000000 120.405000  8.400000 120.555000 ;
      RECT  0.000000 120.555000  8.550000 120.705000 ;
      RECT  0.000000 120.705000  8.700000 120.855000 ;
      RECT  0.000000 120.855000  8.850000 121.005000 ;
      RECT  0.000000 121.005000  9.000000 121.155000 ;
      RECT  0.000000 121.155000  9.150000 121.305000 ;
      RECT  0.000000 121.305000  9.300000 121.455000 ;
      RECT  0.000000 121.455000  9.450000 121.605000 ;
      RECT  0.000000 121.550000 80.000000 175.385000 ;
      RECT  0.000000 121.605000  9.600000 121.650000 ;
      RECT  0.000000 121.650000 15.900000 124.655000 ;
      RECT  0.000000 124.655000  3.005000 172.380000 ;
      RECT  0.000000 172.380000  4.670000 175.385000 ;
      RECT  1.365000  14.535000  4.675000  18.785000 ;
      RECT  1.365000  14.535000 78.635000  18.785000 ;
      RECT  1.455000  70.310000  4.675000  94.885000 ;
      RECT  1.570000  47.435000 78.430000  57.035000 ;
      RECT  1.670000   1.635000 78.330000   4.640000 ;
      RECT  1.670000   1.635000 78.330000   7.885000 ;
      RECT  1.670000   4.640000  4.675000   7.885000 ;
      RECT  1.670000   8.485000  4.675000  13.935000 ;
      RECT  1.670000   8.485000 78.330000  13.935000 ;
      RECT  1.670000  19.385000  4.675000  24.835000 ;
      RECT  1.670000  19.385000 78.330000  24.835000 ;
      RECT  1.670000  25.435000  4.675000  30.885000 ;
      RECT  1.670000  25.435000 78.330000  30.885000 ;
      RECT  1.670000  31.485000  4.675000  35.735000 ;
      RECT  1.670000  31.485000 78.330000  35.735000 ;
      RECT  1.670000  36.335000  4.675000  40.585000 ;
      RECT  1.670000  36.335000 78.330000  40.585000 ;
      RECT  1.670000  41.185000  4.675000  46.635000 ;
      RECT  1.670000  41.185000 78.330000  46.635000 ;
      RECT  1.670000  47.335000  4.675000  57.135000 ;
      RECT  1.670000  57.835000  4.675000  63.085000 ;
      RECT  1.670000  57.835000 78.330000  63.085000 ;
      RECT  1.670000  63.685000  4.675000  68.935000 ;
      RECT  1.670000  63.685000 78.330000  68.935000 ;
      RECT  1.670000  69.635000  4.675000  70.310000 ;
      RECT  1.670000  69.635000 78.330000  95.400000 ;
      RECT  1.670000  94.885000 78.330000 104.215000 ;
      RECT  1.670000 175.385000  4.675000 196.995000 ;
      RECT  1.670000 175.385000 78.330000 200.000000 ;
      RECT  1.670000 196.995000 78.330000 200.000000 ;
      RECT  3.000000  98.400000 77.000000 101.210000 ;
      RECT  3.000000 101.210000  8.245000 101.360000 ;
      RECT  3.000000 101.210000  8.245000 101.360000 ;
      RECT  3.000000 101.360000  8.095000 101.510000 ;
      RECT  3.000000 101.360000  8.095000 101.510000 ;
      RECT  3.000000 101.510000  7.940000 101.660000 ;
      RECT  3.000000 101.510000  7.940000 101.660000 ;
      RECT  3.000000 101.660000  7.795000 101.810000 ;
      RECT  3.000000 101.660000  7.795000 101.810000 ;
      RECT  3.000000 101.810000  7.645000 101.960000 ;
      RECT  3.000000 101.810000  7.645000 101.960000 ;
      RECT  3.000000 101.960000  7.495000 102.110000 ;
      RECT  3.000000 101.960000  7.495000 102.110000 ;
      RECT  3.000000 102.110000  7.345000 102.260000 ;
      RECT  3.000000 102.110000  7.345000 102.260000 ;
      RECT  3.000000 102.260000  7.190000 102.410000 ;
      RECT  3.000000 102.260000  7.190000 102.410000 ;
      RECT  3.000000 102.410000  7.045000 102.560000 ;
      RECT  3.000000 102.410000  7.045000 102.560000 ;
      RECT  3.000000 102.560000  6.895000 102.710000 ;
      RECT  3.000000 102.560000  6.895000 102.710000 ;
      RECT  3.000000 102.710000  6.745000 102.860000 ;
      RECT  3.000000 102.710000  6.745000 102.860000 ;
      RECT  3.000000 102.860000  6.595000 103.010000 ;
      RECT  3.000000 102.860000  6.595000 103.010000 ;
      RECT  3.000000 103.010000  6.440000 103.160000 ;
      RECT  3.000000 103.010000  6.440000 103.160000 ;
      RECT  3.000000 103.160000  6.420000 103.185000 ;
      RECT  3.000000 103.160000  6.420000 103.185000 ;
      RECT  3.000000 122.355000  6.105000 122.505000 ;
      RECT  3.000000 122.355000  6.105000 122.505000 ;
      RECT  3.000000 122.505000  6.255000 122.655000 ;
      RECT  3.000000 122.505000  6.255000 122.655000 ;
      RECT  3.000000 122.655000  6.400000 122.805000 ;
      RECT  3.000000 122.655000  6.400000 122.805000 ;
      RECT  3.000000 122.805000  6.555000 122.955000 ;
      RECT  3.000000 122.805000  6.555000 122.955000 ;
      RECT  3.000000 122.955000  6.705000 123.105000 ;
      RECT  3.000000 122.955000  6.705000 123.105000 ;
      RECT  3.000000 123.105000  6.850000 123.255000 ;
      RECT  3.000000 123.105000  6.850000 123.255000 ;
      RECT  3.000000 123.255000  7.005000 123.405000 ;
      RECT  3.000000 123.255000  7.005000 123.405000 ;
      RECT  3.000000 123.405000  7.150000 123.555000 ;
      RECT  3.000000 123.405000  7.150000 123.555000 ;
      RECT  3.000000 123.555000  7.305000 123.705000 ;
      RECT  3.000000 123.555000  7.305000 123.705000 ;
      RECT  3.000000 123.705000  7.455000 123.855000 ;
      RECT  3.000000 123.705000  7.455000 123.855000 ;
      RECT  3.000000 123.855000  7.600000 124.005000 ;
      RECT  3.000000 123.855000  7.600000 124.005000 ;
      RECT  3.000000 124.005000  7.755000 124.155000 ;
      RECT  3.000000 124.005000  7.755000 124.155000 ;
      RECT  3.000000 124.155000  7.900000 124.305000 ;
      RECT  3.000000 124.155000  7.900000 124.305000 ;
      RECT  3.000000 124.305000  8.055000 124.455000 ;
      RECT  3.000000 124.305000  8.055000 124.455000 ;
      RECT  3.000000 124.455000  8.205000 124.605000 ;
      RECT  3.000000 124.455000  8.205000 124.605000 ;
      RECT  3.000000 124.605000  8.355000 124.650000 ;
      RECT  3.000000 124.605000  8.355000 124.650000 ;
      RECT  3.000000 124.650000 77.000000 172.385000 ;
      RECT  4.455000  73.310000 75.330000  91.880000 ;
      RECT  4.670000   3.000000 75.330000  73.310000 ;
      RECT  4.670000  91.880000 75.330000  98.400000 ;
      RECT  4.670000 172.385000 75.330000 197.000000 ;
      RECT  9.880000 121.400000 12.460000 121.650000 ;
      RECT 12.800000 104.315000 80.000000 121.550000 ;
      RECT 12.900000  95.400000 80.000000 121.650000 ;
      RECT 15.900000 101.210000 77.000000 124.650000 ;
      RECT 75.325000   4.640000 78.330000   7.885000 ;
      RECT 75.325000   7.885000 80.000000   8.485000 ;
      RECT 75.325000   8.485000 78.330000  13.935000 ;
      RECT 75.325000  13.935000 80.000000  14.535000 ;
      RECT 75.325000  14.535000 78.635000  18.785000 ;
      RECT 75.325000  18.785000 80.000000  19.385000 ;
      RECT 75.325000  19.385000 78.330000  24.835000 ;
      RECT 75.325000  24.835000 80.000000  25.435000 ;
      RECT 75.325000  25.435000 78.330000  30.885000 ;
      RECT 75.325000  30.885000 80.000000  31.485000 ;
      RECT 75.325000  31.485000 78.330000  35.735000 ;
      RECT 75.325000  35.735000 80.000000  36.335000 ;
      RECT 75.325000  36.335000 78.330000  40.585000 ;
      RECT 75.325000  40.585000 80.000000  41.185000 ;
      RECT 75.325000  41.185000 78.330000  46.635000 ;
      RECT 75.325000  46.635000 80.000000  47.335000 ;
      RECT 75.325000  47.335000 78.330000  57.135000 ;
      RECT 75.325000  57.135000 80.000000  57.835000 ;
      RECT 75.325000  57.835000 78.330000  63.085000 ;
      RECT 75.325000  63.085000 80.000000  63.685000 ;
      RECT 75.325000  63.685000 78.330000  68.935000 ;
      RECT 75.325000  68.935000 80.000000  69.635000 ;
      RECT 75.325000  69.635000 78.330000  94.885000 ;
      RECT 75.325000 175.385000 78.330000 196.995000 ;
      RECT 75.330000 172.380000 80.000000 175.385000 ;
      RECT 76.995000 121.650000 80.000000 172.380000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000 80.000000 106.585000 ;
      RECT  0.000000 118.955000 80.000000 124.670000 ;
      RECT  0.000000 124.670000 31.315000 147.815000 ;
      RECT  0.000000 147.815000 80.000000 200.000000 ;
      RECT  2.000000 106.585000 80.000000 118.955000 ;
      RECT 54.455000 124.670000 80.000000 147.815000 ;
  END
END sky130_fd_io__top_gpiov2


MACRO sky130_fd_io__overlay_vssd_lvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.500000 39.590000 24.500000 44.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 39.590000 74.700000 44.230000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 24.475000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.590000 39.660000  0.790000 39.860000 ;
        RECT  0.590000 40.090000  0.790000 40.290000 ;
        RECT  0.590000 40.520000  0.790000 40.720000 ;
        RECT  0.590000 40.950000  0.790000 41.150000 ;
        RECT  0.590000 41.380000  0.790000 41.580000 ;
        RECT  0.590000 41.810000  0.790000 42.010000 ;
        RECT  0.590000 42.240000  0.790000 42.440000 ;
        RECT  0.590000 42.670000  0.790000 42.870000 ;
        RECT  0.590000 43.100000  0.790000 43.300000 ;
        RECT  0.590000 43.530000  0.790000 43.730000 ;
        RECT  0.590000 43.960000  0.790000 44.160000 ;
        RECT  0.995000 39.660000  1.195000 39.860000 ;
        RECT  0.995000 40.090000  1.195000 40.290000 ;
        RECT  0.995000 40.520000  1.195000 40.720000 ;
        RECT  0.995000 40.950000  1.195000 41.150000 ;
        RECT  0.995000 41.380000  1.195000 41.580000 ;
        RECT  0.995000 41.810000  1.195000 42.010000 ;
        RECT  0.995000 42.240000  1.195000 42.440000 ;
        RECT  0.995000 42.670000  1.195000 42.870000 ;
        RECT  0.995000 43.100000  1.195000 43.300000 ;
        RECT  0.995000 43.530000  1.195000 43.730000 ;
        RECT  0.995000 43.960000  1.195000 44.160000 ;
        RECT  1.400000 39.660000  1.600000 39.860000 ;
        RECT  1.400000 40.090000  1.600000 40.290000 ;
        RECT  1.400000 40.520000  1.600000 40.720000 ;
        RECT  1.400000 40.950000  1.600000 41.150000 ;
        RECT  1.400000 41.380000  1.600000 41.580000 ;
        RECT  1.400000 41.810000  1.600000 42.010000 ;
        RECT  1.400000 42.240000  1.600000 42.440000 ;
        RECT  1.400000 42.670000  1.600000 42.870000 ;
        RECT  1.400000 43.100000  1.600000 43.300000 ;
        RECT  1.400000 43.530000  1.600000 43.730000 ;
        RECT  1.400000 43.960000  1.600000 44.160000 ;
        RECT  1.805000 39.660000  2.005000 39.860000 ;
        RECT  1.805000 40.090000  2.005000 40.290000 ;
        RECT  1.805000 40.520000  2.005000 40.720000 ;
        RECT  1.805000 40.950000  2.005000 41.150000 ;
        RECT  1.805000 41.380000  2.005000 41.580000 ;
        RECT  1.805000 41.810000  2.005000 42.010000 ;
        RECT  1.805000 42.240000  2.005000 42.440000 ;
        RECT  1.805000 42.670000  2.005000 42.870000 ;
        RECT  1.805000 43.100000  2.005000 43.300000 ;
        RECT  1.805000 43.530000  2.005000 43.730000 ;
        RECT  1.805000 43.960000  2.005000 44.160000 ;
        RECT  2.210000 39.660000  2.410000 39.860000 ;
        RECT  2.210000 40.090000  2.410000 40.290000 ;
        RECT  2.210000 40.520000  2.410000 40.720000 ;
        RECT  2.210000 40.950000  2.410000 41.150000 ;
        RECT  2.210000 41.380000  2.410000 41.580000 ;
        RECT  2.210000 41.810000  2.410000 42.010000 ;
        RECT  2.210000 42.240000  2.410000 42.440000 ;
        RECT  2.210000 42.670000  2.410000 42.870000 ;
        RECT  2.210000 43.100000  2.410000 43.300000 ;
        RECT  2.210000 43.530000  2.410000 43.730000 ;
        RECT  2.210000 43.960000  2.410000 44.160000 ;
        RECT  2.610000 39.660000  2.810000 39.860000 ;
        RECT  2.610000 40.090000  2.810000 40.290000 ;
        RECT  2.610000 40.520000  2.810000 40.720000 ;
        RECT  2.610000 40.950000  2.810000 41.150000 ;
        RECT  2.610000 41.380000  2.810000 41.580000 ;
        RECT  2.610000 41.810000  2.810000 42.010000 ;
        RECT  2.610000 42.240000  2.810000 42.440000 ;
        RECT  2.610000 42.670000  2.810000 42.870000 ;
        RECT  2.610000 43.100000  2.810000 43.300000 ;
        RECT  2.610000 43.530000  2.810000 43.730000 ;
        RECT  2.610000 43.960000  2.810000 44.160000 ;
        RECT  3.010000 39.660000  3.210000 39.860000 ;
        RECT  3.010000 40.090000  3.210000 40.290000 ;
        RECT  3.010000 40.520000  3.210000 40.720000 ;
        RECT  3.010000 40.950000  3.210000 41.150000 ;
        RECT  3.010000 41.380000  3.210000 41.580000 ;
        RECT  3.010000 41.810000  3.210000 42.010000 ;
        RECT  3.010000 42.240000  3.210000 42.440000 ;
        RECT  3.010000 42.670000  3.210000 42.870000 ;
        RECT  3.010000 43.100000  3.210000 43.300000 ;
        RECT  3.010000 43.530000  3.210000 43.730000 ;
        RECT  3.010000 43.960000  3.210000 44.160000 ;
        RECT  3.410000 39.660000  3.610000 39.860000 ;
        RECT  3.410000 40.090000  3.610000 40.290000 ;
        RECT  3.410000 40.520000  3.610000 40.720000 ;
        RECT  3.410000 40.950000  3.610000 41.150000 ;
        RECT  3.410000 41.380000  3.610000 41.580000 ;
        RECT  3.410000 41.810000  3.610000 42.010000 ;
        RECT  3.410000 42.240000  3.610000 42.440000 ;
        RECT  3.410000 42.670000  3.610000 42.870000 ;
        RECT  3.410000 43.100000  3.610000 43.300000 ;
        RECT  3.410000 43.530000  3.610000 43.730000 ;
        RECT  3.410000 43.960000  3.610000 44.160000 ;
        RECT  3.810000 39.660000  4.010000 39.860000 ;
        RECT  3.810000 40.090000  4.010000 40.290000 ;
        RECT  3.810000 40.520000  4.010000 40.720000 ;
        RECT  3.810000 40.950000  4.010000 41.150000 ;
        RECT  3.810000 41.380000  4.010000 41.580000 ;
        RECT  3.810000 41.810000  4.010000 42.010000 ;
        RECT  3.810000 42.240000  4.010000 42.440000 ;
        RECT  3.810000 42.670000  4.010000 42.870000 ;
        RECT  3.810000 43.100000  4.010000 43.300000 ;
        RECT  3.810000 43.530000  4.010000 43.730000 ;
        RECT  3.810000 43.960000  4.010000 44.160000 ;
        RECT  4.210000 39.660000  4.410000 39.860000 ;
        RECT  4.210000 40.090000  4.410000 40.290000 ;
        RECT  4.210000 40.520000  4.410000 40.720000 ;
        RECT  4.210000 40.950000  4.410000 41.150000 ;
        RECT  4.210000 41.380000  4.410000 41.580000 ;
        RECT  4.210000 41.810000  4.410000 42.010000 ;
        RECT  4.210000 42.240000  4.410000 42.440000 ;
        RECT  4.210000 42.670000  4.410000 42.870000 ;
        RECT  4.210000 43.100000  4.410000 43.300000 ;
        RECT  4.210000 43.530000  4.410000 43.730000 ;
        RECT  4.210000 43.960000  4.410000 44.160000 ;
        RECT  4.610000 39.660000  4.810000 39.860000 ;
        RECT  4.610000 40.090000  4.810000 40.290000 ;
        RECT  4.610000 40.520000  4.810000 40.720000 ;
        RECT  4.610000 40.950000  4.810000 41.150000 ;
        RECT  4.610000 41.380000  4.810000 41.580000 ;
        RECT  4.610000 41.810000  4.810000 42.010000 ;
        RECT  4.610000 42.240000  4.810000 42.440000 ;
        RECT  4.610000 42.670000  4.810000 42.870000 ;
        RECT  4.610000 43.100000  4.810000 43.300000 ;
        RECT  4.610000 43.530000  4.810000 43.730000 ;
        RECT  4.610000 43.960000  4.810000 44.160000 ;
        RECT  5.010000 39.660000  5.210000 39.860000 ;
        RECT  5.010000 40.090000  5.210000 40.290000 ;
        RECT  5.010000 40.520000  5.210000 40.720000 ;
        RECT  5.010000 40.950000  5.210000 41.150000 ;
        RECT  5.010000 41.380000  5.210000 41.580000 ;
        RECT  5.010000 41.810000  5.210000 42.010000 ;
        RECT  5.010000 42.240000  5.210000 42.440000 ;
        RECT  5.010000 42.670000  5.210000 42.870000 ;
        RECT  5.010000 43.100000  5.210000 43.300000 ;
        RECT  5.010000 43.530000  5.210000 43.730000 ;
        RECT  5.010000 43.960000  5.210000 44.160000 ;
        RECT  5.410000 39.660000  5.610000 39.860000 ;
        RECT  5.410000 40.090000  5.610000 40.290000 ;
        RECT  5.410000 40.520000  5.610000 40.720000 ;
        RECT  5.410000 40.950000  5.610000 41.150000 ;
        RECT  5.410000 41.380000  5.610000 41.580000 ;
        RECT  5.410000 41.810000  5.610000 42.010000 ;
        RECT  5.410000 42.240000  5.610000 42.440000 ;
        RECT  5.410000 42.670000  5.610000 42.870000 ;
        RECT  5.410000 43.100000  5.610000 43.300000 ;
        RECT  5.410000 43.530000  5.610000 43.730000 ;
        RECT  5.410000 43.960000  5.610000 44.160000 ;
        RECT  5.810000 39.660000  6.010000 39.860000 ;
        RECT  5.810000 40.090000  6.010000 40.290000 ;
        RECT  5.810000 40.520000  6.010000 40.720000 ;
        RECT  5.810000 40.950000  6.010000 41.150000 ;
        RECT  5.810000 41.380000  6.010000 41.580000 ;
        RECT  5.810000 41.810000  6.010000 42.010000 ;
        RECT  5.810000 42.240000  6.010000 42.440000 ;
        RECT  5.810000 42.670000  6.010000 42.870000 ;
        RECT  5.810000 43.100000  6.010000 43.300000 ;
        RECT  5.810000 43.530000  6.010000 43.730000 ;
        RECT  5.810000 43.960000  6.010000 44.160000 ;
        RECT  6.210000 39.660000  6.410000 39.860000 ;
        RECT  6.210000 40.090000  6.410000 40.290000 ;
        RECT  6.210000 40.520000  6.410000 40.720000 ;
        RECT  6.210000 40.950000  6.410000 41.150000 ;
        RECT  6.210000 41.380000  6.410000 41.580000 ;
        RECT  6.210000 41.810000  6.410000 42.010000 ;
        RECT  6.210000 42.240000  6.410000 42.440000 ;
        RECT  6.210000 42.670000  6.410000 42.870000 ;
        RECT  6.210000 43.100000  6.410000 43.300000 ;
        RECT  6.210000 43.530000  6.410000 43.730000 ;
        RECT  6.210000 43.960000  6.410000 44.160000 ;
        RECT  6.610000 39.660000  6.810000 39.860000 ;
        RECT  6.610000 40.090000  6.810000 40.290000 ;
        RECT  6.610000 40.520000  6.810000 40.720000 ;
        RECT  6.610000 40.950000  6.810000 41.150000 ;
        RECT  6.610000 41.380000  6.810000 41.580000 ;
        RECT  6.610000 41.810000  6.810000 42.010000 ;
        RECT  6.610000 42.240000  6.810000 42.440000 ;
        RECT  6.610000 42.670000  6.810000 42.870000 ;
        RECT  6.610000 43.100000  6.810000 43.300000 ;
        RECT  6.610000 43.530000  6.810000 43.730000 ;
        RECT  6.610000 43.960000  6.810000 44.160000 ;
        RECT  7.010000 39.660000  7.210000 39.860000 ;
        RECT  7.010000 40.090000  7.210000 40.290000 ;
        RECT  7.010000 40.520000  7.210000 40.720000 ;
        RECT  7.010000 40.950000  7.210000 41.150000 ;
        RECT  7.010000 41.380000  7.210000 41.580000 ;
        RECT  7.010000 41.810000  7.210000 42.010000 ;
        RECT  7.010000 42.240000  7.210000 42.440000 ;
        RECT  7.010000 42.670000  7.210000 42.870000 ;
        RECT  7.010000 43.100000  7.210000 43.300000 ;
        RECT  7.010000 43.530000  7.210000 43.730000 ;
        RECT  7.010000 43.960000  7.210000 44.160000 ;
        RECT  7.410000 39.660000  7.610000 39.860000 ;
        RECT  7.410000 40.090000  7.610000 40.290000 ;
        RECT  7.410000 40.520000  7.610000 40.720000 ;
        RECT  7.410000 40.950000  7.610000 41.150000 ;
        RECT  7.410000 41.380000  7.610000 41.580000 ;
        RECT  7.410000 41.810000  7.610000 42.010000 ;
        RECT  7.410000 42.240000  7.610000 42.440000 ;
        RECT  7.410000 42.670000  7.610000 42.870000 ;
        RECT  7.410000 43.100000  7.610000 43.300000 ;
        RECT  7.410000 43.530000  7.610000 43.730000 ;
        RECT  7.410000 43.960000  7.610000 44.160000 ;
        RECT  7.810000 39.660000  8.010000 39.860000 ;
        RECT  7.810000 40.090000  8.010000 40.290000 ;
        RECT  7.810000 40.520000  8.010000 40.720000 ;
        RECT  7.810000 40.950000  8.010000 41.150000 ;
        RECT  7.810000 41.380000  8.010000 41.580000 ;
        RECT  7.810000 41.810000  8.010000 42.010000 ;
        RECT  7.810000 42.240000  8.010000 42.440000 ;
        RECT  7.810000 42.670000  8.010000 42.870000 ;
        RECT  7.810000 43.100000  8.010000 43.300000 ;
        RECT  7.810000 43.530000  8.010000 43.730000 ;
        RECT  7.810000 43.960000  8.010000 44.160000 ;
        RECT  8.210000 39.660000  8.410000 39.860000 ;
        RECT  8.210000 40.090000  8.410000 40.290000 ;
        RECT  8.210000 40.520000  8.410000 40.720000 ;
        RECT  8.210000 40.950000  8.410000 41.150000 ;
        RECT  8.210000 41.380000  8.410000 41.580000 ;
        RECT  8.210000 41.810000  8.410000 42.010000 ;
        RECT  8.210000 42.240000  8.410000 42.440000 ;
        RECT  8.210000 42.670000  8.410000 42.870000 ;
        RECT  8.210000 43.100000  8.410000 43.300000 ;
        RECT  8.210000 43.530000  8.410000 43.730000 ;
        RECT  8.210000 43.960000  8.410000 44.160000 ;
        RECT  8.610000 39.660000  8.810000 39.860000 ;
        RECT  8.610000 40.090000  8.810000 40.290000 ;
        RECT  8.610000 40.520000  8.810000 40.720000 ;
        RECT  8.610000 40.950000  8.810000 41.150000 ;
        RECT  8.610000 41.380000  8.810000 41.580000 ;
        RECT  8.610000 41.810000  8.810000 42.010000 ;
        RECT  8.610000 42.240000  8.810000 42.440000 ;
        RECT  8.610000 42.670000  8.810000 42.870000 ;
        RECT  8.610000 43.100000  8.810000 43.300000 ;
        RECT  8.610000 43.530000  8.810000 43.730000 ;
        RECT  8.610000 43.960000  8.810000 44.160000 ;
        RECT  9.010000 39.660000  9.210000 39.860000 ;
        RECT  9.010000 40.090000  9.210000 40.290000 ;
        RECT  9.010000 40.520000  9.210000 40.720000 ;
        RECT  9.010000 40.950000  9.210000 41.150000 ;
        RECT  9.010000 41.380000  9.210000 41.580000 ;
        RECT  9.010000 41.810000  9.210000 42.010000 ;
        RECT  9.010000 42.240000  9.210000 42.440000 ;
        RECT  9.010000 42.670000  9.210000 42.870000 ;
        RECT  9.010000 43.100000  9.210000 43.300000 ;
        RECT  9.010000 43.530000  9.210000 43.730000 ;
        RECT  9.010000 43.960000  9.210000 44.160000 ;
        RECT  9.410000 39.660000  9.610000 39.860000 ;
        RECT  9.410000 40.090000  9.610000 40.290000 ;
        RECT  9.410000 40.520000  9.610000 40.720000 ;
        RECT  9.410000 40.950000  9.610000 41.150000 ;
        RECT  9.410000 41.380000  9.610000 41.580000 ;
        RECT  9.410000 41.810000  9.610000 42.010000 ;
        RECT  9.410000 42.240000  9.610000 42.440000 ;
        RECT  9.410000 42.670000  9.610000 42.870000 ;
        RECT  9.410000 43.100000  9.610000 43.300000 ;
        RECT  9.410000 43.530000  9.610000 43.730000 ;
        RECT  9.410000 43.960000  9.610000 44.160000 ;
        RECT  9.810000 39.660000 10.010000 39.860000 ;
        RECT  9.810000 40.090000 10.010000 40.290000 ;
        RECT  9.810000 40.520000 10.010000 40.720000 ;
        RECT  9.810000 40.950000 10.010000 41.150000 ;
        RECT  9.810000 41.380000 10.010000 41.580000 ;
        RECT  9.810000 41.810000 10.010000 42.010000 ;
        RECT  9.810000 42.240000 10.010000 42.440000 ;
        RECT  9.810000 42.670000 10.010000 42.870000 ;
        RECT  9.810000 43.100000 10.010000 43.300000 ;
        RECT  9.810000 43.530000 10.010000 43.730000 ;
        RECT  9.810000 43.960000 10.010000 44.160000 ;
        RECT 10.210000 39.660000 10.410000 39.860000 ;
        RECT 10.210000 40.090000 10.410000 40.290000 ;
        RECT 10.210000 40.520000 10.410000 40.720000 ;
        RECT 10.210000 40.950000 10.410000 41.150000 ;
        RECT 10.210000 41.380000 10.410000 41.580000 ;
        RECT 10.210000 41.810000 10.410000 42.010000 ;
        RECT 10.210000 42.240000 10.410000 42.440000 ;
        RECT 10.210000 42.670000 10.410000 42.870000 ;
        RECT 10.210000 43.100000 10.410000 43.300000 ;
        RECT 10.210000 43.530000 10.410000 43.730000 ;
        RECT 10.210000 43.960000 10.410000 44.160000 ;
        RECT 10.610000 39.660000 10.810000 39.860000 ;
        RECT 10.610000 40.090000 10.810000 40.290000 ;
        RECT 10.610000 40.520000 10.810000 40.720000 ;
        RECT 10.610000 40.950000 10.810000 41.150000 ;
        RECT 10.610000 41.380000 10.810000 41.580000 ;
        RECT 10.610000 41.810000 10.810000 42.010000 ;
        RECT 10.610000 42.240000 10.810000 42.440000 ;
        RECT 10.610000 42.670000 10.810000 42.870000 ;
        RECT 10.610000 43.100000 10.810000 43.300000 ;
        RECT 10.610000 43.530000 10.810000 43.730000 ;
        RECT 10.610000 43.960000 10.810000 44.160000 ;
        RECT 11.010000 39.660000 11.210000 39.860000 ;
        RECT 11.010000 40.090000 11.210000 40.290000 ;
        RECT 11.010000 40.520000 11.210000 40.720000 ;
        RECT 11.010000 40.950000 11.210000 41.150000 ;
        RECT 11.010000 41.380000 11.210000 41.580000 ;
        RECT 11.010000 41.810000 11.210000 42.010000 ;
        RECT 11.010000 42.240000 11.210000 42.440000 ;
        RECT 11.010000 42.670000 11.210000 42.870000 ;
        RECT 11.010000 43.100000 11.210000 43.300000 ;
        RECT 11.010000 43.530000 11.210000 43.730000 ;
        RECT 11.010000 43.960000 11.210000 44.160000 ;
        RECT 11.410000 39.660000 11.610000 39.860000 ;
        RECT 11.410000 40.090000 11.610000 40.290000 ;
        RECT 11.410000 40.520000 11.610000 40.720000 ;
        RECT 11.410000 40.950000 11.610000 41.150000 ;
        RECT 11.410000 41.380000 11.610000 41.580000 ;
        RECT 11.410000 41.810000 11.610000 42.010000 ;
        RECT 11.410000 42.240000 11.610000 42.440000 ;
        RECT 11.410000 42.670000 11.610000 42.870000 ;
        RECT 11.410000 43.100000 11.610000 43.300000 ;
        RECT 11.410000 43.530000 11.610000 43.730000 ;
        RECT 11.410000 43.960000 11.610000 44.160000 ;
        RECT 11.810000 39.660000 12.010000 39.860000 ;
        RECT 11.810000 40.090000 12.010000 40.290000 ;
        RECT 11.810000 40.520000 12.010000 40.720000 ;
        RECT 11.810000 40.950000 12.010000 41.150000 ;
        RECT 11.810000 41.380000 12.010000 41.580000 ;
        RECT 11.810000 41.810000 12.010000 42.010000 ;
        RECT 11.810000 42.240000 12.010000 42.440000 ;
        RECT 11.810000 42.670000 12.010000 42.870000 ;
        RECT 11.810000 43.100000 12.010000 43.300000 ;
        RECT 11.810000 43.530000 12.010000 43.730000 ;
        RECT 11.810000 43.960000 12.010000 44.160000 ;
        RECT 12.210000 39.660000 12.410000 39.860000 ;
        RECT 12.210000 40.090000 12.410000 40.290000 ;
        RECT 12.210000 40.520000 12.410000 40.720000 ;
        RECT 12.210000 40.950000 12.410000 41.150000 ;
        RECT 12.210000 41.380000 12.410000 41.580000 ;
        RECT 12.210000 41.810000 12.410000 42.010000 ;
        RECT 12.210000 42.240000 12.410000 42.440000 ;
        RECT 12.210000 42.670000 12.410000 42.870000 ;
        RECT 12.210000 43.100000 12.410000 43.300000 ;
        RECT 12.210000 43.530000 12.410000 43.730000 ;
        RECT 12.210000 43.960000 12.410000 44.160000 ;
        RECT 12.610000 39.660000 12.810000 39.860000 ;
        RECT 12.610000 40.090000 12.810000 40.290000 ;
        RECT 12.610000 40.520000 12.810000 40.720000 ;
        RECT 12.610000 40.950000 12.810000 41.150000 ;
        RECT 12.610000 41.380000 12.810000 41.580000 ;
        RECT 12.610000 41.810000 12.810000 42.010000 ;
        RECT 12.610000 42.240000 12.810000 42.440000 ;
        RECT 12.610000 42.670000 12.810000 42.870000 ;
        RECT 12.610000 43.100000 12.810000 43.300000 ;
        RECT 12.610000 43.530000 12.810000 43.730000 ;
        RECT 12.610000 43.960000 12.810000 44.160000 ;
        RECT 13.010000 39.660000 13.210000 39.860000 ;
        RECT 13.010000 40.090000 13.210000 40.290000 ;
        RECT 13.010000 40.520000 13.210000 40.720000 ;
        RECT 13.010000 40.950000 13.210000 41.150000 ;
        RECT 13.010000 41.380000 13.210000 41.580000 ;
        RECT 13.010000 41.810000 13.210000 42.010000 ;
        RECT 13.010000 42.240000 13.210000 42.440000 ;
        RECT 13.010000 42.670000 13.210000 42.870000 ;
        RECT 13.010000 43.100000 13.210000 43.300000 ;
        RECT 13.010000 43.530000 13.210000 43.730000 ;
        RECT 13.010000 43.960000 13.210000 44.160000 ;
        RECT 13.410000 39.660000 13.610000 39.860000 ;
        RECT 13.410000 40.090000 13.610000 40.290000 ;
        RECT 13.410000 40.520000 13.610000 40.720000 ;
        RECT 13.410000 40.950000 13.610000 41.150000 ;
        RECT 13.410000 41.380000 13.610000 41.580000 ;
        RECT 13.410000 41.810000 13.610000 42.010000 ;
        RECT 13.410000 42.240000 13.610000 42.440000 ;
        RECT 13.410000 42.670000 13.610000 42.870000 ;
        RECT 13.410000 43.100000 13.610000 43.300000 ;
        RECT 13.410000 43.530000 13.610000 43.730000 ;
        RECT 13.410000 43.960000 13.610000 44.160000 ;
        RECT 13.810000 39.660000 14.010000 39.860000 ;
        RECT 13.810000 40.090000 14.010000 40.290000 ;
        RECT 13.810000 40.520000 14.010000 40.720000 ;
        RECT 13.810000 40.950000 14.010000 41.150000 ;
        RECT 13.810000 41.380000 14.010000 41.580000 ;
        RECT 13.810000 41.810000 14.010000 42.010000 ;
        RECT 13.810000 42.240000 14.010000 42.440000 ;
        RECT 13.810000 42.670000 14.010000 42.870000 ;
        RECT 13.810000 43.100000 14.010000 43.300000 ;
        RECT 13.810000 43.530000 14.010000 43.730000 ;
        RECT 13.810000 43.960000 14.010000 44.160000 ;
        RECT 14.210000 39.660000 14.410000 39.860000 ;
        RECT 14.210000 40.090000 14.410000 40.290000 ;
        RECT 14.210000 40.520000 14.410000 40.720000 ;
        RECT 14.210000 40.950000 14.410000 41.150000 ;
        RECT 14.210000 41.380000 14.410000 41.580000 ;
        RECT 14.210000 41.810000 14.410000 42.010000 ;
        RECT 14.210000 42.240000 14.410000 42.440000 ;
        RECT 14.210000 42.670000 14.410000 42.870000 ;
        RECT 14.210000 43.100000 14.410000 43.300000 ;
        RECT 14.210000 43.530000 14.410000 43.730000 ;
        RECT 14.210000 43.960000 14.410000 44.160000 ;
        RECT 14.610000 39.660000 14.810000 39.860000 ;
        RECT 14.610000 40.090000 14.810000 40.290000 ;
        RECT 14.610000 40.520000 14.810000 40.720000 ;
        RECT 14.610000 40.950000 14.810000 41.150000 ;
        RECT 14.610000 41.380000 14.810000 41.580000 ;
        RECT 14.610000 41.810000 14.810000 42.010000 ;
        RECT 14.610000 42.240000 14.810000 42.440000 ;
        RECT 14.610000 42.670000 14.810000 42.870000 ;
        RECT 14.610000 43.100000 14.810000 43.300000 ;
        RECT 14.610000 43.530000 14.810000 43.730000 ;
        RECT 14.610000 43.960000 14.810000 44.160000 ;
        RECT 15.010000 39.660000 15.210000 39.860000 ;
        RECT 15.010000 40.090000 15.210000 40.290000 ;
        RECT 15.010000 40.520000 15.210000 40.720000 ;
        RECT 15.010000 40.950000 15.210000 41.150000 ;
        RECT 15.010000 41.380000 15.210000 41.580000 ;
        RECT 15.010000 41.810000 15.210000 42.010000 ;
        RECT 15.010000 42.240000 15.210000 42.440000 ;
        RECT 15.010000 42.670000 15.210000 42.870000 ;
        RECT 15.010000 43.100000 15.210000 43.300000 ;
        RECT 15.010000 43.530000 15.210000 43.730000 ;
        RECT 15.010000 43.960000 15.210000 44.160000 ;
        RECT 15.410000 39.660000 15.610000 39.860000 ;
        RECT 15.410000 40.090000 15.610000 40.290000 ;
        RECT 15.410000 40.520000 15.610000 40.720000 ;
        RECT 15.410000 40.950000 15.610000 41.150000 ;
        RECT 15.410000 41.380000 15.610000 41.580000 ;
        RECT 15.410000 41.810000 15.610000 42.010000 ;
        RECT 15.410000 42.240000 15.610000 42.440000 ;
        RECT 15.410000 42.670000 15.610000 42.870000 ;
        RECT 15.410000 43.100000 15.610000 43.300000 ;
        RECT 15.410000 43.530000 15.610000 43.730000 ;
        RECT 15.410000 43.960000 15.610000 44.160000 ;
        RECT 15.810000 39.660000 16.010000 39.860000 ;
        RECT 15.810000 40.090000 16.010000 40.290000 ;
        RECT 15.810000 40.520000 16.010000 40.720000 ;
        RECT 15.810000 40.950000 16.010000 41.150000 ;
        RECT 15.810000 41.380000 16.010000 41.580000 ;
        RECT 15.810000 41.810000 16.010000 42.010000 ;
        RECT 15.810000 42.240000 16.010000 42.440000 ;
        RECT 15.810000 42.670000 16.010000 42.870000 ;
        RECT 15.810000 43.100000 16.010000 43.300000 ;
        RECT 15.810000 43.530000 16.010000 43.730000 ;
        RECT 15.810000 43.960000 16.010000 44.160000 ;
        RECT 16.210000 39.660000 16.410000 39.860000 ;
        RECT 16.210000 40.090000 16.410000 40.290000 ;
        RECT 16.210000 40.520000 16.410000 40.720000 ;
        RECT 16.210000 40.950000 16.410000 41.150000 ;
        RECT 16.210000 41.380000 16.410000 41.580000 ;
        RECT 16.210000 41.810000 16.410000 42.010000 ;
        RECT 16.210000 42.240000 16.410000 42.440000 ;
        RECT 16.210000 42.670000 16.410000 42.870000 ;
        RECT 16.210000 43.100000 16.410000 43.300000 ;
        RECT 16.210000 43.530000 16.410000 43.730000 ;
        RECT 16.210000 43.960000 16.410000 44.160000 ;
        RECT 16.610000 39.660000 16.810000 39.860000 ;
        RECT 16.610000 40.090000 16.810000 40.290000 ;
        RECT 16.610000 40.520000 16.810000 40.720000 ;
        RECT 16.610000 40.950000 16.810000 41.150000 ;
        RECT 16.610000 41.380000 16.810000 41.580000 ;
        RECT 16.610000 41.810000 16.810000 42.010000 ;
        RECT 16.610000 42.240000 16.810000 42.440000 ;
        RECT 16.610000 42.670000 16.810000 42.870000 ;
        RECT 16.610000 43.100000 16.810000 43.300000 ;
        RECT 16.610000 43.530000 16.810000 43.730000 ;
        RECT 16.610000 43.960000 16.810000 44.160000 ;
        RECT 17.010000 39.660000 17.210000 39.860000 ;
        RECT 17.010000 40.090000 17.210000 40.290000 ;
        RECT 17.010000 40.520000 17.210000 40.720000 ;
        RECT 17.010000 40.950000 17.210000 41.150000 ;
        RECT 17.010000 41.380000 17.210000 41.580000 ;
        RECT 17.010000 41.810000 17.210000 42.010000 ;
        RECT 17.010000 42.240000 17.210000 42.440000 ;
        RECT 17.010000 42.670000 17.210000 42.870000 ;
        RECT 17.010000 43.100000 17.210000 43.300000 ;
        RECT 17.010000 43.530000 17.210000 43.730000 ;
        RECT 17.010000 43.960000 17.210000 44.160000 ;
        RECT 17.410000 39.660000 17.610000 39.860000 ;
        RECT 17.410000 40.090000 17.610000 40.290000 ;
        RECT 17.410000 40.520000 17.610000 40.720000 ;
        RECT 17.410000 40.950000 17.610000 41.150000 ;
        RECT 17.410000 41.380000 17.610000 41.580000 ;
        RECT 17.410000 41.810000 17.610000 42.010000 ;
        RECT 17.410000 42.240000 17.610000 42.440000 ;
        RECT 17.410000 42.670000 17.610000 42.870000 ;
        RECT 17.410000 43.100000 17.610000 43.300000 ;
        RECT 17.410000 43.530000 17.610000 43.730000 ;
        RECT 17.410000 43.960000 17.610000 44.160000 ;
        RECT 17.810000 39.660000 18.010000 39.860000 ;
        RECT 17.810000 40.090000 18.010000 40.290000 ;
        RECT 17.810000 40.520000 18.010000 40.720000 ;
        RECT 17.810000 40.950000 18.010000 41.150000 ;
        RECT 17.810000 41.380000 18.010000 41.580000 ;
        RECT 17.810000 41.810000 18.010000 42.010000 ;
        RECT 17.810000 42.240000 18.010000 42.440000 ;
        RECT 17.810000 42.670000 18.010000 42.870000 ;
        RECT 17.810000 43.100000 18.010000 43.300000 ;
        RECT 17.810000 43.530000 18.010000 43.730000 ;
        RECT 17.810000 43.960000 18.010000 44.160000 ;
        RECT 18.210000 39.660000 18.410000 39.860000 ;
        RECT 18.210000 40.090000 18.410000 40.290000 ;
        RECT 18.210000 40.520000 18.410000 40.720000 ;
        RECT 18.210000 40.950000 18.410000 41.150000 ;
        RECT 18.210000 41.380000 18.410000 41.580000 ;
        RECT 18.210000 41.810000 18.410000 42.010000 ;
        RECT 18.210000 42.240000 18.410000 42.440000 ;
        RECT 18.210000 42.670000 18.410000 42.870000 ;
        RECT 18.210000 43.100000 18.410000 43.300000 ;
        RECT 18.210000 43.530000 18.410000 43.730000 ;
        RECT 18.210000 43.960000 18.410000 44.160000 ;
        RECT 18.610000 39.660000 18.810000 39.860000 ;
        RECT 18.610000 40.090000 18.810000 40.290000 ;
        RECT 18.610000 40.520000 18.810000 40.720000 ;
        RECT 18.610000 40.950000 18.810000 41.150000 ;
        RECT 18.610000 41.380000 18.810000 41.580000 ;
        RECT 18.610000 41.810000 18.810000 42.010000 ;
        RECT 18.610000 42.240000 18.810000 42.440000 ;
        RECT 18.610000 42.670000 18.810000 42.870000 ;
        RECT 18.610000 43.100000 18.810000 43.300000 ;
        RECT 18.610000 43.530000 18.810000 43.730000 ;
        RECT 18.610000 43.960000 18.810000 44.160000 ;
        RECT 19.010000 39.660000 19.210000 39.860000 ;
        RECT 19.010000 40.090000 19.210000 40.290000 ;
        RECT 19.010000 40.520000 19.210000 40.720000 ;
        RECT 19.010000 40.950000 19.210000 41.150000 ;
        RECT 19.010000 41.380000 19.210000 41.580000 ;
        RECT 19.010000 41.810000 19.210000 42.010000 ;
        RECT 19.010000 42.240000 19.210000 42.440000 ;
        RECT 19.010000 42.670000 19.210000 42.870000 ;
        RECT 19.010000 43.100000 19.210000 43.300000 ;
        RECT 19.010000 43.530000 19.210000 43.730000 ;
        RECT 19.010000 43.960000 19.210000 44.160000 ;
        RECT 19.410000 39.660000 19.610000 39.860000 ;
        RECT 19.410000 40.090000 19.610000 40.290000 ;
        RECT 19.410000 40.520000 19.610000 40.720000 ;
        RECT 19.410000 40.950000 19.610000 41.150000 ;
        RECT 19.410000 41.380000 19.610000 41.580000 ;
        RECT 19.410000 41.810000 19.610000 42.010000 ;
        RECT 19.410000 42.240000 19.610000 42.440000 ;
        RECT 19.410000 42.670000 19.610000 42.870000 ;
        RECT 19.410000 43.100000 19.610000 43.300000 ;
        RECT 19.410000 43.530000 19.610000 43.730000 ;
        RECT 19.410000 43.960000 19.610000 44.160000 ;
        RECT 19.810000 39.660000 20.010000 39.860000 ;
        RECT 19.810000 40.090000 20.010000 40.290000 ;
        RECT 19.810000 40.520000 20.010000 40.720000 ;
        RECT 19.810000 40.950000 20.010000 41.150000 ;
        RECT 19.810000 41.380000 20.010000 41.580000 ;
        RECT 19.810000 41.810000 20.010000 42.010000 ;
        RECT 19.810000 42.240000 20.010000 42.440000 ;
        RECT 19.810000 42.670000 20.010000 42.870000 ;
        RECT 19.810000 43.100000 20.010000 43.300000 ;
        RECT 19.810000 43.530000 20.010000 43.730000 ;
        RECT 19.810000 43.960000 20.010000 44.160000 ;
        RECT 20.210000 39.660000 20.410000 39.860000 ;
        RECT 20.210000 40.090000 20.410000 40.290000 ;
        RECT 20.210000 40.520000 20.410000 40.720000 ;
        RECT 20.210000 40.950000 20.410000 41.150000 ;
        RECT 20.210000 41.380000 20.410000 41.580000 ;
        RECT 20.210000 41.810000 20.410000 42.010000 ;
        RECT 20.210000 42.240000 20.410000 42.440000 ;
        RECT 20.210000 42.670000 20.410000 42.870000 ;
        RECT 20.210000 43.100000 20.410000 43.300000 ;
        RECT 20.210000 43.530000 20.410000 43.730000 ;
        RECT 20.210000 43.960000 20.410000 44.160000 ;
        RECT 20.610000 39.660000 20.810000 39.860000 ;
        RECT 20.610000 40.090000 20.810000 40.290000 ;
        RECT 20.610000 40.520000 20.810000 40.720000 ;
        RECT 20.610000 40.950000 20.810000 41.150000 ;
        RECT 20.610000 41.380000 20.810000 41.580000 ;
        RECT 20.610000 41.810000 20.810000 42.010000 ;
        RECT 20.610000 42.240000 20.810000 42.440000 ;
        RECT 20.610000 42.670000 20.810000 42.870000 ;
        RECT 20.610000 43.100000 20.810000 43.300000 ;
        RECT 20.610000 43.530000 20.810000 43.730000 ;
        RECT 20.610000 43.960000 20.810000 44.160000 ;
        RECT 21.010000 39.660000 21.210000 39.860000 ;
        RECT 21.010000 40.090000 21.210000 40.290000 ;
        RECT 21.010000 40.520000 21.210000 40.720000 ;
        RECT 21.010000 40.950000 21.210000 41.150000 ;
        RECT 21.010000 41.380000 21.210000 41.580000 ;
        RECT 21.010000 41.810000 21.210000 42.010000 ;
        RECT 21.010000 42.240000 21.210000 42.440000 ;
        RECT 21.010000 42.670000 21.210000 42.870000 ;
        RECT 21.010000 43.100000 21.210000 43.300000 ;
        RECT 21.010000 43.530000 21.210000 43.730000 ;
        RECT 21.010000 43.960000 21.210000 44.160000 ;
        RECT 21.410000 39.660000 21.610000 39.860000 ;
        RECT 21.410000 40.090000 21.610000 40.290000 ;
        RECT 21.410000 40.520000 21.610000 40.720000 ;
        RECT 21.410000 40.950000 21.610000 41.150000 ;
        RECT 21.410000 41.380000 21.610000 41.580000 ;
        RECT 21.410000 41.810000 21.610000 42.010000 ;
        RECT 21.410000 42.240000 21.610000 42.440000 ;
        RECT 21.410000 42.670000 21.610000 42.870000 ;
        RECT 21.410000 43.100000 21.610000 43.300000 ;
        RECT 21.410000 43.530000 21.610000 43.730000 ;
        RECT 21.410000 43.960000 21.610000 44.160000 ;
        RECT 21.810000 39.660000 22.010000 39.860000 ;
        RECT 21.810000 40.090000 22.010000 40.290000 ;
        RECT 21.810000 40.520000 22.010000 40.720000 ;
        RECT 21.810000 40.950000 22.010000 41.150000 ;
        RECT 21.810000 41.380000 22.010000 41.580000 ;
        RECT 21.810000 41.810000 22.010000 42.010000 ;
        RECT 21.810000 42.240000 22.010000 42.440000 ;
        RECT 21.810000 42.670000 22.010000 42.870000 ;
        RECT 21.810000 43.100000 22.010000 43.300000 ;
        RECT 21.810000 43.530000 22.010000 43.730000 ;
        RECT 21.810000 43.960000 22.010000 44.160000 ;
        RECT 22.210000 39.660000 22.410000 39.860000 ;
        RECT 22.210000 40.090000 22.410000 40.290000 ;
        RECT 22.210000 40.520000 22.410000 40.720000 ;
        RECT 22.210000 40.950000 22.410000 41.150000 ;
        RECT 22.210000 41.380000 22.410000 41.580000 ;
        RECT 22.210000 41.810000 22.410000 42.010000 ;
        RECT 22.210000 42.240000 22.410000 42.440000 ;
        RECT 22.210000 42.670000 22.410000 42.870000 ;
        RECT 22.210000 43.100000 22.410000 43.300000 ;
        RECT 22.210000 43.530000 22.410000 43.730000 ;
        RECT 22.210000 43.960000 22.410000 44.160000 ;
        RECT 22.610000 39.660000 22.810000 39.860000 ;
        RECT 22.610000 40.090000 22.810000 40.290000 ;
        RECT 22.610000 40.520000 22.810000 40.720000 ;
        RECT 22.610000 40.950000 22.810000 41.150000 ;
        RECT 22.610000 41.380000 22.810000 41.580000 ;
        RECT 22.610000 41.810000 22.810000 42.010000 ;
        RECT 22.610000 42.240000 22.810000 42.440000 ;
        RECT 22.610000 42.670000 22.810000 42.870000 ;
        RECT 22.610000 43.100000 22.810000 43.300000 ;
        RECT 22.610000 43.530000 22.810000 43.730000 ;
        RECT 22.610000 43.960000 22.810000 44.160000 ;
        RECT 23.010000 39.660000 23.210000 39.860000 ;
        RECT 23.010000 40.090000 23.210000 40.290000 ;
        RECT 23.010000 40.520000 23.210000 40.720000 ;
        RECT 23.010000 40.950000 23.210000 41.150000 ;
        RECT 23.010000 41.380000 23.210000 41.580000 ;
        RECT 23.010000 41.810000 23.210000 42.010000 ;
        RECT 23.010000 42.240000 23.210000 42.440000 ;
        RECT 23.010000 42.670000 23.210000 42.870000 ;
        RECT 23.010000 43.100000 23.210000 43.300000 ;
        RECT 23.010000 43.530000 23.210000 43.730000 ;
        RECT 23.010000 43.960000 23.210000 44.160000 ;
        RECT 23.410000 39.660000 23.610000 39.860000 ;
        RECT 23.410000 40.090000 23.610000 40.290000 ;
        RECT 23.410000 40.520000 23.610000 40.720000 ;
        RECT 23.410000 40.950000 23.610000 41.150000 ;
        RECT 23.410000 41.380000 23.610000 41.580000 ;
        RECT 23.410000 41.810000 23.610000 42.010000 ;
        RECT 23.410000 42.240000 23.610000 42.440000 ;
        RECT 23.410000 42.670000 23.610000 42.870000 ;
        RECT 23.410000 43.100000 23.610000 43.300000 ;
        RECT 23.410000 43.530000 23.610000 43.730000 ;
        RECT 23.410000 43.960000 23.610000 44.160000 ;
        RECT 23.810000 39.660000 24.010000 39.860000 ;
        RECT 23.810000 40.090000 24.010000 40.290000 ;
        RECT 23.810000 40.520000 24.010000 40.720000 ;
        RECT 23.810000 40.950000 24.010000 41.150000 ;
        RECT 23.810000 41.380000 24.010000 41.580000 ;
        RECT 23.810000 41.810000 24.010000 42.010000 ;
        RECT 23.810000 42.240000 24.010000 42.440000 ;
        RECT 23.810000 42.670000 24.010000 42.870000 ;
        RECT 23.810000 43.100000 24.010000 43.300000 ;
        RECT 23.810000 43.530000 24.010000 43.730000 ;
        RECT 23.810000 43.960000 24.010000 44.160000 ;
        RECT 24.210000 39.660000 24.410000 39.860000 ;
        RECT 24.210000 40.090000 24.410000 40.290000 ;
        RECT 24.210000 40.520000 24.410000 40.720000 ;
        RECT 24.210000 40.950000 24.410000 41.150000 ;
        RECT 24.210000 41.380000 24.410000 41.580000 ;
        RECT 24.210000 41.810000 24.410000 42.010000 ;
        RECT 24.210000 42.240000 24.410000 42.440000 ;
        RECT 24.210000 42.670000 24.410000 42.870000 ;
        RECT 24.210000 43.100000 24.410000 43.300000 ;
        RECT 24.210000 43.530000 24.410000 43.730000 ;
        RECT 24.210000 43.960000 24.410000 44.160000 ;
        RECT 50.845000 39.660000 51.045000 39.860000 ;
        RECT 50.845000 40.090000 51.045000 40.290000 ;
        RECT 50.845000 40.520000 51.045000 40.720000 ;
        RECT 50.845000 40.950000 51.045000 41.150000 ;
        RECT 50.845000 41.380000 51.045000 41.580000 ;
        RECT 50.845000 41.810000 51.045000 42.010000 ;
        RECT 50.845000 42.240000 51.045000 42.440000 ;
        RECT 50.845000 42.670000 51.045000 42.870000 ;
        RECT 50.845000 43.100000 51.045000 43.300000 ;
        RECT 50.845000 43.530000 51.045000 43.730000 ;
        RECT 50.845000 43.960000 51.045000 44.160000 ;
        RECT 51.255000 39.660000 51.455000 39.860000 ;
        RECT 51.255000 40.090000 51.455000 40.290000 ;
        RECT 51.255000 40.520000 51.455000 40.720000 ;
        RECT 51.255000 40.950000 51.455000 41.150000 ;
        RECT 51.255000 41.380000 51.455000 41.580000 ;
        RECT 51.255000 41.810000 51.455000 42.010000 ;
        RECT 51.255000 42.240000 51.455000 42.440000 ;
        RECT 51.255000 42.670000 51.455000 42.870000 ;
        RECT 51.255000 43.100000 51.455000 43.300000 ;
        RECT 51.255000 43.530000 51.455000 43.730000 ;
        RECT 51.255000 43.960000 51.455000 44.160000 ;
        RECT 51.665000 39.660000 51.865000 39.860000 ;
        RECT 51.665000 40.090000 51.865000 40.290000 ;
        RECT 51.665000 40.520000 51.865000 40.720000 ;
        RECT 51.665000 40.950000 51.865000 41.150000 ;
        RECT 51.665000 41.380000 51.865000 41.580000 ;
        RECT 51.665000 41.810000 51.865000 42.010000 ;
        RECT 51.665000 42.240000 51.865000 42.440000 ;
        RECT 51.665000 42.670000 51.865000 42.870000 ;
        RECT 51.665000 43.100000 51.865000 43.300000 ;
        RECT 51.665000 43.530000 51.865000 43.730000 ;
        RECT 51.665000 43.960000 51.865000 44.160000 ;
        RECT 52.075000 39.660000 52.275000 39.860000 ;
        RECT 52.075000 40.090000 52.275000 40.290000 ;
        RECT 52.075000 40.520000 52.275000 40.720000 ;
        RECT 52.075000 40.950000 52.275000 41.150000 ;
        RECT 52.075000 41.380000 52.275000 41.580000 ;
        RECT 52.075000 41.810000 52.275000 42.010000 ;
        RECT 52.075000 42.240000 52.275000 42.440000 ;
        RECT 52.075000 42.670000 52.275000 42.870000 ;
        RECT 52.075000 43.100000 52.275000 43.300000 ;
        RECT 52.075000 43.530000 52.275000 43.730000 ;
        RECT 52.075000 43.960000 52.275000 44.160000 ;
        RECT 52.485000 39.660000 52.685000 39.860000 ;
        RECT 52.485000 40.090000 52.685000 40.290000 ;
        RECT 52.485000 40.520000 52.685000 40.720000 ;
        RECT 52.485000 40.950000 52.685000 41.150000 ;
        RECT 52.485000 41.380000 52.685000 41.580000 ;
        RECT 52.485000 41.810000 52.685000 42.010000 ;
        RECT 52.485000 42.240000 52.685000 42.440000 ;
        RECT 52.485000 42.670000 52.685000 42.870000 ;
        RECT 52.485000 43.100000 52.685000 43.300000 ;
        RECT 52.485000 43.530000 52.685000 43.730000 ;
        RECT 52.485000 43.960000 52.685000 44.160000 ;
        RECT 52.895000 39.660000 53.095000 39.860000 ;
        RECT 52.895000 40.090000 53.095000 40.290000 ;
        RECT 52.895000 40.520000 53.095000 40.720000 ;
        RECT 52.895000 40.950000 53.095000 41.150000 ;
        RECT 52.895000 41.380000 53.095000 41.580000 ;
        RECT 52.895000 41.810000 53.095000 42.010000 ;
        RECT 52.895000 42.240000 53.095000 42.440000 ;
        RECT 52.895000 42.670000 53.095000 42.870000 ;
        RECT 52.895000 43.100000 53.095000 43.300000 ;
        RECT 52.895000 43.530000 53.095000 43.730000 ;
        RECT 52.895000 43.960000 53.095000 44.160000 ;
        RECT 53.305000 39.660000 53.505000 39.860000 ;
        RECT 53.305000 40.090000 53.505000 40.290000 ;
        RECT 53.305000 40.520000 53.505000 40.720000 ;
        RECT 53.305000 40.950000 53.505000 41.150000 ;
        RECT 53.305000 41.380000 53.505000 41.580000 ;
        RECT 53.305000 41.810000 53.505000 42.010000 ;
        RECT 53.305000 42.240000 53.505000 42.440000 ;
        RECT 53.305000 42.670000 53.505000 42.870000 ;
        RECT 53.305000 43.100000 53.505000 43.300000 ;
        RECT 53.305000 43.530000 53.505000 43.730000 ;
        RECT 53.305000 43.960000 53.505000 44.160000 ;
        RECT 53.715000 39.660000 53.915000 39.860000 ;
        RECT 53.715000 40.090000 53.915000 40.290000 ;
        RECT 53.715000 40.520000 53.915000 40.720000 ;
        RECT 53.715000 40.950000 53.915000 41.150000 ;
        RECT 53.715000 41.380000 53.915000 41.580000 ;
        RECT 53.715000 41.810000 53.915000 42.010000 ;
        RECT 53.715000 42.240000 53.915000 42.440000 ;
        RECT 53.715000 42.670000 53.915000 42.870000 ;
        RECT 53.715000 43.100000 53.915000 43.300000 ;
        RECT 53.715000 43.530000 53.915000 43.730000 ;
        RECT 53.715000 43.960000 53.915000 44.160000 ;
        RECT 54.125000 39.660000 54.325000 39.860000 ;
        RECT 54.125000 40.090000 54.325000 40.290000 ;
        RECT 54.125000 40.520000 54.325000 40.720000 ;
        RECT 54.125000 40.950000 54.325000 41.150000 ;
        RECT 54.125000 41.380000 54.325000 41.580000 ;
        RECT 54.125000 41.810000 54.325000 42.010000 ;
        RECT 54.125000 42.240000 54.325000 42.440000 ;
        RECT 54.125000 42.670000 54.325000 42.870000 ;
        RECT 54.125000 43.100000 54.325000 43.300000 ;
        RECT 54.125000 43.530000 54.325000 43.730000 ;
        RECT 54.125000 43.960000 54.325000 44.160000 ;
        RECT 54.535000 39.660000 54.735000 39.860000 ;
        RECT 54.535000 40.090000 54.735000 40.290000 ;
        RECT 54.535000 40.520000 54.735000 40.720000 ;
        RECT 54.535000 40.950000 54.735000 41.150000 ;
        RECT 54.535000 41.380000 54.735000 41.580000 ;
        RECT 54.535000 41.810000 54.735000 42.010000 ;
        RECT 54.535000 42.240000 54.735000 42.440000 ;
        RECT 54.535000 42.670000 54.735000 42.870000 ;
        RECT 54.535000 43.100000 54.735000 43.300000 ;
        RECT 54.535000 43.530000 54.735000 43.730000 ;
        RECT 54.535000 43.960000 54.735000 44.160000 ;
        RECT 54.945000 39.660000 55.145000 39.860000 ;
        RECT 54.945000 40.090000 55.145000 40.290000 ;
        RECT 54.945000 40.520000 55.145000 40.720000 ;
        RECT 54.945000 40.950000 55.145000 41.150000 ;
        RECT 54.945000 41.380000 55.145000 41.580000 ;
        RECT 54.945000 41.810000 55.145000 42.010000 ;
        RECT 54.945000 42.240000 55.145000 42.440000 ;
        RECT 54.945000 42.670000 55.145000 42.870000 ;
        RECT 54.945000 43.100000 55.145000 43.300000 ;
        RECT 54.945000 43.530000 55.145000 43.730000 ;
        RECT 54.945000 43.960000 55.145000 44.160000 ;
        RECT 55.355000 39.660000 55.555000 39.860000 ;
        RECT 55.355000 40.090000 55.555000 40.290000 ;
        RECT 55.355000 40.520000 55.555000 40.720000 ;
        RECT 55.355000 40.950000 55.555000 41.150000 ;
        RECT 55.355000 41.380000 55.555000 41.580000 ;
        RECT 55.355000 41.810000 55.555000 42.010000 ;
        RECT 55.355000 42.240000 55.555000 42.440000 ;
        RECT 55.355000 42.670000 55.555000 42.870000 ;
        RECT 55.355000 43.100000 55.555000 43.300000 ;
        RECT 55.355000 43.530000 55.555000 43.730000 ;
        RECT 55.355000 43.960000 55.555000 44.160000 ;
        RECT 55.765000 39.660000 55.965000 39.860000 ;
        RECT 55.765000 40.090000 55.965000 40.290000 ;
        RECT 55.765000 40.520000 55.965000 40.720000 ;
        RECT 55.765000 40.950000 55.965000 41.150000 ;
        RECT 55.765000 41.380000 55.965000 41.580000 ;
        RECT 55.765000 41.810000 55.965000 42.010000 ;
        RECT 55.765000 42.240000 55.965000 42.440000 ;
        RECT 55.765000 42.670000 55.965000 42.870000 ;
        RECT 55.765000 43.100000 55.965000 43.300000 ;
        RECT 55.765000 43.530000 55.965000 43.730000 ;
        RECT 55.765000 43.960000 55.965000 44.160000 ;
        RECT 56.175000 39.660000 56.375000 39.860000 ;
        RECT 56.175000 40.090000 56.375000 40.290000 ;
        RECT 56.175000 40.520000 56.375000 40.720000 ;
        RECT 56.175000 40.950000 56.375000 41.150000 ;
        RECT 56.175000 41.380000 56.375000 41.580000 ;
        RECT 56.175000 41.810000 56.375000 42.010000 ;
        RECT 56.175000 42.240000 56.375000 42.440000 ;
        RECT 56.175000 42.670000 56.375000 42.870000 ;
        RECT 56.175000 43.100000 56.375000 43.300000 ;
        RECT 56.175000 43.530000 56.375000 43.730000 ;
        RECT 56.175000 43.960000 56.375000 44.160000 ;
        RECT 56.585000 39.660000 56.785000 39.860000 ;
        RECT 56.585000 40.090000 56.785000 40.290000 ;
        RECT 56.585000 40.520000 56.785000 40.720000 ;
        RECT 56.585000 40.950000 56.785000 41.150000 ;
        RECT 56.585000 41.380000 56.785000 41.580000 ;
        RECT 56.585000 41.810000 56.785000 42.010000 ;
        RECT 56.585000 42.240000 56.785000 42.440000 ;
        RECT 56.585000 42.670000 56.785000 42.870000 ;
        RECT 56.585000 43.100000 56.785000 43.300000 ;
        RECT 56.585000 43.530000 56.785000 43.730000 ;
        RECT 56.585000 43.960000 56.785000 44.160000 ;
        RECT 56.995000 39.660000 57.195000 39.860000 ;
        RECT 56.995000 40.090000 57.195000 40.290000 ;
        RECT 56.995000 40.520000 57.195000 40.720000 ;
        RECT 56.995000 40.950000 57.195000 41.150000 ;
        RECT 56.995000 41.380000 57.195000 41.580000 ;
        RECT 56.995000 41.810000 57.195000 42.010000 ;
        RECT 56.995000 42.240000 57.195000 42.440000 ;
        RECT 56.995000 42.670000 57.195000 42.870000 ;
        RECT 56.995000 43.100000 57.195000 43.300000 ;
        RECT 56.995000 43.530000 57.195000 43.730000 ;
        RECT 56.995000 43.960000 57.195000 44.160000 ;
        RECT 57.400000 39.660000 57.600000 39.860000 ;
        RECT 57.400000 40.090000 57.600000 40.290000 ;
        RECT 57.400000 40.520000 57.600000 40.720000 ;
        RECT 57.400000 40.950000 57.600000 41.150000 ;
        RECT 57.400000 41.380000 57.600000 41.580000 ;
        RECT 57.400000 41.810000 57.600000 42.010000 ;
        RECT 57.400000 42.240000 57.600000 42.440000 ;
        RECT 57.400000 42.670000 57.600000 42.870000 ;
        RECT 57.400000 43.100000 57.600000 43.300000 ;
        RECT 57.400000 43.530000 57.600000 43.730000 ;
        RECT 57.400000 43.960000 57.600000 44.160000 ;
        RECT 57.805000 39.660000 58.005000 39.860000 ;
        RECT 57.805000 40.090000 58.005000 40.290000 ;
        RECT 57.805000 40.520000 58.005000 40.720000 ;
        RECT 57.805000 40.950000 58.005000 41.150000 ;
        RECT 57.805000 41.380000 58.005000 41.580000 ;
        RECT 57.805000 41.810000 58.005000 42.010000 ;
        RECT 57.805000 42.240000 58.005000 42.440000 ;
        RECT 57.805000 42.670000 58.005000 42.870000 ;
        RECT 57.805000 43.100000 58.005000 43.300000 ;
        RECT 57.805000 43.530000 58.005000 43.730000 ;
        RECT 57.805000 43.960000 58.005000 44.160000 ;
        RECT 58.210000 39.660000 58.410000 39.860000 ;
        RECT 58.210000 40.090000 58.410000 40.290000 ;
        RECT 58.210000 40.520000 58.410000 40.720000 ;
        RECT 58.210000 40.950000 58.410000 41.150000 ;
        RECT 58.210000 41.380000 58.410000 41.580000 ;
        RECT 58.210000 41.810000 58.410000 42.010000 ;
        RECT 58.210000 42.240000 58.410000 42.440000 ;
        RECT 58.210000 42.670000 58.410000 42.870000 ;
        RECT 58.210000 43.100000 58.410000 43.300000 ;
        RECT 58.210000 43.530000 58.410000 43.730000 ;
        RECT 58.210000 43.960000 58.410000 44.160000 ;
        RECT 58.615000 39.660000 58.815000 39.860000 ;
        RECT 58.615000 40.090000 58.815000 40.290000 ;
        RECT 58.615000 40.520000 58.815000 40.720000 ;
        RECT 58.615000 40.950000 58.815000 41.150000 ;
        RECT 58.615000 41.380000 58.815000 41.580000 ;
        RECT 58.615000 41.810000 58.815000 42.010000 ;
        RECT 58.615000 42.240000 58.815000 42.440000 ;
        RECT 58.615000 42.670000 58.815000 42.870000 ;
        RECT 58.615000 43.100000 58.815000 43.300000 ;
        RECT 58.615000 43.530000 58.815000 43.730000 ;
        RECT 58.615000 43.960000 58.815000 44.160000 ;
        RECT 59.020000 39.660000 59.220000 39.860000 ;
        RECT 59.020000 40.090000 59.220000 40.290000 ;
        RECT 59.020000 40.520000 59.220000 40.720000 ;
        RECT 59.020000 40.950000 59.220000 41.150000 ;
        RECT 59.020000 41.380000 59.220000 41.580000 ;
        RECT 59.020000 41.810000 59.220000 42.010000 ;
        RECT 59.020000 42.240000 59.220000 42.440000 ;
        RECT 59.020000 42.670000 59.220000 42.870000 ;
        RECT 59.020000 43.100000 59.220000 43.300000 ;
        RECT 59.020000 43.530000 59.220000 43.730000 ;
        RECT 59.020000 43.960000 59.220000 44.160000 ;
        RECT 59.425000 39.660000 59.625000 39.860000 ;
        RECT 59.425000 40.090000 59.625000 40.290000 ;
        RECT 59.425000 40.520000 59.625000 40.720000 ;
        RECT 59.425000 40.950000 59.625000 41.150000 ;
        RECT 59.425000 41.380000 59.625000 41.580000 ;
        RECT 59.425000 41.810000 59.625000 42.010000 ;
        RECT 59.425000 42.240000 59.625000 42.440000 ;
        RECT 59.425000 42.670000 59.625000 42.870000 ;
        RECT 59.425000 43.100000 59.625000 43.300000 ;
        RECT 59.425000 43.530000 59.625000 43.730000 ;
        RECT 59.425000 43.960000 59.625000 44.160000 ;
        RECT 59.830000 39.660000 60.030000 39.860000 ;
        RECT 59.830000 40.090000 60.030000 40.290000 ;
        RECT 59.830000 40.520000 60.030000 40.720000 ;
        RECT 59.830000 40.950000 60.030000 41.150000 ;
        RECT 59.830000 41.380000 60.030000 41.580000 ;
        RECT 59.830000 41.810000 60.030000 42.010000 ;
        RECT 59.830000 42.240000 60.030000 42.440000 ;
        RECT 59.830000 42.670000 60.030000 42.870000 ;
        RECT 59.830000 43.100000 60.030000 43.300000 ;
        RECT 59.830000 43.530000 60.030000 43.730000 ;
        RECT 59.830000 43.960000 60.030000 44.160000 ;
        RECT 60.235000 39.660000 60.435000 39.860000 ;
        RECT 60.235000 40.090000 60.435000 40.290000 ;
        RECT 60.235000 40.520000 60.435000 40.720000 ;
        RECT 60.235000 40.950000 60.435000 41.150000 ;
        RECT 60.235000 41.380000 60.435000 41.580000 ;
        RECT 60.235000 41.810000 60.435000 42.010000 ;
        RECT 60.235000 42.240000 60.435000 42.440000 ;
        RECT 60.235000 42.670000 60.435000 42.870000 ;
        RECT 60.235000 43.100000 60.435000 43.300000 ;
        RECT 60.235000 43.530000 60.435000 43.730000 ;
        RECT 60.235000 43.960000 60.435000 44.160000 ;
        RECT 60.640000 39.660000 60.840000 39.860000 ;
        RECT 60.640000 40.090000 60.840000 40.290000 ;
        RECT 60.640000 40.520000 60.840000 40.720000 ;
        RECT 60.640000 40.950000 60.840000 41.150000 ;
        RECT 60.640000 41.380000 60.840000 41.580000 ;
        RECT 60.640000 41.810000 60.840000 42.010000 ;
        RECT 60.640000 42.240000 60.840000 42.440000 ;
        RECT 60.640000 42.670000 60.840000 42.870000 ;
        RECT 60.640000 43.100000 60.840000 43.300000 ;
        RECT 60.640000 43.530000 60.840000 43.730000 ;
        RECT 60.640000 43.960000 60.840000 44.160000 ;
        RECT 61.045000 39.660000 61.245000 39.860000 ;
        RECT 61.045000 40.090000 61.245000 40.290000 ;
        RECT 61.045000 40.520000 61.245000 40.720000 ;
        RECT 61.045000 40.950000 61.245000 41.150000 ;
        RECT 61.045000 41.380000 61.245000 41.580000 ;
        RECT 61.045000 41.810000 61.245000 42.010000 ;
        RECT 61.045000 42.240000 61.245000 42.440000 ;
        RECT 61.045000 42.670000 61.245000 42.870000 ;
        RECT 61.045000 43.100000 61.245000 43.300000 ;
        RECT 61.045000 43.530000 61.245000 43.730000 ;
        RECT 61.045000 43.960000 61.245000 44.160000 ;
        RECT 61.450000 39.660000 61.650000 39.860000 ;
        RECT 61.450000 40.090000 61.650000 40.290000 ;
        RECT 61.450000 40.520000 61.650000 40.720000 ;
        RECT 61.450000 40.950000 61.650000 41.150000 ;
        RECT 61.450000 41.380000 61.650000 41.580000 ;
        RECT 61.450000 41.810000 61.650000 42.010000 ;
        RECT 61.450000 42.240000 61.650000 42.440000 ;
        RECT 61.450000 42.670000 61.650000 42.870000 ;
        RECT 61.450000 43.100000 61.650000 43.300000 ;
        RECT 61.450000 43.530000 61.650000 43.730000 ;
        RECT 61.450000 43.960000 61.650000 44.160000 ;
        RECT 61.855000 39.660000 62.055000 39.860000 ;
        RECT 61.855000 40.090000 62.055000 40.290000 ;
        RECT 61.855000 40.520000 62.055000 40.720000 ;
        RECT 61.855000 40.950000 62.055000 41.150000 ;
        RECT 61.855000 41.380000 62.055000 41.580000 ;
        RECT 61.855000 41.810000 62.055000 42.010000 ;
        RECT 61.855000 42.240000 62.055000 42.440000 ;
        RECT 61.855000 42.670000 62.055000 42.870000 ;
        RECT 61.855000 43.100000 62.055000 43.300000 ;
        RECT 61.855000 43.530000 62.055000 43.730000 ;
        RECT 61.855000 43.960000 62.055000 44.160000 ;
        RECT 62.260000 39.660000 62.460000 39.860000 ;
        RECT 62.260000 40.090000 62.460000 40.290000 ;
        RECT 62.260000 40.520000 62.460000 40.720000 ;
        RECT 62.260000 40.950000 62.460000 41.150000 ;
        RECT 62.260000 41.380000 62.460000 41.580000 ;
        RECT 62.260000 41.810000 62.460000 42.010000 ;
        RECT 62.260000 42.240000 62.460000 42.440000 ;
        RECT 62.260000 42.670000 62.460000 42.870000 ;
        RECT 62.260000 43.100000 62.460000 43.300000 ;
        RECT 62.260000 43.530000 62.460000 43.730000 ;
        RECT 62.260000 43.960000 62.460000 44.160000 ;
        RECT 62.665000 39.660000 62.865000 39.860000 ;
        RECT 62.665000 40.090000 62.865000 40.290000 ;
        RECT 62.665000 40.520000 62.865000 40.720000 ;
        RECT 62.665000 40.950000 62.865000 41.150000 ;
        RECT 62.665000 41.380000 62.865000 41.580000 ;
        RECT 62.665000 41.810000 62.865000 42.010000 ;
        RECT 62.665000 42.240000 62.865000 42.440000 ;
        RECT 62.665000 42.670000 62.865000 42.870000 ;
        RECT 62.665000 43.100000 62.865000 43.300000 ;
        RECT 62.665000 43.530000 62.865000 43.730000 ;
        RECT 62.665000 43.960000 62.865000 44.160000 ;
        RECT 63.070000 39.660000 63.270000 39.860000 ;
        RECT 63.070000 40.090000 63.270000 40.290000 ;
        RECT 63.070000 40.520000 63.270000 40.720000 ;
        RECT 63.070000 40.950000 63.270000 41.150000 ;
        RECT 63.070000 41.380000 63.270000 41.580000 ;
        RECT 63.070000 41.810000 63.270000 42.010000 ;
        RECT 63.070000 42.240000 63.270000 42.440000 ;
        RECT 63.070000 42.670000 63.270000 42.870000 ;
        RECT 63.070000 43.100000 63.270000 43.300000 ;
        RECT 63.070000 43.530000 63.270000 43.730000 ;
        RECT 63.070000 43.960000 63.270000 44.160000 ;
        RECT 63.475000 39.660000 63.675000 39.860000 ;
        RECT 63.475000 40.090000 63.675000 40.290000 ;
        RECT 63.475000 40.520000 63.675000 40.720000 ;
        RECT 63.475000 40.950000 63.675000 41.150000 ;
        RECT 63.475000 41.380000 63.675000 41.580000 ;
        RECT 63.475000 41.810000 63.675000 42.010000 ;
        RECT 63.475000 42.240000 63.675000 42.440000 ;
        RECT 63.475000 42.670000 63.675000 42.870000 ;
        RECT 63.475000 43.100000 63.675000 43.300000 ;
        RECT 63.475000 43.530000 63.675000 43.730000 ;
        RECT 63.475000 43.960000 63.675000 44.160000 ;
        RECT 63.880000 39.660000 64.080000 39.860000 ;
        RECT 63.880000 40.090000 64.080000 40.290000 ;
        RECT 63.880000 40.520000 64.080000 40.720000 ;
        RECT 63.880000 40.950000 64.080000 41.150000 ;
        RECT 63.880000 41.380000 64.080000 41.580000 ;
        RECT 63.880000 41.810000 64.080000 42.010000 ;
        RECT 63.880000 42.240000 64.080000 42.440000 ;
        RECT 63.880000 42.670000 64.080000 42.870000 ;
        RECT 63.880000 43.100000 64.080000 43.300000 ;
        RECT 63.880000 43.530000 64.080000 43.730000 ;
        RECT 63.880000 43.960000 64.080000 44.160000 ;
        RECT 64.285000 39.660000 64.485000 39.860000 ;
        RECT 64.285000 40.090000 64.485000 40.290000 ;
        RECT 64.285000 40.520000 64.485000 40.720000 ;
        RECT 64.285000 40.950000 64.485000 41.150000 ;
        RECT 64.285000 41.380000 64.485000 41.580000 ;
        RECT 64.285000 41.810000 64.485000 42.010000 ;
        RECT 64.285000 42.240000 64.485000 42.440000 ;
        RECT 64.285000 42.670000 64.485000 42.870000 ;
        RECT 64.285000 43.100000 64.485000 43.300000 ;
        RECT 64.285000 43.530000 64.485000 43.730000 ;
        RECT 64.285000 43.960000 64.485000 44.160000 ;
        RECT 64.690000 39.660000 64.890000 39.860000 ;
        RECT 64.690000 40.090000 64.890000 40.290000 ;
        RECT 64.690000 40.520000 64.890000 40.720000 ;
        RECT 64.690000 40.950000 64.890000 41.150000 ;
        RECT 64.690000 41.380000 64.890000 41.580000 ;
        RECT 64.690000 41.810000 64.890000 42.010000 ;
        RECT 64.690000 42.240000 64.890000 42.440000 ;
        RECT 64.690000 42.670000 64.890000 42.870000 ;
        RECT 64.690000 43.100000 64.890000 43.300000 ;
        RECT 64.690000 43.530000 64.890000 43.730000 ;
        RECT 64.690000 43.960000 64.890000 44.160000 ;
        RECT 65.095000 39.660000 65.295000 39.860000 ;
        RECT 65.095000 40.090000 65.295000 40.290000 ;
        RECT 65.095000 40.520000 65.295000 40.720000 ;
        RECT 65.095000 40.950000 65.295000 41.150000 ;
        RECT 65.095000 41.380000 65.295000 41.580000 ;
        RECT 65.095000 41.810000 65.295000 42.010000 ;
        RECT 65.095000 42.240000 65.295000 42.440000 ;
        RECT 65.095000 42.670000 65.295000 42.870000 ;
        RECT 65.095000 43.100000 65.295000 43.300000 ;
        RECT 65.095000 43.530000 65.295000 43.730000 ;
        RECT 65.095000 43.960000 65.295000 44.160000 ;
        RECT 65.500000 39.660000 65.700000 39.860000 ;
        RECT 65.500000 40.090000 65.700000 40.290000 ;
        RECT 65.500000 40.520000 65.700000 40.720000 ;
        RECT 65.500000 40.950000 65.700000 41.150000 ;
        RECT 65.500000 41.380000 65.700000 41.580000 ;
        RECT 65.500000 41.810000 65.700000 42.010000 ;
        RECT 65.500000 42.240000 65.700000 42.440000 ;
        RECT 65.500000 42.670000 65.700000 42.870000 ;
        RECT 65.500000 43.100000 65.700000 43.300000 ;
        RECT 65.500000 43.530000 65.700000 43.730000 ;
        RECT 65.500000 43.960000 65.700000 44.160000 ;
        RECT 65.905000 39.660000 66.105000 39.860000 ;
        RECT 65.905000 40.090000 66.105000 40.290000 ;
        RECT 65.905000 40.520000 66.105000 40.720000 ;
        RECT 65.905000 40.950000 66.105000 41.150000 ;
        RECT 65.905000 41.380000 66.105000 41.580000 ;
        RECT 65.905000 41.810000 66.105000 42.010000 ;
        RECT 65.905000 42.240000 66.105000 42.440000 ;
        RECT 65.905000 42.670000 66.105000 42.870000 ;
        RECT 65.905000 43.100000 66.105000 43.300000 ;
        RECT 65.905000 43.530000 66.105000 43.730000 ;
        RECT 65.905000 43.960000 66.105000 44.160000 ;
        RECT 66.310000 39.660000 66.510000 39.860000 ;
        RECT 66.310000 40.090000 66.510000 40.290000 ;
        RECT 66.310000 40.520000 66.510000 40.720000 ;
        RECT 66.310000 40.950000 66.510000 41.150000 ;
        RECT 66.310000 41.380000 66.510000 41.580000 ;
        RECT 66.310000 41.810000 66.510000 42.010000 ;
        RECT 66.310000 42.240000 66.510000 42.440000 ;
        RECT 66.310000 42.670000 66.510000 42.870000 ;
        RECT 66.310000 43.100000 66.510000 43.300000 ;
        RECT 66.310000 43.530000 66.510000 43.730000 ;
        RECT 66.310000 43.960000 66.510000 44.160000 ;
        RECT 66.715000 39.660000 66.915000 39.860000 ;
        RECT 66.715000 40.090000 66.915000 40.290000 ;
        RECT 66.715000 40.520000 66.915000 40.720000 ;
        RECT 66.715000 40.950000 66.915000 41.150000 ;
        RECT 66.715000 41.380000 66.915000 41.580000 ;
        RECT 66.715000 41.810000 66.915000 42.010000 ;
        RECT 66.715000 42.240000 66.915000 42.440000 ;
        RECT 66.715000 42.670000 66.915000 42.870000 ;
        RECT 66.715000 43.100000 66.915000 43.300000 ;
        RECT 66.715000 43.530000 66.915000 43.730000 ;
        RECT 66.715000 43.960000 66.915000 44.160000 ;
        RECT 67.120000 39.660000 67.320000 39.860000 ;
        RECT 67.120000 40.090000 67.320000 40.290000 ;
        RECT 67.120000 40.520000 67.320000 40.720000 ;
        RECT 67.120000 40.950000 67.320000 41.150000 ;
        RECT 67.120000 41.380000 67.320000 41.580000 ;
        RECT 67.120000 41.810000 67.320000 42.010000 ;
        RECT 67.120000 42.240000 67.320000 42.440000 ;
        RECT 67.120000 42.670000 67.320000 42.870000 ;
        RECT 67.120000 43.100000 67.320000 43.300000 ;
        RECT 67.120000 43.530000 67.320000 43.730000 ;
        RECT 67.120000 43.960000 67.320000 44.160000 ;
        RECT 67.525000 39.660000 67.725000 39.860000 ;
        RECT 67.525000 40.090000 67.725000 40.290000 ;
        RECT 67.525000 40.520000 67.725000 40.720000 ;
        RECT 67.525000 40.950000 67.725000 41.150000 ;
        RECT 67.525000 41.380000 67.725000 41.580000 ;
        RECT 67.525000 41.810000 67.725000 42.010000 ;
        RECT 67.525000 42.240000 67.725000 42.440000 ;
        RECT 67.525000 42.670000 67.725000 42.870000 ;
        RECT 67.525000 43.100000 67.725000 43.300000 ;
        RECT 67.525000 43.530000 67.725000 43.730000 ;
        RECT 67.525000 43.960000 67.725000 44.160000 ;
        RECT 67.930000 39.660000 68.130000 39.860000 ;
        RECT 67.930000 40.090000 68.130000 40.290000 ;
        RECT 67.930000 40.520000 68.130000 40.720000 ;
        RECT 67.930000 40.950000 68.130000 41.150000 ;
        RECT 67.930000 41.380000 68.130000 41.580000 ;
        RECT 67.930000 41.810000 68.130000 42.010000 ;
        RECT 67.930000 42.240000 68.130000 42.440000 ;
        RECT 67.930000 42.670000 68.130000 42.870000 ;
        RECT 67.930000 43.100000 68.130000 43.300000 ;
        RECT 67.930000 43.530000 68.130000 43.730000 ;
        RECT 67.930000 43.960000 68.130000 44.160000 ;
        RECT 68.335000 39.660000 68.535000 39.860000 ;
        RECT 68.335000 40.090000 68.535000 40.290000 ;
        RECT 68.335000 40.520000 68.535000 40.720000 ;
        RECT 68.335000 40.950000 68.535000 41.150000 ;
        RECT 68.335000 41.380000 68.535000 41.580000 ;
        RECT 68.335000 41.810000 68.535000 42.010000 ;
        RECT 68.335000 42.240000 68.535000 42.440000 ;
        RECT 68.335000 42.670000 68.535000 42.870000 ;
        RECT 68.335000 43.100000 68.535000 43.300000 ;
        RECT 68.335000 43.530000 68.535000 43.730000 ;
        RECT 68.335000 43.960000 68.535000 44.160000 ;
        RECT 68.740000 39.660000 68.940000 39.860000 ;
        RECT 68.740000 40.090000 68.940000 40.290000 ;
        RECT 68.740000 40.520000 68.940000 40.720000 ;
        RECT 68.740000 40.950000 68.940000 41.150000 ;
        RECT 68.740000 41.380000 68.940000 41.580000 ;
        RECT 68.740000 41.810000 68.940000 42.010000 ;
        RECT 68.740000 42.240000 68.940000 42.440000 ;
        RECT 68.740000 42.670000 68.940000 42.870000 ;
        RECT 68.740000 43.100000 68.940000 43.300000 ;
        RECT 68.740000 43.530000 68.940000 43.730000 ;
        RECT 68.740000 43.960000 68.940000 44.160000 ;
        RECT 69.145000 39.660000 69.345000 39.860000 ;
        RECT 69.145000 40.090000 69.345000 40.290000 ;
        RECT 69.145000 40.520000 69.345000 40.720000 ;
        RECT 69.145000 40.950000 69.345000 41.150000 ;
        RECT 69.145000 41.380000 69.345000 41.580000 ;
        RECT 69.145000 41.810000 69.345000 42.010000 ;
        RECT 69.145000 42.240000 69.345000 42.440000 ;
        RECT 69.145000 42.670000 69.345000 42.870000 ;
        RECT 69.145000 43.100000 69.345000 43.300000 ;
        RECT 69.145000 43.530000 69.345000 43.730000 ;
        RECT 69.145000 43.960000 69.345000 44.160000 ;
        RECT 69.550000 39.660000 69.750000 39.860000 ;
        RECT 69.550000 40.090000 69.750000 40.290000 ;
        RECT 69.550000 40.520000 69.750000 40.720000 ;
        RECT 69.550000 40.950000 69.750000 41.150000 ;
        RECT 69.550000 41.380000 69.750000 41.580000 ;
        RECT 69.550000 41.810000 69.750000 42.010000 ;
        RECT 69.550000 42.240000 69.750000 42.440000 ;
        RECT 69.550000 42.670000 69.750000 42.870000 ;
        RECT 69.550000 43.100000 69.750000 43.300000 ;
        RECT 69.550000 43.530000 69.750000 43.730000 ;
        RECT 69.550000 43.960000 69.750000 44.160000 ;
        RECT 69.955000 39.660000 70.155000 39.860000 ;
        RECT 69.955000 40.090000 70.155000 40.290000 ;
        RECT 69.955000 40.520000 70.155000 40.720000 ;
        RECT 69.955000 40.950000 70.155000 41.150000 ;
        RECT 69.955000 41.380000 70.155000 41.580000 ;
        RECT 69.955000 41.810000 70.155000 42.010000 ;
        RECT 69.955000 42.240000 70.155000 42.440000 ;
        RECT 69.955000 42.670000 70.155000 42.870000 ;
        RECT 69.955000 43.100000 70.155000 43.300000 ;
        RECT 69.955000 43.530000 70.155000 43.730000 ;
        RECT 69.955000 43.960000 70.155000 44.160000 ;
        RECT 70.360000 39.660000 70.560000 39.860000 ;
        RECT 70.360000 40.090000 70.560000 40.290000 ;
        RECT 70.360000 40.520000 70.560000 40.720000 ;
        RECT 70.360000 40.950000 70.560000 41.150000 ;
        RECT 70.360000 41.380000 70.560000 41.580000 ;
        RECT 70.360000 41.810000 70.560000 42.010000 ;
        RECT 70.360000 42.240000 70.560000 42.440000 ;
        RECT 70.360000 42.670000 70.560000 42.870000 ;
        RECT 70.360000 43.100000 70.560000 43.300000 ;
        RECT 70.360000 43.530000 70.560000 43.730000 ;
        RECT 70.360000 43.960000 70.560000 44.160000 ;
        RECT 70.765000 39.660000 70.965000 39.860000 ;
        RECT 70.765000 40.090000 70.965000 40.290000 ;
        RECT 70.765000 40.520000 70.965000 40.720000 ;
        RECT 70.765000 40.950000 70.965000 41.150000 ;
        RECT 70.765000 41.380000 70.965000 41.580000 ;
        RECT 70.765000 41.810000 70.965000 42.010000 ;
        RECT 70.765000 42.240000 70.965000 42.440000 ;
        RECT 70.765000 42.670000 70.965000 42.870000 ;
        RECT 70.765000 43.100000 70.965000 43.300000 ;
        RECT 70.765000 43.530000 70.965000 43.730000 ;
        RECT 70.765000 43.960000 70.965000 44.160000 ;
        RECT 71.170000 39.660000 71.370000 39.860000 ;
        RECT 71.170000 40.090000 71.370000 40.290000 ;
        RECT 71.170000 40.520000 71.370000 40.720000 ;
        RECT 71.170000 40.950000 71.370000 41.150000 ;
        RECT 71.170000 41.380000 71.370000 41.580000 ;
        RECT 71.170000 41.810000 71.370000 42.010000 ;
        RECT 71.170000 42.240000 71.370000 42.440000 ;
        RECT 71.170000 42.670000 71.370000 42.870000 ;
        RECT 71.170000 43.100000 71.370000 43.300000 ;
        RECT 71.170000 43.530000 71.370000 43.730000 ;
        RECT 71.170000 43.960000 71.370000 44.160000 ;
        RECT 71.575000 39.660000 71.775000 39.860000 ;
        RECT 71.575000 40.090000 71.775000 40.290000 ;
        RECT 71.575000 40.520000 71.775000 40.720000 ;
        RECT 71.575000 40.950000 71.775000 41.150000 ;
        RECT 71.575000 41.380000 71.775000 41.580000 ;
        RECT 71.575000 41.810000 71.775000 42.010000 ;
        RECT 71.575000 42.240000 71.775000 42.440000 ;
        RECT 71.575000 42.670000 71.775000 42.870000 ;
        RECT 71.575000 43.100000 71.775000 43.300000 ;
        RECT 71.575000 43.530000 71.775000 43.730000 ;
        RECT 71.575000 43.960000 71.775000 44.160000 ;
        RECT 71.980000 39.660000 72.180000 39.860000 ;
        RECT 71.980000 40.090000 72.180000 40.290000 ;
        RECT 71.980000 40.520000 72.180000 40.720000 ;
        RECT 71.980000 40.950000 72.180000 41.150000 ;
        RECT 71.980000 41.380000 72.180000 41.580000 ;
        RECT 71.980000 41.810000 72.180000 42.010000 ;
        RECT 71.980000 42.240000 72.180000 42.440000 ;
        RECT 71.980000 42.670000 72.180000 42.870000 ;
        RECT 71.980000 43.100000 72.180000 43.300000 ;
        RECT 71.980000 43.530000 72.180000 43.730000 ;
        RECT 71.980000 43.960000 72.180000 44.160000 ;
        RECT 72.385000 39.660000 72.585000 39.860000 ;
        RECT 72.385000 40.090000 72.585000 40.290000 ;
        RECT 72.385000 40.520000 72.585000 40.720000 ;
        RECT 72.385000 40.950000 72.585000 41.150000 ;
        RECT 72.385000 41.380000 72.585000 41.580000 ;
        RECT 72.385000 41.810000 72.585000 42.010000 ;
        RECT 72.385000 42.240000 72.585000 42.440000 ;
        RECT 72.385000 42.670000 72.585000 42.870000 ;
        RECT 72.385000 43.100000 72.585000 43.300000 ;
        RECT 72.385000 43.530000 72.585000 43.730000 ;
        RECT 72.385000 43.960000 72.585000 44.160000 ;
        RECT 72.790000 39.660000 72.990000 39.860000 ;
        RECT 72.790000 40.090000 72.990000 40.290000 ;
        RECT 72.790000 40.520000 72.990000 40.720000 ;
        RECT 72.790000 40.950000 72.990000 41.150000 ;
        RECT 72.790000 41.380000 72.990000 41.580000 ;
        RECT 72.790000 41.810000 72.990000 42.010000 ;
        RECT 72.790000 42.240000 72.990000 42.440000 ;
        RECT 72.790000 42.670000 72.990000 42.870000 ;
        RECT 72.790000 43.100000 72.990000 43.300000 ;
        RECT 72.790000 43.530000 72.990000 43.730000 ;
        RECT 72.790000 43.960000 72.990000 44.160000 ;
        RECT 73.195000 39.660000 73.395000 39.860000 ;
        RECT 73.195000 40.090000 73.395000 40.290000 ;
        RECT 73.195000 40.520000 73.395000 40.720000 ;
        RECT 73.195000 40.950000 73.395000 41.150000 ;
        RECT 73.195000 41.380000 73.395000 41.580000 ;
        RECT 73.195000 41.810000 73.395000 42.010000 ;
        RECT 73.195000 42.240000 73.395000 42.440000 ;
        RECT 73.195000 42.670000 73.395000 42.870000 ;
        RECT 73.195000 43.100000 73.395000 43.300000 ;
        RECT 73.195000 43.530000 73.395000 43.730000 ;
        RECT 73.195000 43.960000 73.395000 44.160000 ;
        RECT 73.600000 39.660000 73.800000 39.860000 ;
        RECT 73.600000 40.090000 73.800000 40.290000 ;
        RECT 73.600000 40.520000 73.800000 40.720000 ;
        RECT 73.600000 40.950000 73.800000 41.150000 ;
        RECT 73.600000 41.380000 73.800000 41.580000 ;
        RECT 73.600000 41.810000 73.800000 42.010000 ;
        RECT 73.600000 42.240000 73.800000 42.440000 ;
        RECT 73.600000 42.670000 73.800000 42.870000 ;
        RECT 73.600000 43.100000 73.800000 43.300000 ;
        RECT 73.600000 43.530000 73.800000 43.730000 ;
        RECT 73.600000 43.960000 73.800000 44.160000 ;
        RECT 74.005000 39.660000 74.205000 39.860000 ;
        RECT 74.005000 40.090000 74.205000 40.290000 ;
        RECT 74.005000 40.520000 74.205000 40.720000 ;
        RECT 74.005000 40.950000 74.205000 41.150000 ;
        RECT 74.005000 41.380000 74.205000 41.580000 ;
        RECT 74.005000 41.810000 74.205000 42.010000 ;
        RECT 74.005000 42.240000 74.205000 42.440000 ;
        RECT 74.005000 42.670000 74.205000 42.870000 ;
        RECT 74.005000 43.100000 74.205000 43.300000 ;
        RECT 74.005000 43.530000 74.205000 43.730000 ;
        RECT 74.005000 43.960000 74.205000 44.160000 ;
        RECT 74.410000 39.660000 74.610000 39.860000 ;
        RECT 74.410000 40.090000 74.610000 40.290000 ;
        RECT 74.410000 40.520000 74.610000 40.720000 ;
        RECT 74.410000 40.950000 74.610000 41.150000 ;
        RECT 74.410000 41.380000 74.610000 41.580000 ;
        RECT 74.410000 41.810000 74.610000 42.010000 ;
        RECT 74.410000 42.240000 74.610000 42.440000 ;
        RECT 74.410000 42.670000 74.610000 42.870000 ;
        RECT 74.410000 43.100000 74.610000 43.300000 ;
        RECT 74.410000 43.530000 74.610000 43.730000 ;
        RECT 74.410000 43.960000 74.610000 44.160000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 75.000000  39.190000 ;
      RECT  0.000000 44.630000 75.000000 198.000000 ;
      RECT 24.900000 39.190000 50.355000  44.630000 ;
    LAYER met4 ;
      RECT  0.000000   5.885000  1.670000   6.485000 ;
      RECT  0.000000  11.935000  1.365000  12.535000 ;
      RECT  0.000000  16.785000  1.365000  17.385000 ;
      RECT  0.000000  22.835000  1.670000  23.435000 ;
      RECT  0.000000  28.885000  1.670000  29.485000 ;
      RECT  0.000000  33.735000  1.670000  34.335000 ;
      RECT  0.000000  38.585000  1.670000  39.185000 ;
      RECT  0.000000  44.635000  1.670000  45.335000 ;
      RECT  0.000000  55.135000  1.670000  55.835000 ;
      RECT  0.000000  61.085000  1.670000  61.685000 ;
      RECT  0.000000  66.935000  1.670000  67.635000 ;
      RECT  0.000000  93.400000 75.000000 173.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.670000   0.000000 73.330000  11.935000 ;
      RECT  1.670000  17.385000 73.330000  39.185000 ;
      RECT  1.670000  44.635000 73.330000  93.400000 ;
      RECT  1.670000 173.385000 73.330000 198.000000 ;
      RECT 24.875000  39.185000 50.380000  44.635000 ;
      RECT 73.330000   5.885000 75.000000   6.485000 ;
      RECT 73.330000  22.835000 75.000000  23.435000 ;
      RECT 73.330000  28.885000 75.000000  29.485000 ;
      RECT 73.330000  33.735000 75.000000  34.335000 ;
      RECT 73.330000  38.585000 75.000000  39.185000 ;
      RECT 73.330000  44.635000 75.000000  45.335000 ;
      RECT 73.330000  55.135000 75.000000  55.835000 ;
      RECT 73.330000  61.085000 75.000000  61.685000 ;
      RECT 73.330000  66.935000 75.000000  67.635000 ;
      RECT 73.635000  11.935000 75.000000  12.535000 ;
      RECT 73.635000  16.785000 75.000000  17.385000 ;
    LAYER met5 ;
      RECT 0.000000  93.785000 75.000000 172.985000 ;
      RECT 1.765000  12.235000 73.235000  17.085000 ;
      RECT 2.070000   0.000000 72.930000  12.235000 ;
      RECT 2.070000  17.085000 72.930000  93.785000 ;
      RECT 2.070000 172.985000 72.930000 198.000000 ;
  END
END sky130_fd_io__overlay_vssd_lvc


MACRO sky130_fd_io__overlay_gpiov2
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 80 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 53.125000 80.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 48.365000 80.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN PAD
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 31.870000 127.605000 53.410000 149.150000 ;
    END
  END PAD
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT  0.000000  8.885000  1.270000  9.105000 ;
        RECT  0.000000  9.105000 80.000000 13.315000 ;
        RECT  0.000000 13.315000  1.270000 13.535000 ;
        RECT 78.730000  8.885000 80.000000  9.105000 ;
        RECT 78.730000 13.315000 80.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 80.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT  0.000000 2.035000  1.270000 2.255000 ;
        RECT  0.000000 2.255000 80.000000 7.265000 ;
        RECT  0.000000 7.265000  1.270000 7.485000 ;
        RECT 78.730000 2.035000 80.000000 2.255000 ;
        RECT 78.730000 7.265000 80.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 80.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000  0.965000 15.155000 ;
        RECT 0.000000 15.155000 78.970000 18.165000 ;
        RECT 0.000000 18.165000  0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.035000 14.935000 80.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 80.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT  0.000000 19.785000  1.270000 20.005000 ;
        RECT  0.000000 20.005000 80.000000 24.215000 ;
        RECT  0.000000 24.215000  1.270000 24.435000 ;
        RECT 78.730000 19.785000 80.000000 20.005000 ;
        RECT 78.730000 24.215000 80.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT  0.000000 70.035000  1.270000 70.155000 ;
        RECT  0.000000 70.155000 80.000000 94.865000 ;
        RECT  0.000000 94.865000  1.270000 95.000000 ;
        RECT 78.730000 70.035000 80.000000 70.155000 ;
        RECT 78.730000 94.865000 80.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 80.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 80.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT  0.000000 64.085000  1.270000 64.305000 ;
        RECT  0.000000 64.305000 80.000000 68.315000 ;
        RECT  0.000000 68.315000  1.270000 68.535000 ;
        RECT 78.730000 64.085000 80.000000 64.305000 ;
        RECT 78.730000 68.315000 80.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 80.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT  0.000000 36.735000  1.270000 36.955000 ;
        RECT  0.000000 36.955000 80.000000 39.965000 ;
        RECT  0.000000 39.965000  1.270000 40.185000 ;
        RECT 78.730000 36.735000 80.000000 36.955000 ;
        RECT 78.730000 39.965000 80.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 80.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 47.735000 80.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 56.405000 80.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.835000 80.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 80.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT  0.000000 41.585000  1.270000 41.805000 ;
        RECT  0.000000 41.805000 80.000000 46.015000 ;
        RECT  0.000000 46.015000  1.270000 46.235000 ;
        RECT 78.730000 41.585000 80.000000 41.805000 ;
        RECT 78.730000 46.015000 80.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 80.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT  0.000000 175.785000  1.270000 175.910000 ;
        RECT  0.000000 175.910000 80.000000 199.880000 ;
        RECT  0.000000 199.880000  1.270000 200.000000 ;
        RECT 78.730000 175.785000 80.000000 175.910000 ;
        RECT 78.730000 199.880000 80.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT  0.000000 25.835000  1.270000 26.055000 ;
        RECT  0.000000 26.055000 80.000000 30.265000 ;
        RECT  0.000000 30.265000  1.270000 30.485000 ;
        RECT 78.730000 25.835000 80.000000 26.055000 ;
        RECT 78.730000 30.265000 80.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 80.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 80.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT  0.000000 58.235000  1.270000 58.455000 ;
        RECT  0.000000 58.455000 80.000000 62.465000 ;
        RECT  0.000000 62.465000  1.270000 62.685000 ;
        RECT 78.730000 58.235000 80.000000 58.455000 ;
        RECT 78.730000 62.465000 80.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 80.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT  0.000000 31.885000  1.270000 32.105000 ;
        RECT  0.000000 32.105000 80.000000 35.115000 ;
        RECT  0.000000 35.115000  1.270000 35.335000 ;
        RECT 78.730000 31.885000 80.000000 32.105000 ;
        RECT 78.730000 35.115000 80.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 80.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER via4 ;
      RECT  0.995000  20.195000  1.795000  20.995000 ;
      RECT  0.995000  23.225000  1.795000  24.025000 ;
      RECT  0.995000  26.245000  1.795000  27.045000 ;
      RECT  0.995000  29.275000  1.795000  30.075000 ;
      RECT  1.000000   2.450000  1.800000   3.250000 ;
      RECT  1.000000   4.360000  1.800000   5.160000 ;
      RECT  1.000000   6.270000  1.800000   7.070000 ;
      RECT  1.000000  15.345000  1.800000  16.145000 ;
      RECT  1.000000  17.175000  1.800000  17.975000 ;
      RECT  1.000000  32.295000  1.800000  33.095000 ;
      RECT  1.000000  34.125000  1.800000  34.925000 ;
      RECT  1.000000  37.145000  1.800000  37.945000 ;
      RECT  1.000000  38.975000  1.800000  39.775000 ;
      RECT  1.000000  41.995000  1.800000  42.795000 ;
      RECT  1.000000  45.025000  1.800000  45.825000 ;
      RECT  1.000000  51.835000  1.800000  52.635000 ;
      RECT  1.000000  58.645000  1.800000  59.445000 ;
      RECT  1.000000  61.475000  1.800000  62.275000 ;
      RECT  1.000000  64.495000  1.800000  65.295000 ;
      RECT  1.000000  67.325000  1.800000  68.125000 ;
      RECT  1.000000  70.350000  1.800000  71.150000 ;
      RECT  1.000000  72.030000  1.800000  72.830000 ;
      RECT  1.000000  73.710000  1.800000  74.510000 ;
      RECT  1.000000  75.390000  1.800000  76.190000 ;
      RECT  1.000000  77.070000  1.800000  77.870000 ;
      RECT  1.000000  78.750000  1.800000  79.550000 ;
      RECT  1.000000  80.430000  1.800000  81.230000 ;
      RECT  1.000000  82.110000  1.800000  82.910000 ;
      RECT  1.000000  83.790000  1.800000  84.590000 ;
      RECT  1.000000  85.470000  1.800000  86.270000 ;
      RECT  1.000000  87.150000  1.800000  87.950000 ;
      RECT  1.000000  88.830000  1.800000  89.630000 ;
      RECT  1.000000  90.510000  1.800000  91.310000 ;
      RECT  1.000000  92.190000  1.800000  92.990000 ;
      RECT  1.000000  93.870000  1.800000  94.670000 ;
      RECT  1.000000 176.155000  1.800000 176.955000 ;
      RECT  1.000000 177.775000  1.800000 178.575000 ;
      RECT  1.000000 179.395000  1.800000 180.195000 ;
      RECT  1.000000 181.015000  1.800000 181.815000 ;
      RECT  1.000000 182.635000  1.800000 183.435000 ;
      RECT  1.000000 184.255000  1.800000 185.055000 ;
      RECT  1.000000 185.875000  1.800000 186.675000 ;
      RECT  1.000000 187.495000  1.800000 188.295000 ;
      RECT  1.000000 189.115000  1.800000 189.915000 ;
      RECT  1.000000 190.735000  1.800000 191.535000 ;
      RECT  1.000000 192.355000  1.800000 193.155000 ;
      RECT  1.000000 193.975000  1.800000 194.775000 ;
      RECT  1.000000 195.595000  1.800000 196.395000 ;
      RECT  1.000000 197.215000  1.800000 198.015000 ;
      RECT  1.000000 198.835000  1.800000 199.635000 ;
      RECT  1.005000   9.295000  1.805000  10.095000 ;
      RECT  1.005000  12.325000  1.805000  13.125000 ;
      RECT  2.600000  20.195000  3.400000  20.995000 ;
      RECT  2.600000  23.225000  3.400000  24.025000 ;
      RECT  2.600000  26.245000  3.400000  27.045000 ;
      RECT  2.600000  29.275000  3.400000  30.075000 ;
      RECT  2.605000   2.450000  3.405000   3.250000 ;
      RECT  2.605000   4.360000  3.405000   5.160000 ;
      RECT  2.605000   6.270000  3.405000   7.070000 ;
      RECT  2.605000  15.345000  3.405000  16.145000 ;
      RECT  2.605000  17.175000  3.405000  17.975000 ;
      RECT  2.605000  32.295000  3.405000  33.095000 ;
      RECT  2.605000  34.125000  3.405000  34.925000 ;
      RECT  2.605000  37.145000  3.405000  37.945000 ;
      RECT  2.605000  38.975000  3.405000  39.775000 ;
      RECT  2.605000  41.995000  3.405000  42.795000 ;
      RECT  2.605000  45.025000  3.405000  45.825000 ;
      RECT  2.605000  51.835000  3.405000  52.635000 ;
      RECT  2.605000  58.645000  3.405000  59.445000 ;
      RECT  2.605000  61.475000  3.405000  62.275000 ;
      RECT  2.605000  64.495000  3.405000  65.295000 ;
      RECT  2.605000  67.325000  3.405000  68.125000 ;
      RECT  2.605000  70.350000  3.405000  71.150000 ;
      RECT  2.605000  72.030000  3.405000  72.830000 ;
      RECT  2.605000  73.710000  3.405000  74.510000 ;
      RECT  2.605000  75.390000  3.405000  76.190000 ;
      RECT  2.605000  77.070000  3.405000  77.870000 ;
      RECT  2.605000  78.750000  3.405000  79.550000 ;
      RECT  2.605000  80.430000  3.405000  81.230000 ;
      RECT  2.605000  82.110000  3.405000  82.910000 ;
      RECT  2.605000  83.790000  3.405000  84.590000 ;
      RECT  2.605000  85.470000  3.405000  86.270000 ;
      RECT  2.605000  87.150000  3.405000  87.950000 ;
      RECT  2.605000  88.830000  3.405000  89.630000 ;
      RECT  2.605000  90.510000  3.405000  91.310000 ;
      RECT  2.605000  92.190000  3.405000  92.990000 ;
      RECT  2.605000  93.870000  3.405000  94.670000 ;
      RECT  2.605000 176.155000  3.405000 176.955000 ;
      RECT  2.605000 177.775000  3.405000 178.575000 ;
      RECT  2.605000 179.395000  3.405000 180.195000 ;
      RECT  2.605000 181.015000  3.405000 181.815000 ;
      RECT  2.605000 182.635000  3.405000 183.435000 ;
      RECT  2.605000 184.255000  3.405000 185.055000 ;
      RECT  2.605000 185.875000  3.405000 186.675000 ;
      RECT  2.605000 187.495000  3.405000 188.295000 ;
      RECT  2.605000 189.115000  3.405000 189.915000 ;
      RECT  2.605000 190.735000  3.405000 191.535000 ;
      RECT  2.605000 192.355000  3.405000 193.155000 ;
      RECT  2.605000 193.975000  3.405000 194.775000 ;
      RECT  2.605000 195.595000  3.405000 196.395000 ;
      RECT  2.605000 197.215000  3.405000 198.015000 ;
      RECT  2.605000 198.835000  3.405000 199.635000 ;
      RECT  2.610000   9.295000  3.410000  10.095000 ;
      RECT  2.610000  12.325000  3.410000  13.125000 ;
      RECT  4.205000  20.195000  5.005000  20.995000 ;
      RECT  4.205000  23.225000  5.005000  24.025000 ;
      RECT  4.205000  26.245000  5.005000  27.045000 ;
      RECT  4.205000  29.275000  5.005000  30.075000 ;
      RECT  4.210000   2.450000  5.010000   3.250000 ;
      RECT  4.210000   4.360000  5.010000   5.160000 ;
      RECT  4.210000   6.270000  5.010000   7.070000 ;
      RECT  4.210000  15.345000  5.010000  16.145000 ;
      RECT  4.210000  17.175000  5.010000  17.975000 ;
      RECT  4.210000  32.295000  5.010000  33.095000 ;
      RECT  4.210000  34.125000  5.010000  34.925000 ;
      RECT  4.210000  37.145000  5.010000  37.945000 ;
      RECT  4.210000  38.975000  5.010000  39.775000 ;
      RECT  4.210000  41.995000  5.010000  42.795000 ;
      RECT  4.210000  45.025000  5.010000  45.825000 ;
      RECT  4.210000  51.835000  5.010000  52.635000 ;
      RECT  4.210000  58.645000  5.010000  59.445000 ;
      RECT  4.210000  61.475000  5.010000  62.275000 ;
      RECT  4.210000  64.495000  5.010000  65.295000 ;
      RECT  4.210000  67.325000  5.010000  68.125000 ;
      RECT  4.210000  70.350000  5.010000  71.150000 ;
      RECT  4.210000  72.030000  5.010000  72.830000 ;
      RECT  4.210000  73.710000  5.010000  74.510000 ;
      RECT  4.210000  75.390000  5.010000  76.190000 ;
      RECT  4.210000  77.070000  5.010000  77.870000 ;
      RECT  4.210000  78.750000  5.010000  79.550000 ;
      RECT  4.210000  80.430000  5.010000  81.230000 ;
      RECT  4.210000  82.110000  5.010000  82.910000 ;
      RECT  4.210000  83.790000  5.010000  84.590000 ;
      RECT  4.210000  85.470000  5.010000  86.270000 ;
      RECT  4.210000  87.150000  5.010000  87.950000 ;
      RECT  4.210000  88.830000  5.010000  89.630000 ;
      RECT  4.210000  90.510000  5.010000  91.310000 ;
      RECT  4.210000  92.190000  5.010000  92.990000 ;
      RECT  4.210000  93.870000  5.010000  94.670000 ;
      RECT  4.210000 176.155000  5.010000 176.955000 ;
      RECT  4.210000 177.775000  5.010000 178.575000 ;
      RECT  4.210000 179.395000  5.010000 180.195000 ;
      RECT  4.210000 181.015000  5.010000 181.815000 ;
      RECT  4.210000 182.635000  5.010000 183.435000 ;
      RECT  4.210000 184.255000  5.010000 185.055000 ;
      RECT  4.210000 185.875000  5.010000 186.675000 ;
      RECT  4.210000 187.495000  5.010000 188.295000 ;
      RECT  4.210000 189.115000  5.010000 189.915000 ;
      RECT  4.210000 190.735000  5.010000 191.535000 ;
      RECT  4.210000 192.355000  5.010000 193.155000 ;
      RECT  4.210000 193.975000  5.010000 194.775000 ;
      RECT  4.210000 195.595000  5.010000 196.395000 ;
      RECT  4.210000 197.215000  5.010000 198.015000 ;
      RECT  4.210000 198.835000  5.010000 199.635000 ;
      RECT  4.215000   9.295000  5.015000  10.095000 ;
      RECT  4.215000  12.325000  5.015000  13.125000 ;
      RECT  5.810000  20.195000  6.610000  20.995000 ;
      RECT  5.810000  23.225000  6.610000  24.025000 ;
      RECT  5.810000  26.245000  6.610000  27.045000 ;
      RECT  5.810000  29.275000  6.610000  30.075000 ;
      RECT  5.815000   2.450000  6.615000   3.250000 ;
      RECT  5.815000   4.360000  6.615000   5.160000 ;
      RECT  5.815000   6.270000  6.615000   7.070000 ;
      RECT  5.815000  15.345000  6.615000  16.145000 ;
      RECT  5.815000  17.175000  6.615000  17.975000 ;
      RECT  5.815000  32.295000  6.615000  33.095000 ;
      RECT  5.815000  34.125000  6.615000  34.925000 ;
      RECT  5.815000  37.145000  6.615000  37.945000 ;
      RECT  5.815000  38.975000  6.615000  39.775000 ;
      RECT  5.815000  41.995000  6.615000  42.795000 ;
      RECT  5.815000  45.025000  6.615000  45.825000 ;
      RECT  5.815000  51.835000  6.615000  52.635000 ;
      RECT  5.815000  58.645000  6.615000  59.445000 ;
      RECT  5.815000  61.475000  6.615000  62.275000 ;
      RECT  5.815000  64.495000  6.615000  65.295000 ;
      RECT  5.815000  67.325000  6.615000  68.125000 ;
      RECT  5.815000  70.350000  6.615000  71.150000 ;
      RECT  5.815000  72.030000  6.615000  72.830000 ;
      RECT  5.815000  73.710000  6.615000  74.510000 ;
      RECT  5.815000  75.390000  6.615000  76.190000 ;
      RECT  5.815000  77.070000  6.615000  77.870000 ;
      RECT  5.815000  78.750000  6.615000  79.550000 ;
      RECT  5.815000  80.430000  6.615000  81.230000 ;
      RECT  5.815000  82.110000  6.615000  82.910000 ;
      RECT  5.815000  83.790000  6.615000  84.590000 ;
      RECT  5.815000  85.470000  6.615000  86.270000 ;
      RECT  5.815000  87.150000  6.615000  87.950000 ;
      RECT  5.815000  88.830000  6.615000  89.630000 ;
      RECT  5.815000  90.510000  6.615000  91.310000 ;
      RECT  5.815000  92.190000  6.615000  92.990000 ;
      RECT  5.815000  93.870000  6.615000  94.670000 ;
      RECT  5.815000 176.155000  6.615000 176.955000 ;
      RECT  5.815000 177.775000  6.615000 178.575000 ;
      RECT  5.815000 179.395000  6.615000 180.195000 ;
      RECT  5.815000 181.015000  6.615000 181.815000 ;
      RECT  5.815000 182.635000  6.615000 183.435000 ;
      RECT  5.815000 184.255000  6.615000 185.055000 ;
      RECT  5.815000 185.875000  6.615000 186.675000 ;
      RECT  5.815000 187.495000  6.615000 188.295000 ;
      RECT  5.815000 189.115000  6.615000 189.915000 ;
      RECT  5.815000 190.735000  6.615000 191.535000 ;
      RECT  5.815000 192.355000  6.615000 193.155000 ;
      RECT  5.815000 193.975000  6.615000 194.775000 ;
      RECT  5.815000 195.595000  6.615000 196.395000 ;
      RECT  5.815000 197.215000  6.615000 198.015000 ;
      RECT  5.815000 198.835000  6.615000 199.635000 ;
      RECT  5.820000   9.295000  6.620000  10.095000 ;
      RECT  5.820000  12.325000  6.620000  13.125000 ;
      RECT  7.415000  20.195000  8.215000  20.995000 ;
      RECT  7.415000  23.225000  8.215000  24.025000 ;
      RECT  7.415000  26.245000  8.215000  27.045000 ;
      RECT  7.415000  29.275000  8.215000  30.075000 ;
      RECT  7.420000   2.450000  8.220000   3.250000 ;
      RECT  7.420000   4.360000  8.220000   5.160000 ;
      RECT  7.420000   6.270000  8.220000   7.070000 ;
      RECT  7.420000  15.345000  8.220000  16.145000 ;
      RECT  7.420000  17.175000  8.220000  17.975000 ;
      RECT  7.420000  32.295000  8.220000  33.095000 ;
      RECT  7.420000  34.125000  8.220000  34.925000 ;
      RECT  7.420000  37.145000  8.220000  37.945000 ;
      RECT  7.420000  38.975000  8.220000  39.775000 ;
      RECT  7.420000  41.995000  8.220000  42.795000 ;
      RECT  7.420000  45.025000  8.220000  45.825000 ;
      RECT  7.420000  51.835000  8.220000  52.635000 ;
      RECT  7.420000  58.645000  8.220000  59.445000 ;
      RECT  7.420000  61.475000  8.220000  62.275000 ;
      RECT  7.420000  64.495000  8.220000  65.295000 ;
      RECT  7.420000  67.325000  8.220000  68.125000 ;
      RECT  7.420000  70.350000  8.220000  71.150000 ;
      RECT  7.420000  72.030000  8.220000  72.830000 ;
      RECT  7.420000  73.710000  8.220000  74.510000 ;
      RECT  7.420000  75.390000  8.220000  76.190000 ;
      RECT  7.420000  77.070000  8.220000  77.870000 ;
      RECT  7.420000  78.750000  8.220000  79.550000 ;
      RECT  7.420000  80.430000  8.220000  81.230000 ;
      RECT  7.420000  82.110000  8.220000  82.910000 ;
      RECT  7.420000  83.790000  8.220000  84.590000 ;
      RECT  7.420000  85.470000  8.220000  86.270000 ;
      RECT  7.420000  87.150000  8.220000  87.950000 ;
      RECT  7.420000  88.830000  8.220000  89.630000 ;
      RECT  7.420000  90.510000  8.220000  91.310000 ;
      RECT  7.420000  92.190000  8.220000  92.990000 ;
      RECT  7.420000  93.870000  8.220000  94.670000 ;
      RECT  7.420000 176.155000  8.220000 176.955000 ;
      RECT  7.420000 177.775000  8.220000 178.575000 ;
      RECT  7.420000 179.395000  8.220000 180.195000 ;
      RECT  7.420000 181.015000  8.220000 181.815000 ;
      RECT  7.420000 182.635000  8.220000 183.435000 ;
      RECT  7.420000 184.255000  8.220000 185.055000 ;
      RECT  7.420000 185.875000  8.220000 186.675000 ;
      RECT  7.420000 187.495000  8.220000 188.295000 ;
      RECT  7.420000 189.115000  8.220000 189.915000 ;
      RECT  7.420000 190.735000  8.220000 191.535000 ;
      RECT  7.420000 192.355000  8.220000 193.155000 ;
      RECT  7.420000 193.975000  8.220000 194.775000 ;
      RECT  7.420000 195.595000  8.220000 196.395000 ;
      RECT  7.420000 197.215000  8.220000 198.015000 ;
      RECT  7.420000 198.835000  8.220000 199.635000 ;
      RECT  7.425000   9.295000  8.225000  10.095000 ;
      RECT  7.425000  12.325000  8.225000  13.125000 ;
      RECT  9.020000  20.195000  9.820000  20.995000 ;
      RECT  9.020000  23.225000  9.820000  24.025000 ;
      RECT  9.020000  26.245000  9.820000  27.045000 ;
      RECT  9.020000  29.275000  9.820000  30.075000 ;
      RECT  9.025000   2.450000  9.825000   3.250000 ;
      RECT  9.025000   4.360000  9.825000   5.160000 ;
      RECT  9.025000   6.270000  9.825000   7.070000 ;
      RECT  9.025000  15.345000  9.825000  16.145000 ;
      RECT  9.025000  17.175000  9.825000  17.975000 ;
      RECT  9.025000  32.295000  9.825000  33.095000 ;
      RECT  9.025000  34.125000  9.825000  34.925000 ;
      RECT  9.025000  37.145000  9.825000  37.945000 ;
      RECT  9.025000  38.975000  9.825000  39.775000 ;
      RECT  9.025000  41.995000  9.825000  42.795000 ;
      RECT  9.025000  45.025000  9.825000  45.825000 ;
      RECT  9.025000  51.835000  9.825000  52.635000 ;
      RECT  9.025000  58.645000  9.825000  59.445000 ;
      RECT  9.025000  61.475000  9.825000  62.275000 ;
      RECT  9.025000  64.495000  9.825000  65.295000 ;
      RECT  9.025000  67.325000  9.825000  68.125000 ;
      RECT  9.025000  70.350000  9.825000  71.150000 ;
      RECT  9.025000  72.030000  9.825000  72.830000 ;
      RECT  9.025000  73.710000  9.825000  74.510000 ;
      RECT  9.025000  75.390000  9.825000  76.190000 ;
      RECT  9.025000  77.070000  9.825000  77.870000 ;
      RECT  9.025000  78.750000  9.825000  79.550000 ;
      RECT  9.025000  80.430000  9.825000  81.230000 ;
      RECT  9.025000  82.110000  9.825000  82.910000 ;
      RECT  9.025000  83.790000  9.825000  84.590000 ;
      RECT  9.025000  85.470000  9.825000  86.270000 ;
      RECT  9.025000  87.150000  9.825000  87.950000 ;
      RECT  9.025000  88.830000  9.825000  89.630000 ;
      RECT  9.025000  90.510000  9.825000  91.310000 ;
      RECT  9.025000  92.190000  9.825000  92.990000 ;
      RECT  9.025000  93.870000  9.825000  94.670000 ;
      RECT  9.025000 176.155000  9.825000 176.955000 ;
      RECT  9.025000 177.775000  9.825000 178.575000 ;
      RECT  9.025000 179.395000  9.825000 180.195000 ;
      RECT  9.025000 181.015000  9.825000 181.815000 ;
      RECT  9.025000 182.635000  9.825000 183.435000 ;
      RECT  9.025000 184.255000  9.825000 185.055000 ;
      RECT  9.025000 185.875000  9.825000 186.675000 ;
      RECT  9.025000 187.495000  9.825000 188.295000 ;
      RECT  9.025000 189.115000  9.825000 189.915000 ;
      RECT  9.025000 190.735000  9.825000 191.535000 ;
      RECT  9.025000 192.355000  9.825000 193.155000 ;
      RECT  9.025000 193.975000  9.825000 194.775000 ;
      RECT  9.025000 195.595000  9.825000 196.395000 ;
      RECT  9.025000 197.215000  9.825000 198.015000 ;
      RECT  9.025000 198.835000  9.825000 199.635000 ;
      RECT  9.030000   9.295000  9.830000  10.095000 ;
      RECT  9.030000  12.325000  9.830000  13.125000 ;
      RECT 10.625000  20.195000 11.425000  20.995000 ;
      RECT 10.625000  23.225000 11.425000  24.025000 ;
      RECT 10.625000  26.245000 11.425000  27.045000 ;
      RECT 10.625000  29.275000 11.425000  30.075000 ;
      RECT 10.630000   2.450000 11.430000   3.250000 ;
      RECT 10.630000   4.360000 11.430000   5.160000 ;
      RECT 10.630000   6.270000 11.430000   7.070000 ;
      RECT 10.630000  15.345000 11.430000  16.145000 ;
      RECT 10.630000  17.175000 11.430000  17.975000 ;
      RECT 10.630000  32.295000 11.430000  33.095000 ;
      RECT 10.630000  34.125000 11.430000  34.925000 ;
      RECT 10.630000  37.145000 11.430000  37.945000 ;
      RECT 10.630000  38.975000 11.430000  39.775000 ;
      RECT 10.630000  41.995000 11.430000  42.795000 ;
      RECT 10.630000  45.025000 11.430000  45.825000 ;
      RECT 10.630000  51.835000 11.430000  52.635000 ;
      RECT 10.630000  58.645000 11.430000  59.445000 ;
      RECT 10.630000  61.475000 11.430000  62.275000 ;
      RECT 10.630000  64.495000 11.430000  65.295000 ;
      RECT 10.630000  67.325000 11.430000  68.125000 ;
      RECT 10.630000  70.350000 11.430000  71.150000 ;
      RECT 10.630000  72.030000 11.430000  72.830000 ;
      RECT 10.630000  73.710000 11.430000  74.510000 ;
      RECT 10.630000  75.390000 11.430000  76.190000 ;
      RECT 10.630000  77.070000 11.430000  77.870000 ;
      RECT 10.630000  78.750000 11.430000  79.550000 ;
      RECT 10.630000  80.430000 11.430000  81.230000 ;
      RECT 10.630000  82.110000 11.430000  82.910000 ;
      RECT 10.630000  83.790000 11.430000  84.590000 ;
      RECT 10.630000  85.470000 11.430000  86.270000 ;
      RECT 10.630000  87.150000 11.430000  87.950000 ;
      RECT 10.630000  88.830000 11.430000  89.630000 ;
      RECT 10.630000  90.510000 11.430000  91.310000 ;
      RECT 10.630000  92.190000 11.430000  92.990000 ;
      RECT 10.630000  93.870000 11.430000  94.670000 ;
      RECT 10.630000 176.155000 11.430000 176.955000 ;
      RECT 10.630000 177.775000 11.430000 178.575000 ;
      RECT 10.630000 179.395000 11.430000 180.195000 ;
      RECT 10.630000 181.015000 11.430000 181.815000 ;
      RECT 10.630000 182.635000 11.430000 183.435000 ;
      RECT 10.630000 184.255000 11.430000 185.055000 ;
      RECT 10.630000 185.875000 11.430000 186.675000 ;
      RECT 10.630000 187.495000 11.430000 188.295000 ;
      RECT 10.630000 189.115000 11.430000 189.915000 ;
      RECT 10.630000 190.735000 11.430000 191.535000 ;
      RECT 10.630000 192.355000 11.430000 193.155000 ;
      RECT 10.630000 193.975000 11.430000 194.775000 ;
      RECT 10.630000 195.595000 11.430000 196.395000 ;
      RECT 10.630000 197.215000 11.430000 198.015000 ;
      RECT 10.630000 198.835000 11.430000 199.635000 ;
      RECT 10.635000   9.295000 11.435000  10.095000 ;
      RECT 10.635000  12.325000 11.435000  13.125000 ;
      RECT 12.230000  20.195000 13.030000  20.995000 ;
      RECT 12.230000  23.225000 13.030000  24.025000 ;
      RECT 12.230000  26.245000 13.030000  27.045000 ;
      RECT 12.230000  29.275000 13.030000  30.075000 ;
      RECT 12.235000   2.450000 13.035000   3.250000 ;
      RECT 12.235000   4.360000 13.035000   5.160000 ;
      RECT 12.235000   6.270000 13.035000   7.070000 ;
      RECT 12.235000  15.345000 13.035000  16.145000 ;
      RECT 12.235000  17.175000 13.035000  17.975000 ;
      RECT 12.235000  32.295000 13.035000  33.095000 ;
      RECT 12.235000  34.125000 13.035000  34.925000 ;
      RECT 12.235000  37.145000 13.035000  37.945000 ;
      RECT 12.235000  38.975000 13.035000  39.775000 ;
      RECT 12.235000  41.995000 13.035000  42.795000 ;
      RECT 12.235000  45.025000 13.035000  45.825000 ;
      RECT 12.235000  51.835000 13.035000  52.635000 ;
      RECT 12.235000  58.645000 13.035000  59.445000 ;
      RECT 12.235000  61.475000 13.035000  62.275000 ;
      RECT 12.235000  64.495000 13.035000  65.295000 ;
      RECT 12.235000  67.325000 13.035000  68.125000 ;
      RECT 12.235000  70.350000 13.035000  71.150000 ;
      RECT 12.235000  72.030000 13.035000  72.830000 ;
      RECT 12.235000  73.710000 13.035000  74.510000 ;
      RECT 12.235000  75.390000 13.035000  76.190000 ;
      RECT 12.235000  77.070000 13.035000  77.870000 ;
      RECT 12.235000  78.750000 13.035000  79.550000 ;
      RECT 12.235000  80.430000 13.035000  81.230000 ;
      RECT 12.235000  82.110000 13.035000  82.910000 ;
      RECT 12.235000  83.790000 13.035000  84.590000 ;
      RECT 12.235000  85.470000 13.035000  86.270000 ;
      RECT 12.235000  87.150000 13.035000  87.950000 ;
      RECT 12.235000  88.830000 13.035000  89.630000 ;
      RECT 12.235000  90.510000 13.035000  91.310000 ;
      RECT 12.235000  92.190000 13.035000  92.990000 ;
      RECT 12.235000  93.870000 13.035000  94.670000 ;
      RECT 12.235000 176.155000 13.035000 176.955000 ;
      RECT 12.235000 177.775000 13.035000 178.575000 ;
      RECT 12.235000 179.395000 13.035000 180.195000 ;
      RECT 12.235000 181.015000 13.035000 181.815000 ;
      RECT 12.235000 182.635000 13.035000 183.435000 ;
      RECT 12.235000 184.255000 13.035000 185.055000 ;
      RECT 12.235000 185.875000 13.035000 186.675000 ;
      RECT 12.235000 187.495000 13.035000 188.295000 ;
      RECT 12.235000 189.115000 13.035000 189.915000 ;
      RECT 12.235000 190.735000 13.035000 191.535000 ;
      RECT 12.235000 192.355000 13.035000 193.155000 ;
      RECT 12.235000 193.975000 13.035000 194.775000 ;
      RECT 12.235000 195.595000 13.035000 196.395000 ;
      RECT 12.235000 197.215000 13.035000 198.015000 ;
      RECT 12.235000 198.835000 13.035000 199.635000 ;
      RECT 12.240000   9.295000 13.040000  10.095000 ;
      RECT 12.240000  12.325000 13.040000  13.125000 ;
      RECT 13.835000  20.195000 14.635000  20.995000 ;
      RECT 13.835000  23.225000 14.635000  24.025000 ;
      RECT 13.835000  26.245000 14.635000  27.045000 ;
      RECT 13.835000  29.275000 14.635000  30.075000 ;
      RECT 13.840000   2.450000 14.640000   3.250000 ;
      RECT 13.840000   4.360000 14.640000   5.160000 ;
      RECT 13.840000   6.270000 14.640000   7.070000 ;
      RECT 13.840000  15.345000 14.640000  16.145000 ;
      RECT 13.840000  17.175000 14.640000  17.975000 ;
      RECT 13.840000  32.295000 14.640000  33.095000 ;
      RECT 13.840000  34.125000 14.640000  34.925000 ;
      RECT 13.840000  37.145000 14.640000  37.945000 ;
      RECT 13.840000  38.975000 14.640000  39.775000 ;
      RECT 13.840000  41.995000 14.640000  42.795000 ;
      RECT 13.840000  45.025000 14.640000  45.825000 ;
      RECT 13.840000  51.835000 14.640000  52.635000 ;
      RECT 13.840000  58.645000 14.640000  59.445000 ;
      RECT 13.840000  61.475000 14.640000  62.275000 ;
      RECT 13.840000  64.495000 14.640000  65.295000 ;
      RECT 13.840000  67.325000 14.640000  68.125000 ;
      RECT 13.840000  70.350000 14.640000  71.150000 ;
      RECT 13.840000  72.030000 14.640000  72.830000 ;
      RECT 13.840000  73.710000 14.640000  74.510000 ;
      RECT 13.840000  75.390000 14.640000  76.190000 ;
      RECT 13.840000  77.070000 14.640000  77.870000 ;
      RECT 13.840000  78.750000 14.640000  79.550000 ;
      RECT 13.840000  80.430000 14.640000  81.230000 ;
      RECT 13.840000  82.110000 14.640000  82.910000 ;
      RECT 13.840000  83.790000 14.640000  84.590000 ;
      RECT 13.840000  85.470000 14.640000  86.270000 ;
      RECT 13.840000  87.150000 14.640000  87.950000 ;
      RECT 13.840000  88.830000 14.640000  89.630000 ;
      RECT 13.840000  90.510000 14.640000  91.310000 ;
      RECT 13.840000  92.190000 14.640000  92.990000 ;
      RECT 13.840000  93.870000 14.640000  94.670000 ;
      RECT 13.840000 176.155000 14.640000 176.955000 ;
      RECT 13.840000 177.775000 14.640000 178.575000 ;
      RECT 13.840000 179.395000 14.640000 180.195000 ;
      RECT 13.840000 181.015000 14.640000 181.815000 ;
      RECT 13.840000 182.635000 14.640000 183.435000 ;
      RECT 13.840000 184.255000 14.640000 185.055000 ;
      RECT 13.840000 185.875000 14.640000 186.675000 ;
      RECT 13.840000 187.495000 14.640000 188.295000 ;
      RECT 13.840000 189.115000 14.640000 189.915000 ;
      RECT 13.840000 190.735000 14.640000 191.535000 ;
      RECT 13.840000 192.355000 14.640000 193.155000 ;
      RECT 13.840000 193.975000 14.640000 194.775000 ;
      RECT 13.840000 195.595000 14.640000 196.395000 ;
      RECT 13.840000 197.215000 14.640000 198.015000 ;
      RECT 13.840000 198.835000 14.640000 199.635000 ;
      RECT 13.845000   9.295000 14.645000  10.095000 ;
      RECT 13.845000  12.325000 14.645000  13.125000 ;
      RECT 15.440000  20.195000 16.240000  20.995000 ;
      RECT 15.440000  23.225000 16.240000  24.025000 ;
      RECT 15.440000  26.245000 16.240000  27.045000 ;
      RECT 15.440000  29.275000 16.240000  30.075000 ;
      RECT 15.445000   2.450000 16.245000   3.250000 ;
      RECT 15.445000   4.360000 16.245000   5.160000 ;
      RECT 15.445000   6.270000 16.245000   7.070000 ;
      RECT 15.445000  15.345000 16.245000  16.145000 ;
      RECT 15.445000  17.175000 16.245000  17.975000 ;
      RECT 15.445000  32.295000 16.245000  33.095000 ;
      RECT 15.445000  34.125000 16.245000  34.925000 ;
      RECT 15.445000  37.145000 16.245000  37.945000 ;
      RECT 15.445000  38.975000 16.245000  39.775000 ;
      RECT 15.445000  41.995000 16.245000  42.795000 ;
      RECT 15.445000  45.025000 16.245000  45.825000 ;
      RECT 15.445000  51.835000 16.245000  52.635000 ;
      RECT 15.445000  58.645000 16.245000  59.445000 ;
      RECT 15.445000  61.475000 16.245000  62.275000 ;
      RECT 15.445000  64.495000 16.245000  65.295000 ;
      RECT 15.445000  67.325000 16.245000  68.125000 ;
      RECT 15.445000  70.350000 16.245000  71.150000 ;
      RECT 15.445000  72.030000 16.245000  72.830000 ;
      RECT 15.445000  73.710000 16.245000  74.510000 ;
      RECT 15.445000  75.390000 16.245000  76.190000 ;
      RECT 15.445000  77.070000 16.245000  77.870000 ;
      RECT 15.445000  78.750000 16.245000  79.550000 ;
      RECT 15.445000  80.430000 16.245000  81.230000 ;
      RECT 15.445000  82.110000 16.245000  82.910000 ;
      RECT 15.445000  83.790000 16.245000  84.590000 ;
      RECT 15.445000  85.470000 16.245000  86.270000 ;
      RECT 15.445000  87.150000 16.245000  87.950000 ;
      RECT 15.445000  88.830000 16.245000  89.630000 ;
      RECT 15.445000  90.510000 16.245000  91.310000 ;
      RECT 15.445000  92.190000 16.245000  92.990000 ;
      RECT 15.445000  93.870000 16.245000  94.670000 ;
      RECT 15.445000 176.155000 16.245000 176.955000 ;
      RECT 15.445000 177.775000 16.245000 178.575000 ;
      RECT 15.445000 179.395000 16.245000 180.195000 ;
      RECT 15.445000 181.015000 16.245000 181.815000 ;
      RECT 15.445000 182.635000 16.245000 183.435000 ;
      RECT 15.445000 184.255000 16.245000 185.055000 ;
      RECT 15.445000 185.875000 16.245000 186.675000 ;
      RECT 15.445000 187.495000 16.245000 188.295000 ;
      RECT 15.445000 189.115000 16.245000 189.915000 ;
      RECT 15.445000 190.735000 16.245000 191.535000 ;
      RECT 15.445000 192.355000 16.245000 193.155000 ;
      RECT 15.445000 193.975000 16.245000 194.775000 ;
      RECT 15.445000 195.595000 16.245000 196.395000 ;
      RECT 15.445000 197.215000 16.245000 198.015000 ;
      RECT 15.445000 198.835000 16.245000 199.635000 ;
      RECT 15.450000   9.295000 16.250000  10.095000 ;
      RECT 15.450000  12.325000 16.250000  13.125000 ;
      RECT 17.045000  20.195000 17.845000  20.995000 ;
      RECT 17.045000  23.225000 17.845000  24.025000 ;
      RECT 17.045000  26.245000 17.845000  27.045000 ;
      RECT 17.045000  29.275000 17.845000  30.075000 ;
      RECT 17.050000   2.450000 17.850000   3.250000 ;
      RECT 17.050000   4.360000 17.850000   5.160000 ;
      RECT 17.050000   6.270000 17.850000   7.070000 ;
      RECT 17.050000  15.345000 17.850000  16.145000 ;
      RECT 17.050000  17.175000 17.850000  17.975000 ;
      RECT 17.050000  32.295000 17.850000  33.095000 ;
      RECT 17.050000  34.125000 17.850000  34.925000 ;
      RECT 17.050000  37.145000 17.850000  37.945000 ;
      RECT 17.050000  38.975000 17.850000  39.775000 ;
      RECT 17.050000  41.995000 17.850000  42.795000 ;
      RECT 17.050000  45.025000 17.850000  45.825000 ;
      RECT 17.050000  51.835000 17.850000  52.635000 ;
      RECT 17.050000  58.645000 17.850000  59.445000 ;
      RECT 17.050000  61.475000 17.850000  62.275000 ;
      RECT 17.050000  64.495000 17.850000  65.295000 ;
      RECT 17.050000  67.325000 17.850000  68.125000 ;
      RECT 17.050000  70.350000 17.850000  71.150000 ;
      RECT 17.050000  72.030000 17.850000  72.830000 ;
      RECT 17.050000  73.710000 17.850000  74.510000 ;
      RECT 17.050000  75.390000 17.850000  76.190000 ;
      RECT 17.050000  77.070000 17.850000  77.870000 ;
      RECT 17.050000  78.750000 17.850000  79.550000 ;
      RECT 17.050000  80.430000 17.850000  81.230000 ;
      RECT 17.050000  82.110000 17.850000  82.910000 ;
      RECT 17.050000  83.790000 17.850000  84.590000 ;
      RECT 17.050000  85.470000 17.850000  86.270000 ;
      RECT 17.050000  87.150000 17.850000  87.950000 ;
      RECT 17.050000  88.830000 17.850000  89.630000 ;
      RECT 17.050000  90.510000 17.850000  91.310000 ;
      RECT 17.050000  92.190000 17.850000  92.990000 ;
      RECT 17.050000  93.870000 17.850000  94.670000 ;
      RECT 17.050000 176.155000 17.850000 176.955000 ;
      RECT 17.050000 177.775000 17.850000 178.575000 ;
      RECT 17.050000 179.395000 17.850000 180.195000 ;
      RECT 17.050000 181.015000 17.850000 181.815000 ;
      RECT 17.050000 182.635000 17.850000 183.435000 ;
      RECT 17.050000 184.255000 17.850000 185.055000 ;
      RECT 17.050000 185.875000 17.850000 186.675000 ;
      RECT 17.050000 187.495000 17.850000 188.295000 ;
      RECT 17.050000 189.115000 17.850000 189.915000 ;
      RECT 17.050000 190.735000 17.850000 191.535000 ;
      RECT 17.050000 192.355000 17.850000 193.155000 ;
      RECT 17.050000 193.975000 17.850000 194.775000 ;
      RECT 17.050000 195.595000 17.850000 196.395000 ;
      RECT 17.050000 197.215000 17.850000 198.015000 ;
      RECT 17.050000 198.835000 17.850000 199.635000 ;
      RECT 17.055000   9.295000 17.855000  10.095000 ;
      RECT 17.055000  12.325000 17.855000  13.125000 ;
      RECT 18.650000  20.195000 19.450000  20.995000 ;
      RECT 18.650000  23.225000 19.450000  24.025000 ;
      RECT 18.650000  26.245000 19.450000  27.045000 ;
      RECT 18.650000  29.275000 19.450000  30.075000 ;
      RECT 18.655000   2.450000 19.455000   3.250000 ;
      RECT 18.655000   4.360000 19.455000   5.160000 ;
      RECT 18.655000   6.270000 19.455000   7.070000 ;
      RECT 18.655000  15.345000 19.455000  16.145000 ;
      RECT 18.655000  17.175000 19.455000  17.975000 ;
      RECT 18.655000  32.295000 19.455000  33.095000 ;
      RECT 18.655000  34.125000 19.455000  34.925000 ;
      RECT 18.655000  37.145000 19.455000  37.945000 ;
      RECT 18.655000  38.975000 19.455000  39.775000 ;
      RECT 18.655000  41.995000 19.455000  42.795000 ;
      RECT 18.655000  45.025000 19.455000  45.825000 ;
      RECT 18.655000  51.835000 19.455000  52.635000 ;
      RECT 18.655000  58.645000 19.455000  59.445000 ;
      RECT 18.655000  61.475000 19.455000  62.275000 ;
      RECT 18.655000  64.495000 19.455000  65.295000 ;
      RECT 18.655000  67.325000 19.455000  68.125000 ;
      RECT 18.655000  70.350000 19.455000  71.150000 ;
      RECT 18.655000  72.030000 19.455000  72.830000 ;
      RECT 18.655000  73.710000 19.455000  74.510000 ;
      RECT 18.655000  75.390000 19.455000  76.190000 ;
      RECT 18.655000  77.070000 19.455000  77.870000 ;
      RECT 18.655000  78.750000 19.455000  79.550000 ;
      RECT 18.655000  80.430000 19.455000  81.230000 ;
      RECT 18.655000  82.110000 19.455000  82.910000 ;
      RECT 18.655000  83.790000 19.455000  84.590000 ;
      RECT 18.655000  85.470000 19.455000  86.270000 ;
      RECT 18.655000  87.150000 19.455000  87.950000 ;
      RECT 18.655000  88.830000 19.455000  89.630000 ;
      RECT 18.655000  90.510000 19.455000  91.310000 ;
      RECT 18.655000  92.190000 19.455000  92.990000 ;
      RECT 18.655000  93.870000 19.455000  94.670000 ;
      RECT 18.655000 176.155000 19.455000 176.955000 ;
      RECT 18.655000 177.775000 19.455000 178.575000 ;
      RECT 18.655000 179.395000 19.455000 180.195000 ;
      RECT 18.655000 181.015000 19.455000 181.815000 ;
      RECT 18.655000 182.635000 19.455000 183.435000 ;
      RECT 18.655000 184.255000 19.455000 185.055000 ;
      RECT 18.655000 185.875000 19.455000 186.675000 ;
      RECT 18.655000 187.495000 19.455000 188.295000 ;
      RECT 18.655000 189.115000 19.455000 189.915000 ;
      RECT 18.655000 190.735000 19.455000 191.535000 ;
      RECT 18.655000 192.355000 19.455000 193.155000 ;
      RECT 18.655000 193.975000 19.455000 194.775000 ;
      RECT 18.655000 195.595000 19.455000 196.395000 ;
      RECT 18.655000 197.215000 19.455000 198.015000 ;
      RECT 18.655000 198.835000 19.455000 199.635000 ;
      RECT 18.660000   9.295000 19.460000  10.095000 ;
      RECT 18.660000  12.325000 19.460000  13.125000 ;
      RECT 20.255000  20.195000 21.055000  20.995000 ;
      RECT 20.255000  23.225000 21.055000  24.025000 ;
      RECT 20.255000  26.245000 21.055000  27.045000 ;
      RECT 20.255000  29.275000 21.055000  30.075000 ;
      RECT 20.260000   2.450000 21.060000   3.250000 ;
      RECT 20.260000   4.360000 21.060000   5.160000 ;
      RECT 20.260000   6.270000 21.060000   7.070000 ;
      RECT 20.260000  15.345000 21.060000  16.145000 ;
      RECT 20.260000  17.175000 21.060000  17.975000 ;
      RECT 20.260000  32.295000 21.060000  33.095000 ;
      RECT 20.260000  34.125000 21.060000  34.925000 ;
      RECT 20.260000  37.145000 21.060000  37.945000 ;
      RECT 20.260000  38.975000 21.060000  39.775000 ;
      RECT 20.260000  41.995000 21.060000  42.795000 ;
      RECT 20.260000  45.025000 21.060000  45.825000 ;
      RECT 20.260000  51.835000 21.060000  52.635000 ;
      RECT 20.260000  58.645000 21.060000  59.445000 ;
      RECT 20.260000  61.475000 21.060000  62.275000 ;
      RECT 20.260000  64.495000 21.060000  65.295000 ;
      RECT 20.260000  67.325000 21.060000  68.125000 ;
      RECT 20.260000  70.350000 21.060000  71.150000 ;
      RECT 20.260000  72.030000 21.060000  72.830000 ;
      RECT 20.260000  73.710000 21.060000  74.510000 ;
      RECT 20.260000  75.390000 21.060000  76.190000 ;
      RECT 20.260000  77.070000 21.060000  77.870000 ;
      RECT 20.260000  78.750000 21.060000  79.550000 ;
      RECT 20.260000  80.430000 21.060000  81.230000 ;
      RECT 20.260000  82.110000 21.060000  82.910000 ;
      RECT 20.260000  83.790000 21.060000  84.590000 ;
      RECT 20.260000  85.470000 21.060000  86.270000 ;
      RECT 20.260000  87.150000 21.060000  87.950000 ;
      RECT 20.260000  88.830000 21.060000  89.630000 ;
      RECT 20.260000  90.510000 21.060000  91.310000 ;
      RECT 20.260000  92.190000 21.060000  92.990000 ;
      RECT 20.260000  93.870000 21.060000  94.670000 ;
      RECT 20.260000 176.155000 21.060000 176.955000 ;
      RECT 20.260000 177.775000 21.060000 178.575000 ;
      RECT 20.260000 179.395000 21.060000 180.195000 ;
      RECT 20.260000 181.015000 21.060000 181.815000 ;
      RECT 20.260000 182.635000 21.060000 183.435000 ;
      RECT 20.260000 184.255000 21.060000 185.055000 ;
      RECT 20.260000 185.875000 21.060000 186.675000 ;
      RECT 20.260000 187.495000 21.060000 188.295000 ;
      RECT 20.260000 189.115000 21.060000 189.915000 ;
      RECT 20.260000 190.735000 21.060000 191.535000 ;
      RECT 20.260000 192.355000 21.060000 193.155000 ;
      RECT 20.260000 193.975000 21.060000 194.775000 ;
      RECT 20.260000 195.595000 21.060000 196.395000 ;
      RECT 20.260000 197.215000 21.060000 198.015000 ;
      RECT 20.260000 198.835000 21.060000 199.635000 ;
      RECT 20.265000   9.295000 21.065000  10.095000 ;
      RECT 20.265000  12.325000 21.065000  13.125000 ;
      RECT 21.860000  20.195000 22.660000  20.995000 ;
      RECT 21.860000  23.225000 22.660000  24.025000 ;
      RECT 21.860000  26.245000 22.660000  27.045000 ;
      RECT 21.860000  29.275000 22.660000  30.075000 ;
      RECT 21.865000   2.450000 22.665000   3.250000 ;
      RECT 21.865000   4.360000 22.665000   5.160000 ;
      RECT 21.865000   6.270000 22.665000   7.070000 ;
      RECT 21.865000  15.345000 22.665000  16.145000 ;
      RECT 21.865000  17.175000 22.665000  17.975000 ;
      RECT 21.865000  32.295000 22.665000  33.095000 ;
      RECT 21.865000  34.125000 22.665000  34.925000 ;
      RECT 21.865000  37.145000 22.665000  37.945000 ;
      RECT 21.865000  38.975000 22.665000  39.775000 ;
      RECT 21.865000  41.995000 22.665000  42.795000 ;
      RECT 21.865000  45.025000 22.665000  45.825000 ;
      RECT 21.865000  51.835000 22.665000  52.635000 ;
      RECT 21.865000  58.645000 22.665000  59.445000 ;
      RECT 21.865000  61.475000 22.665000  62.275000 ;
      RECT 21.865000  64.495000 22.665000  65.295000 ;
      RECT 21.865000  67.325000 22.665000  68.125000 ;
      RECT 21.865000  70.350000 22.665000  71.150000 ;
      RECT 21.865000  72.030000 22.665000  72.830000 ;
      RECT 21.865000  73.710000 22.665000  74.510000 ;
      RECT 21.865000  75.390000 22.665000  76.190000 ;
      RECT 21.865000  77.070000 22.665000  77.870000 ;
      RECT 21.865000  78.750000 22.665000  79.550000 ;
      RECT 21.865000  80.430000 22.665000  81.230000 ;
      RECT 21.865000  82.110000 22.665000  82.910000 ;
      RECT 21.865000  83.790000 22.665000  84.590000 ;
      RECT 21.865000  85.470000 22.665000  86.270000 ;
      RECT 21.865000  87.150000 22.665000  87.950000 ;
      RECT 21.865000  88.830000 22.665000  89.630000 ;
      RECT 21.865000  90.510000 22.665000  91.310000 ;
      RECT 21.865000  92.190000 22.665000  92.990000 ;
      RECT 21.865000  93.870000 22.665000  94.670000 ;
      RECT 21.865000 176.155000 22.665000 176.955000 ;
      RECT 21.865000 177.775000 22.665000 178.575000 ;
      RECT 21.865000 179.395000 22.665000 180.195000 ;
      RECT 21.865000 181.015000 22.665000 181.815000 ;
      RECT 21.865000 182.635000 22.665000 183.435000 ;
      RECT 21.865000 184.255000 22.665000 185.055000 ;
      RECT 21.865000 185.875000 22.665000 186.675000 ;
      RECT 21.865000 187.495000 22.665000 188.295000 ;
      RECT 21.865000 189.115000 22.665000 189.915000 ;
      RECT 21.865000 190.735000 22.665000 191.535000 ;
      RECT 21.865000 192.355000 22.665000 193.155000 ;
      RECT 21.865000 193.975000 22.665000 194.775000 ;
      RECT 21.865000 195.595000 22.665000 196.395000 ;
      RECT 21.865000 197.215000 22.665000 198.015000 ;
      RECT 21.865000 198.835000 22.665000 199.635000 ;
      RECT 21.870000   9.295000 22.670000  10.095000 ;
      RECT 21.870000  12.325000 22.670000  13.125000 ;
      RECT 23.465000  20.195000 24.265000  20.995000 ;
      RECT 23.465000  23.225000 24.265000  24.025000 ;
      RECT 23.465000  26.245000 24.265000  27.045000 ;
      RECT 23.465000  29.275000 24.265000  30.075000 ;
      RECT 23.470000   2.450000 24.270000   3.250000 ;
      RECT 23.470000   4.360000 24.270000   5.160000 ;
      RECT 23.470000   6.270000 24.270000   7.070000 ;
      RECT 23.470000  15.345000 24.270000  16.145000 ;
      RECT 23.470000  17.175000 24.270000  17.975000 ;
      RECT 23.470000  32.295000 24.270000  33.095000 ;
      RECT 23.470000  34.125000 24.270000  34.925000 ;
      RECT 23.470000  37.145000 24.270000  37.945000 ;
      RECT 23.470000  38.975000 24.270000  39.775000 ;
      RECT 23.470000  41.995000 24.270000  42.795000 ;
      RECT 23.470000  45.025000 24.270000  45.825000 ;
      RECT 23.470000  51.835000 24.270000  52.635000 ;
      RECT 23.470000  58.645000 24.270000  59.445000 ;
      RECT 23.470000  61.475000 24.270000  62.275000 ;
      RECT 23.470000  64.495000 24.270000  65.295000 ;
      RECT 23.470000  67.325000 24.270000  68.125000 ;
      RECT 23.470000  70.350000 24.270000  71.150000 ;
      RECT 23.470000  72.030000 24.270000  72.830000 ;
      RECT 23.470000  73.710000 24.270000  74.510000 ;
      RECT 23.470000  75.390000 24.270000  76.190000 ;
      RECT 23.470000  77.070000 24.270000  77.870000 ;
      RECT 23.470000  78.750000 24.270000  79.550000 ;
      RECT 23.470000  80.430000 24.270000  81.230000 ;
      RECT 23.470000  82.110000 24.270000  82.910000 ;
      RECT 23.470000  83.790000 24.270000  84.590000 ;
      RECT 23.470000  85.470000 24.270000  86.270000 ;
      RECT 23.470000  87.150000 24.270000  87.950000 ;
      RECT 23.470000  88.830000 24.270000  89.630000 ;
      RECT 23.470000  90.510000 24.270000  91.310000 ;
      RECT 23.470000  92.190000 24.270000  92.990000 ;
      RECT 23.470000  93.870000 24.270000  94.670000 ;
      RECT 23.470000 176.155000 24.270000 176.955000 ;
      RECT 23.470000 177.775000 24.270000 178.575000 ;
      RECT 23.470000 179.395000 24.270000 180.195000 ;
      RECT 23.470000 181.015000 24.270000 181.815000 ;
      RECT 23.470000 182.635000 24.270000 183.435000 ;
      RECT 23.470000 184.255000 24.270000 185.055000 ;
      RECT 23.470000 185.875000 24.270000 186.675000 ;
      RECT 23.470000 187.495000 24.270000 188.295000 ;
      RECT 23.470000 189.115000 24.270000 189.915000 ;
      RECT 23.470000 190.735000 24.270000 191.535000 ;
      RECT 23.470000 192.355000 24.270000 193.155000 ;
      RECT 23.470000 193.975000 24.270000 194.775000 ;
      RECT 23.470000 195.595000 24.270000 196.395000 ;
      RECT 23.470000 197.215000 24.270000 198.015000 ;
      RECT 23.470000 198.835000 24.270000 199.635000 ;
      RECT 23.475000   9.295000 24.275000  10.095000 ;
      RECT 23.475000  12.325000 24.275000  13.125000 ;
      RECT 25.070000  20.195000 25.870000  20.995000 ;
      RECT 25.070000  23.225000 25.870000  24.025000 ;
      RECT 25.070000  26.245000 25.870000  27.045000 ;
      RECT 25.070000  29.275000 25.870000  30.075000 ;
      RECT 25.075000   2.450000 25.875000   3.250000 ;
      RECT 25.075000   4.360000 25.875000   5.160000 ;
      RECT 25.075000   6.270000 25.875000   7.070000 ;
      RECT 25.075000  15.345000 25.875000  16.145000 ;
      RECT 25.075000  17.175000 25.875000  17.975000 ;
      RECT 25.075000  32.295000 25.875000  33.095000 ;
      RECT 25.075000  34.125000 25.875000  34.925000 ;
      RECT 25.075000  37.145000 25.875000  37.945000 ;
      RECT 25.075000  38.975000 25.875000  39.775000 ;
      RECT 25.075000  41.995000 25.875000  42.795000 ;
      RECT 25.075000  45.025000 25.875000  45.825000 ;
      RECT 25.075000  51.835000 25.875000  52.635000 ;
      RECT 25.075000  58.645000 25.875000  59.445000 ;
      RECT 25.075000  61.475000 25.875000  62.275000 ;
      RECT 25.075000  64.495000 25.875000  65.295000 ;
      RECT 25.075000  67.325000 25.875000  68.125000 ;
      RECT 25.075000  70.350000 25.875000  71.150000 ;
      RECT 25.075000  72.030000 25.875000  72.830000 ;
      RECT 25.075000  73.710000 25.875000  74.510000 ;
      RECT 25.075000  75.390000 25.875000  76.190000 ;
      RECT 25.075000  77.070000 25.875000  77.870000 ;
      RECT 25.075000  78.750000 25.875000  79.550000 ;
      RECT 25.075000  80.430000 25.875000  81.230000 ;
      RECT 25.075000  82.110000 25.875000  82.910000 ;
      RECT 25.075000  83.790000 25.875000  84.590000 ;
      RECT 25.075000  85.470000 25.875000  86.270000 ;
      RECT 25.075000  87.150000 25.875000  87.950000 ;
      RECT 25.075000  88.830000 25.875000  89.630000 ;
      RECT 25.075000  90.510000 25.875000  91.310000 ;
      RECT 25.075000  92.190000 25.875000  92.990000 ;
      RECT 25.075000  93.870000 25.875000  94.670000 ;
      RECT 25.075000 176.155000 25.875000 176.955000 ;
      RECT 25.075000 177.775000 25.875000 178.575000 ;
      RECT 25.075000 179.395000 25.875000 180.195000 ;
      RECT 25.075000 181.015000 25.875000 181.815000 ;
      RECT 25.075000 182.635000 25.875000 183.435000 ;
      RECT 25.075000 184.255000 25.875000 185.055000 ;
      RECT 25.075000 185.875000 25.875000 186.675000 ;
      RECT 25.075000 187.495000 25.875000 188.295000 ;
      RECT 25.075000 189.115000 25.875000 189.915000 ;
      RECT 25.075000 190.735000 25.875000 191.535000 ;
      RECT 25.075000 192.355000 25.875000 193.155000 ;
      RECT 25.075000 193.975000 25.875000 194.775000 ;
      RECT 25.075000 195.595000 25.875000 196.395000 ;
      RECT 25.075000 197.215000 25.875000 198.015000 ;
      RECT 25.075000 198.835000 25.875000 199.635000 ;
      RECT 25.080000   9.295000 25.880000  10.095000 ;
      RECT 25.080000  12.325000 25.880000  13.125000 ;
      RECT 26.675000  20.195000 27.475000  20.995000 ;
      RECT 26.675000  23.225000 27.475000  24.025000 ;
      RECT 26.675000  26.245000 27.475000  27.045000 ;
      RECT 26.675000  29.275000 27.475000  30.075000 ;
      RECT 26.680000   2.450000 27.480000   3.250000 ;
      RECT 26.680000   4.360000 27.480000   5.160000 ;
      RECT 26.680000   6.270000 27.480000   7.070000 ;
      RECT 26.680000  15.345000 27.480000  16.145000 ;
      RECT 26.680000  17.175000 27.480000  17.975000 ;
      RECT 26.680000  32.295000 27.480000  33.095000 ;
      RECT 26.680000  34.125000 27.480000  34.925000 ;
      RECT 26.680000  37.145000 27.480000  37.945000 ;
      RECT 26.680000  38.975000 27.480000  39.775000 ;
      RECT 26.680000  41.995000 27.480000  42.795000 ;
      RECT 26.680000  45.025000 27.480000  45.825000 ;
      RECT 26.680000  51.835000 27.480000  52.635000 ;
      RECT 26.680000  58.645000 27.480000  59.445000 ;
      RECT 26.680000  61.475000 27.480000  62.275000 ;
      RECT 26.680000  64.495000 27.480000  65.295000 ;
      RECT 26.680000  67.325000 27.480000  68.125000 ;
      RECT 26.680000  70.350000 27.480000  71.150000 ;
      RECT 26.680000  72.030000 27.480000  72.830000 ;
      RECT 26.680000  73.710000 27.480000  74.510000 ;
      RECT 26.680000  75.390000 27.480000  76.190000 ;
      RECT 26.680000  77.070000 27.480000  77.870000 ;
      RECT 26.680000  78.750000 27.480000  79.550000 ;
      RECT 26.680000  80.430000 27.480000  81.230000 ;
      RECT 26.680000  82.110000 27.480000  82.910000 ;
      RECT 26.680000  83.790000 27.480000  84.590000 ;
      RECT 26.680000  85.470000 27.480000  86.270000 ;
      RECT 26.680000  87.150000 27.480000  87.950000 ;
      RECT 26.680000  88.830000 27.480000  89.630000 ;
      RECT 26.680000  90.510000 27.480000  91.310000 ;
      RECT 26.680000  92.190000 27.480000  92.990000 ;
      RECT 26.680000  93.870000 27.480000  94.670000 ;
      RECT 26.680000 176.155000 27.480000 176.955000 ;
      RECT 26.680000 177.775000 27.480000 178.575000 ;
      RECT 26.680000 179.395000 27.480000 180.195000 ;
      RECT 26.680000 181.015000 27.480000 181.815000 ;
      RECT 26.680000 182.635000 27.480000 183.435000 ;
      RECT 26.680000 184.255000 27.480000 185.055000 ;
      RECT 26.680000 185.875000 27.480000 186.675000 ;
      RECT 26.680000 187.495000 27.480000 188.295000 ;
      RECT 26.680000 189.115000 27.480000 189.915000 ;
      RECT 26.680000 190.735000 27.480000 191.535000 ;
      RECT 26.680000 192.355000 27.480000 193.155000 ;
      RECT 26.680000 193.975000 27.480000 194.775000 ;
      RECT 26.680000 195.595000 27.480000 196.395000 ;
      RECT 26.680000 197.215000 27.480000 198.015000 ;
      RECT 26.680000 198.835000 27.480000 199.635000 ;
      RECT 26.685000   9.295000 27.485000  10.095000 ;
      RECT 26.685000  12.325000 27.485000  13.125000 ;
      RECT 28.280000  20.195000 29.080000  20.995000 ;
      RECT 28.280000  23.225000 29.080000  24.025000 ;
      RECT 28.280000  26.245000 29.080000  27.045000 ;
      RECT 28.280000  29.275000 29.080000  30.075000 ;
      RECT 28.285000   2.450000 29.085000   3.250000 ;
      RECT 28.285000   4.360000 29.085000   5.160000 ;
      RECT 28.285000   6.270000 29.085000   7.070000 ;
      RECT 28.285000  15.345000 29.085000  16.145000 ;
      RECT 28.285000  17.175000 29.085000  17.975000 ;
      RECT 28.285000  32.295000 29.085000  33.095000 ;
      RECT 28.285000  34.125000 29.085000  34.925000 ;
      RECT 28.285000  37.145000 29.085000  37.945000 ;
      RECT 28.285000  38.975000 29.085000  39.775000 ;
      RECT 28.285000  41.995000 29.085000  42.795000 ;
      RECT 28.285000  45.025000 29.085000  45.825000 ;
      RECT 28.285000  51.835000 29.085000  52.635000 ;
      RECT 28.285000  58.645000 29.085000  59.445000 ;
      RECT 28.285000  61.475000 29.085000  62.275000 ;
      RECT 28.285000  64.495000 29.085000  65.295000 ;
      RECT 28.285000  67.325000 29.085000  68.125000 ;
      RECT 28.285000  70.350000 29.085000  71.150000 ;
      RECT 28.285000  72.030000 29.085000  72.830000 ;
      RECT 28.285000  73.710000 29.085000  74.510000 ;
      RECT 28.285000  75.390000 29.085000  76.190000 ;
      RECT 28.285000  77.070000 29.085000  77.870000 ;
      RECT 28.285000  78.750000 29.085000  79.550000 ;
      RECT 28.285000  80.430000 29.085000  81.230000 ;
      RECT 28.285000  82.110000 29.085000  82.910000 ;
      RECT 28.285000  83.790000 29.085000  84.590000 ;
      RECT 28.285000  85.470000 29.085000  86.270000 ;
      RECT 28.285000  87.150000 29.085000  87.950000 ;
      RECT 28.285000  88.830000 29.085000  89.630000 ;
      RECT 28.285000  90.510000 29.085000  91.310000 ;
      RECT 28.285000  92.190000 29.085000  92.990000 ;
      RECT 28.285000  93.870000 29.085000  94.670000 ;
      RECT 28.285000 176.155000 29.085000 176.955000 ;
      RECT 28.285000 177.775000 29.085000 178.575000 ;
      RECT 28.285000 179.395000 29.085000 180.195000 ;
      RECT 28.285000 181.015000 29.085000 181.815000 ;
      RECT 28.285000 182.635000 29.085000 183.435000 ;
      RECT 28.285000 184.255000 29.085000 185.055000 ;
      RECT 28.285000 185.875000 29.085000 186.675000 ;
      RECT 28.285000 187.495000 29.085000 188.295000 ;
      RECT 28.285000 189.115000 29.085000 189.915000 ;
      RECT 28.285000 190.735000 29.085000 191.535000 ;
      RECT 28.285000 192.355000 29.085000 193.155000 ;
      RECT 28.285000 193.975000 29.085000 194.775000 ;
      RECT 28.285000 195.595000 29.085000 196.395000 ;
      RECT 28.285000 197.215000 29.085000 198.015000 ;
      RECT 28.285000 198.835000 29.085000 199.635000 ;
      RECT 28.290000   9.295000 29.090000  10.095000 ;
      RECT 28.290000  12.325000 29.090000  13.125000 ;
      RECT 29.885000  20.195000 30.685000  20.995000 ;
      RECT 29.885000  23.225000 30.685000  24.025000 ;
      RECT 29.885000  26.245000 30.685000  27.045000 ;
      RECT 29.885000  29.275000 30.685000  30.075000 ;
      RECT 29.890000   2.450000 30.690000   3.250000 ;
      RECT 29.890000   4.360000 30.690000   5.160000 ;
      RECT 29.890000   6.270000 30.690000   7.070000 ;
      RECT 29.890000  15.345000 30.690000  16.145000 ;
      RECT 29.890000  17.175000 30.690000  17.975000 ;
      RECT 29.890000  32.295000 30.690000  33.095000 ;
      RECT 29.890000  34.125000 30.690000  34.925000 ;
      RECT 29.890000  37.145000 30.690000  37.945000 ;
      RECT 29.890000  38.975000 30.690000  39.775000 ;
      RECT 29.890000  41.995000 30.690000  42.795000 ;
      RECT 29.890000  45.025000 30.690000  45.825000 ;
      RECT 29.890000  51.835000 30.690000  52.635000 ;
      RECT 29.890000  58.645000 30.690000  59.445000 ;
      RECT 29.890000  61.475000 30.690000  62.275000 ;
      RECT 29.890000  64.495000 30.690000  65.295000 ;
      RECT 29.890000  67.325000 30.690000  68.125000 ;
      RECT 29.890000  70.350000 30.690000  71.150000 ;
      RECT 29.890000  72.030000 30.690000  72.830000 ;
      RECT 29.890000  73.710000 30.690000  74.510000 ;
      RECT 29.890000  75.390000 30.690000  76.190000 ;
      RECT 29.890000  77.070000 30.690000  77.870000 ;
      RECT 29.890000  78.750000 30.690000  79.550000 ;
      RECT 29.890000  80.430000 30.690000  81.230000 ;
      RECT 29.890000  82.110000 30.690000  82.910000 ;
      RECT 29.890000  83.790000 30.690000  84.590000 ;
      RECT 29.890000  85.470000 30.690000  86.270000 ;
      RECT 29.890000  87.150000 30.690000  87.950000 ;
      RECT 29.890000  88.830000 30.690000  89.630000 ;
      RECT 29.890000  90.510000 30.690000  91.310000 ;
      RECT 29.890000  92.190000 30.690000  92.990000 ;
      RECT 29.890000  93.870000 30.690000  94.670000 ;
      RECT 29.890000 176.155000 30.690000 176.955000 ;
      RECT 29.890000 177.775000 30.690000 178.575000 ;
      RECT 29.890000 179.395000 30.690000 180.195000 ;
      RECT 29.890000 181.015000 30.690000 181.815000 ;
      RECT 29.890000 182.635000 30.690000 183.435000 ;
      RECT 29.890000 184.255000 30.690000 185.055000 ;
      RECT 29.890000 185.875000 30.690000 186.675000 ;
      RECT 29.890000 187.495000 30.690000 188.295000 ;
      RECT 29.890000 189.115000 30.690000 189.915000 ;
      RECT 29.890000 190.735000 30.690000 191.535000 ;
      RECT 29.890000 192.355000 30.690000 193.155000 ;
      RECT 29.890000 193.975000 30.690000 194.775000 ;
      RECT 29.890000 195.595000 30.690000 196.395000 ;
      RECT 29.890000 197.215000 30.690000 198.015000 ;
      RECT 29.890000 198.835000 30.690000 199.635000 ;
      RECT 29.895000   9.295000 30.695000  10.095000 ;
      RECT 29.895000  12.325000 30.695000  13.125000 ;
      RECT 31.490000  20.195000 32.290000  20.995000 ;
      RECT 31.490000  23.225000 32.290000  24.025000 ;
      RECT 31.490000  26.245000 32.290000  27.045000 ;
      RECT 31.490000  29.275000 32.290000  30.075000 ;
      RECT 31.495000   2.450000 32.295000   3.250000 ;
      RECT 31.495000   4.360000 32.295000   5.160000 ;
      RECT 31.495000   6.270000 32.295000   7.070000 ;
      RECT 31.495000  15.345000 32.295000  16.145000 ;
      RECT 31.495000  17.175000 32.295000  17.975000 ;
      RECT 31.495000  32.295000 32.295000  33.095000 ;
      RECT 31.495000  34.125000 32.295000  34.925000 ;
      RECT 31.495000  37.145000 32.295000  37.945000 ;
      RECT 31.495000  38.975000 32.295000  39.775000 ;
      RECT 31.495000  41.995000 32.295000  42.795000 ;
      RECT 31.495000  45.025000 32.295000  45.825000 ;
      RECT 31.495000  51.835000 32.295000  52.635000 ;
      RECT 31.495000  58.645000 32.295000  59.445000 ;
      RECT 31.495000  61.475000 32.295000  62.275000 ;
      RECT 31.495000  64.495000 32.295000  65.295000 ;
      RECT 31.495000  67.325000 32.295000  68.125000 ;
      RECT 31.495000  70.350000 32.295000  71.150000 ;
      RECT 31.495000  72.030000 32.295000  72.830000 ;
      RECT 31.495000  73.710000 32.295000  74.510000 ;
      RECT 31.495000  75.390000 32.295000  76.190000 ;
      RECT 31.495000  77.070000 32.295000  77.870000 ;
      RECT 31.495000  78.750000 32.295000  79.550000 ;
      RECT 31.495000  80.430000 32.295000  81.230000 ;
      RECT 31.495000  82.110000 32.295000  82.910000 ;
      RECT 31.495000  83.790000 32.295000  84.590000 ;
      RECT 31.495000  85.470000 32.295000  86.270000 ;
      RECT 31.495000  87.150000 32.295000  87.950000 ;
      RECT 31.495000  88.830000 32.295000  89.630000 ;
      RECT 31.495000  90.510000 32.295000  91.310000 ;
      RECT 31.495000  92.190000 32.295000  92.990000 ;
      RECT 31.495000  93.870000 32.295000  94.670000 ;
      RECT 31.495000 176.155000 32.295000 176.955000 ;
      RECT 31.495000 177.775000 32.295000 178.575000 ;
      RECT 31.495000 179.395000 32.295000 180.195000 ;
      RECT 31.495000 181.015000 32.295000 181.815000 ;
      RECT 31.495000 182.635000 32.295000 183.435000 ;
      RECT 31.495000 184.255000 32.295000 185.055000 ;
      RECT 31.495000 185.875000 32.295000 186.675000 ;
      RECT 31.495000 187.495000 32.295000 188.295000 ;
      RECT 31.495000 189.115000 32.295000 189.915000 ;
      RECT 31.495000 190.735000 32.295000 191.535000 ;
      RECT 31.495000 192.355000 32.295000 193.155000 ;
      RECT 31.495000 193.975000 32.295000 194.775000 ;
      RECT 31.495000 195.595000 32.295000 196.395000 ;
      RECT 31.495000 197.215000 32.295000 198.015000 ;
      RECT 31.495000 198.835000 32.295000 199.635000 ;
      RECT 31.500000   9.295000 32.300000  10.095000 ;
      RECT 31.500000  12.325000 32.300000  13.125000 ;
      RECT 33.095000  20.195000 33.895000  20.995000 ;
      RECT 33.095000  23.225000 33.895000  24.025000 ;
      RECT 33.095000  26.245000 33.895000  27.045000 ;
      RECT 33.095000  29.275000 33.895000  30.075000 ;
      RECT 33.100000   2.450000 33.900000   3.250000 ;
      RECT 33.100000   4.360000 33.900000   5.160000 ;
      RECT 33.100000   6.270000 33.900000   7.070000 ;
      RECT 33.100000  15.345000 33.900000  16.145000 ;
      RECT 33.100000  17.175000 33.900000  17.975000 ;
      RECT 33.100000  32.295000 33.900000  33.095000 ;
      RECT 33.100000  34.125000 33.900000  34.925000 ;
      RECT 33.100000  37.145000 33.900000  37.945000 ;
      RECT 33.100000  38.975000 33.900000  39.775000 ;
      RECT 33.100000  41.995000 33.900000  42.795000 ;
      RECT 33.100000  45.025000 33.900000  45.825000 ;
      RECT 33.100000  51.835000 33.900000  52.635000 ;
      RECT 33.100000  58.645000 33.900000  59.445000 ;
      RECT 33.100000  61.475000 33.900000  62.275000 ;
      RECT 33.100000  64.495000 33.900000  65.295000 ;
      RECT 33.100000  67.325000 33.900000  68.125000 ;
      RECT 33.100000  70.350000 33.900000  71.150000 ;
      RECT 33.100000  72.030000 33.900000  72.830000 ;
      RECT 33.100000  73.710000 33.900000  74.510000 ;
      RECT 33.100000  75.390000 33.900000  76.190000 ;
      RECT 33.100000  77.070000 33.900000  77.870000 ;
      RECT 33.100000  78.750000 33.900000  79.550000 ;
      RECT 33.100000  80.430000 33.900000  81.230000 ;
      RECT 33.100000  82.110000 33.900000  82.910000 ;
      RECT 33.100000  83.790000 33.900000  84.590000 ;
      RECT 33.100000  85.470000 33.900000  86.270000 ;
      RECT 33.100000  87.150000 33.900000  87.950000 ;
      RECT 33.100000  88.830000 33.900000  89.630000 ;
      RECT 33.100000  90.510000 33.900000  91.310000 ;
      RECT 33.100000  92.190000 33.900000  92.990000 ;
      RECT 33.100000  93.870000 33.900000  94.670000 ;
      RECT 33.100000 176.155000 33.900000 176.955000 ;
      RECT 33.100000 177.775000 33.900000 178.575000 ;
      RECT 33.100000 179.395000 33.900000 180.195000 ;
      RECT 33.100000 181.015000 33.900000 181.815000 ;
      RECT 33.100000 182.635000 33.900000 183.435000 ;
      RECT 33.100000 184.255000 33.900000 185.055000 ;
      RECT 33.100000 185.875000 33.900000 186.675000 ;
      RECT 33.100000 187.495000 33.900000 188.295000 ;
      RECT 33.100000 189.115000 33.900000 189.915000 ;
      RECT 33.100000 190.735000 33.900000 191.535000 ;
      RECT 33.100000 192.355000 33.900000 193.155000 ;
      RECT 33.100000 193.975000 33.900000 194.775000 ;
      RECT 33.100000 195.595000 33.900000 196.395000 ;
      RECT 33.100000 197.215000 33.900000 198.015000 ;
      RECT 33.100000 198.835000 33.900000 199.635000 ;
      RECT 33.105000   9.295000 33.905000  10.095000 ;
      RECT 33.105000  12.325000 33.905000  13.125000 ;
      RECT 34.700000  20.195000 35.500000  20.995000 ;
      RECT 34.700000  23.225000 35.500000  24.025000 ;
      RECT 34.700000  26.245000 35.500000  27.045000 ;
      RECT 34.700000  29.275000 35.500000  30.075000 ;
      RECT 34.705000   2.450000 35.505000   3.250000 ;
      RECT 34.705000   4.360000 35.505000   5.160000 ;
      RECT 34.705000   6.270000 35.505000   7.070000 ;
      RECT 34.705000  15.345000 35.505000  16.145000 ;
      RECT 34.705000  17.175000 35.505000  17.975000 ;
      RECT 34.705000  32.295000 35.505000  33.095000 ;
      RECT 34.705000  34.125000 35.505000  34.925000 ;
      RECT 34.705000  37.145000 35.505000  37.945000 ;
      RECT 34.705000  38.975000 35.505000  39.775000 ;
      RECT 34.705000  41.995000 35.505000  42.795000 ;
      RECT 34.705000  45.025000 35.505000  45.825000 ;
      RECT 34.705000  51.835000 35.505000  52.635000 ;
      RECT 34.705000  58.645000 35.505000  59.445000 ;
      RECT 34.705000  61.475000 35.505000  62.275000 ;
      RECT 34.705000  64.495000 35.505000  65.295000 ;
      RECT 34.705000  67.325000 35.505000  68.125000 ;
      RECT 34.705000  70.350000 35.505000  71.150000 ;
      RECT 34.705000  72.030000 35.505000  72.830000 ;
      RECT 34.705000  73.710000 35.505000  74.510000 ;
      RECT 34.705000  75.390000 35.505000  76.190000 ;
      RECT 34.705000  77.070000 35.505000  77.870000 ;
      RECT 34.705000  78.750000 35.505000  79.550000 ;
      RECT 34.705000  80.430000 35.505000  81.230000 ;
      RECT 34.705000  82.110000 35.505000  82.910000 ;
      RECT 34.705000  83.790000 35.505000  84.590000 ;
      RECT 34.705000  85.470000 35.505000  86.270000 ;
      RECT 34.705000  87.150000 35.505000  87.950000 ;
      RECT 34.705000  88.830000 35.505000  89.630000 ;
      RECT 34.705000  90.510000 35.505000  91.310000 ;
      RECT 34.705000  92.190000 35.505000  92.990000 ;
      RECT 34.705000  93.870000 35.505000  94.670000 ;
      RECT 34.705000 176.155000 35.505000 176.955000 ;
      RECT 34.705000 177.775000 35.505000 178.575000 ;
      RECT 34.705000 179.395000 35.505000 180.195000 ;
      RECT 34.705000 181.015000 35.505000 181.815000 ;
      RECT 34.705000 182.635000 35.505000 183.435000 ;
      RECT 34.705000 184.255000 35.505000 185.055000 ;
      RECT 34.705000 185.875000 35.505000 186.675000 ;
      RECT 34.705000 187.495000 35.505000 188.295000 ;
      RECT 34.705000 189.115000 35.505000 189.915000 ;
      RECT 34.705000 190.735000 35.505000 191.535000 ;
      RECT 34.705000 192.355000 35.505000 193.155000 ;
      RECT 34.705000 193.975000 35.505000 194.775000 ;
      RECT 34.705000 195.595000 35.505000 196.395000 ;
      RECT 34.705000 197.215000 35.505000 198.015000 ;
      RECT 34.705000 198.835000 35.505000 199.635000 ;
      RECT 34.710000   9.295000 35.510000  10.095000 ;
      RECT 34.710000  12.325000 35.510000  13.125000 ;
      RECT 36.305000  20.195000 37.105000  20.995000 ;
      RECT 36.305000  23.225000 37.105000  24.025000 ;
      RECT 36.305000  26.245000 37.105000  27.045000 ;
      RECT 36.305000  29.275000 37.105000  30.075000 ;
      RECT 36.310000   2.450000 37.110000   3.250000 ;
      RECT 36.310000   4.360000 37.110000   5.160000 ;
      RECT 36.310000   6.270000 37.110000   7.070000 ;
      RECT 36.310000  15.345000 37.110000  16.145000 ;
      RECT 36.310000  17.175000 37.110000  17.975000 ;
      RECT 36.310000  32.295000 37.110000  33.095000 ;
      RECT 36.310000  34.125000 37.110000  34.925000 ;
      RECT 36.310000  37.145000 37.110000  37.945000 ;
      RECT 36.310000  38.975000 37.110000  39.775000 ;
      RECT 36.310000  41.995000 37.110000  42.795000 ;
      RECT 36.310000  45.025000 37.110000  45.825000 ;
      RECT 36.310000  51.835000 37.110000  52.635000 ;
      RECT 36.310000  58.645000 37.110000  59.445000 ;
      RECT 36.310000  61.475000 37.110000  62.275000 ;
      RECT 36.310000  64.495000 37.110000  65.295000 ;
      RECT 36.310000  67.325000 37.110000  68.125000 ;
      RECT 36.310000  70.350000 37.110000  71.150000 ;
      RECT 36.310000  72.030000 37.110000  72.830000 ;
      RECT 36.310000  73.710000 37.110000  74.510000 ;
      RECT 36.310000  75.390000 37.110000  76.190000 ;
      RECT 36.310000  77.070000 37.110000  77.870000 ;
      RECT 36.310000  78.750000 37.110000  79.550000 ;
      RECT 36.310000  80.430000 37.110000  81.230000 ;
      RECT 36.310000  82.110000 37.110000  82.910000 ;
      RECT 36.310000  83.790000 37.110000  84.590000 ;
      RECT 36.310000  85.470000 37.110000  86.270000 ;
      RECT 36.310000  87.150000 37.110000  87.950000 ;
      RECT 36.310000  88.830000 37.110000  89.630000 ;
      RECT 36.310000  90.510000 37.110000  91.310000 ;
      RECT 36.310000  92.190000 37.110000  92.990000 ;
      RECT 36.310000  93.870000 37.110000  94.670000 ;
      RECT 36.310000 176.155000 37.110000 176.955000 ;
      RECT 36.310000 177.775000 37.110000 178.575000 ;
      RECT 36.310000 179.395000 37.110000 180.195000 ;
      RECT 36.310000 181.015000 37.110000 181.815000 ;
      RECT 36.310000 182.635000 37.110000 183.435000 ;
      RECT 36.310000 184.255000 37.110000 185.055000 ;
      RECT 36.310000 185.875000 37.110000 186.675000 ;
      RECT 36.310000 187.495000 37.110000 188.295000 ;
      RECT 36.310000 189.115000 37.110000 189.915000 ;
      RECT 36.310000 190.735000 37.110000 191.535000 ;
      RECT 36.310000 192.355000 37.110000 193.155000 ;
      RECT 36.310000 193.975000 37.110000 194.775000 ;
      RECT 36.310000 195.595000 37.110000 196.395000 ;
      RECT 36.310000 197.215000 37.110000 198.015000 ;
      RECT 36.310000 198.835000 37.110000 199.635000 ;
      RECT 36.315000   9.295000 37.115000  10.095000 ;
      RECT 36.315000  12.325000 37.115000  13.125000 ;
      RECT 37.910000  20.195000 38.710000  20.995000 ;
      RECT 37.910000  23.225000 38.710000  24.025000 ;
      RECT 37.910000  26.245000 38.710000  27.045000 ;
      RECT 37.910000  29.275000 38.710000  30.075000 ;
      RECT 37.915000   2.450000 38.715000   3.250000 ;
      RECT 37.915000   4.360000 38.715000   5.160000 ;
      RECT 37.915000   6.270000 38.715000   7.070000 ;
      RECT 37.915000  15.345000 38.715000  16.145000 ;
      RECT 37.915000  17.175000 38.715000  17.975000 ;
      RECT 37.915000  32.295000 38.715000  33.095000 ;
      RECT 37.915000  34.125000 38.715000  34.925000 ;
      RECT 37.915000  37.145000 38.715000  37.945000 ;
      RECT 37.915000  38.975000 38.715000  39.775000 ;
      RECT 37.915000  41.995000 38.715000  42.795000 ;
      RECT 37.915000  45.025000 38.715000  45.825000 ;
      RECT 37.915000  51.835000 38.715000  52.635000 ;
      RECT 37.915000  58.645000 38.715000  59.445000 ;
      RECT 37.915000  61.475000 38.715000  62.275000 ;
      RECT 37.915000  64.495000 38.715000  65.295000 ;
      RECT 37.915000  67.325000 38.715000  68.125000 ;
      RECT 37.915000  70.350000 38.715000  71.150000 ;
      RECT 37.915000  72.030000 38.715000  72.830000 ;
      RECT 37.915000  73.710000 38.715000  74.510000 ;
      RECT 37.915000  75.390000 38.715000  76.190000 ;
      RECT 37.915000  77.070000 38.715000  77.870000 ;
      RECT 37.915000  78.750000 38.715000  79.550000 ;
      RECT 37.915000  80.430000 38.715000  81.230000 ;
      RECT 37.915000  82.110000 38.715000  82.910000 ;
      RECT 37.915000  83.790000 38.715000  84.590000 ;
      RECT 37.915000  85.470000 38.715000  86.270000 ;
      RECT 37.915000  87.150000 38.715000  87.950000 ;
      RECT 37.915000  88.830000 38.715000  89.630000 ;
      RECT 37.915000  90.510000 38.715000  91.310000 ;
      RECT 37.915000  92.190000 38.715000  92.990000 ;
      RECT 37.915000  93.870000 38.715000  94.670000 ;
      RECT 37.915000 176.155000 38.715000 176.955000 ;
      RECT 37.915000 177.775000 38.715000 178.575000 ;
      RECT 37.915000 179.395000 38.715000 180.195000 ;
      RECT 37.915000 181.015000 38.715000 181.815000 ;
      RECT 37.915000 182.635000 38.715000 183.435000 ;
      RECT 37.915000 184.255000 38.715000 185.055000 ;
      RECT 37.915000 185.875000 38.715000 186.675000 ;
      RECT 37.915000 187.495000 38.715000 188.295000 ;
      RECT 37.915000 189.115000 38.715000 189.915000 ;
      RECT 37.915000 190.735000 38.715000 191.535000 ;
      RECT 37.915000 192.355000 38.715000 193.155000 ;
      RECT 37.915000 193.975000 38.715000 194.775000 ;
      RECT 37.915000 195.595000 38.715000 196.395000 ;
      RECT 37.915000 197.215000 38.715000 198.015000 ;
      RECT 37.915000 198.835000 38.715000 199.635000 ;
      RECT 37.920000   9.295000 38.720000  10.095000 ;
      RECT 37.920000  12.325000 38.720000  13.125000 ;
      RECT 39.515000  20.195000 40.315000  20.995000 ;
      RECT 39.515000  23.225000 40.315000  24.025000 ;
      RECT 39.515000  26.245000 40.315000  27.045000 ;
      RECT 39.515000  29.275000 40.315000  30.075000 ;
      RECT 39.520000   2.450000 40.320000   3.250000 ;
      RECT 39.520000   4.360000 40.320000   5.160000 ;
      RECT 39.520000   6.270000 40.320000   7.070000 ;
      RECT 39.520000  15.345000 40.320000  16.145000 ;
      RECT 39.520000  17.175000 40.320000  17.975000 ;
      RECT 39.520000  32.295000 40.320000  33.095000 ;
      RECT 39.520000  34.125000 40.320000  34.925000 ;
      RECT 39.520000  37.145000 40.320000  37.945000 ;
      RECT 39.520000  38.975000 40.320000  39.775000 ;
      RECT 39.520000  41.995000 40.320000  42.795000 ;
      RECT 39.520000  45.025000 40.320000  45.825000 ;
      RECT 39.520000  51.835000 40.320000  52.635000 ;
      RECT 39.520000  58.645000 40.320000  59.445000 ;
      RECT 39.520000  61.475000 40.320000  62.275000 ;
      RECT 39.520000  64.495000 40.320000  65.295000 ;
      RECT 39.520000  67.325000 40.320000  68.125000 ;
      RECT 39.520000  70.350000 40.320000  71.150000 ;
      RECT 39.520000  72.030000 40.320000  72.830000 ;
      RECT 39.520000  73.710000 40.320000  74.510000 ;
      RECT 39.520000  75.390000 40.320000  76.190000 ;
      RECT 39.520000  77.070000 40.320000  77.870000 ;
      RECT 39.520000  78.750000 40.320000  79.550000 ;
      RECT 39.520000  80.430000 40.320000  81.230000 ;
      RECT 39.520000  82.110000 40.320000  82.910000 ;
      RECT 39.520000  83.790000 40.320000  84.590000 ;
      RECT 39.520000  85.470000 40.320000  86.270000 ;
      RECT 39.520000  87.150000 40.320000  87.950000 ;
      RECT 39.520000  88.830000 40.320000  89.630000 ;
      RECT 39.520000  90.510000 40.320000  91.310000 ;
      RECT 39.520000  92.190000 40.320000  92.990000 ;
      RECT 39.520000  93.870000 40.320000  94.670000 ;
      RECT 39.520000 176.155000 40.320000 176.955000 ;
      RECT 39.520000 177.775000 40.320000 178.575000 ;
      RECT 39.520000 179.395000 40.320000 180.195000 ;
      RECT 39.520000 181.015000 40.320000 181.815000 ;
      RECT 39.520000 182.635000 40.320000 183.435000 ;
      RECT 39.520000 184.255000 40.320000 185.055000 ;
      RECT 39.520000 185.875000 40.320000 186.675000 ;
      RECT 39.520000 187.495000 40.320000 188.295000 ;
      RECT 39.520000 189.115000 40.320000 189.915000 ;
      RECT 39.520000 190.735000 40.320000 191.535000 ;
      RECT 39.520000 192.355000 40.320000 193.155000 ;
      RECT 39.520000 193.975000 40.320000 194.775000 ;
      RECT 39.520000 195.595000 40.320000 196.395000 ;
      RECT 39.520000 197.215000 40.320000 198.015000 ;
      RECT 39.520000 198.835000 40.320000 199.635000 ;
      RECT 39.525000   9.295000 40.325000  10.095000 ;
      RECT 39.525000  12.325000 40.325000  13.125000 ;
      RECT 41.120000  20.195000 41.920000  20.995000 ;
      RECT 41.120000  23.225000 41.920000  24.025000 ;
      RECT 41.120000  26.245000 41.920000  27.045000 ;
      RECT 41.120000  29.275000 41.920000  30.075000 ;
      RECT 41.125000   2.450000 41.925000   3.250000 ;
      RECT 41.125000   4.360000 41.925000   5.160000 ;
      RECT 41.125000   6.270000 41.925000   7.070000 ;
      RECT 41.125000  15.345000 41.925000  16.145000 ;
      RECT 41.125000  17.175000 41.925000  17.975000 ;
      RECT 41.125000  32.295000 41.925000  33.095000 ;
      RECT 41.125000  34.125000 41.925000  34.925000 ;
      RECT 41.125000  37.145000 41.925000  37.945000 ;
      RECT 41.125000  38.975000 41.925000  39.775000 ;
      RECT 41.125000  41.995000 41.925000  42.795000 ;
      RECT 41.125000  45.025000 41.925000  45.825000 ;
      RECT 41.125000  51.835000 41.925000  52.635000 ;
      RECT 41.125000  58.645000 41.925000  59.445000 ;
      RECT 41.125000  61.475000 41.925000  62.275000 ;
      RECT 41.125000  64.495000 41.925000  65.295000 ;
      RECT 41.125000  67.325000 41.925000  68.125000 ;
      RECT 41.125000  70.350000 41.925000  71.150000 ;
      RECT 41.125000  72.030000 41.925000  72.830000 ;
      RECT 41.125000  73.710000 41.925000  74.510000 ;
      RECT 41.125000  75.390000 41.925000  76.190000 ;
      RECT 41.125000  77.070000 41.925000  77.870000 ;
      RECT 41.125000  78.750000 41.925000  79.550000 ;
      RECT 41.125000  80.430000 41.925000  81.230000 ;
      RECT 41.125000  82.110000 41.925000  82.910000 ;
      RECT 41.125000  83.790000 41.925000  84.590000 ;
      RECT 41.125000  85.470000 41.925000  86.270000 ;
      RECT 41.125000  87.150000 41.925000  87.950000 ;
      RECT 41.125000  88.830000 41.925000  89.630000 ;
      RECT 41.125000  90.510000 41.925000  91.310000 ;
      RECT 41.125000  92.190000 41.925000  92.990000 ;
      RECT 41.125000  93.870000 41.925000  94.670000 ;
      RECT 41.125000 176.155000 41.925000 176.955000 ;
      RECT 41.125000 177.775000 41.925000 178.575000 ;
      RECT 41.125000 179.395000 41.925000 180.195000 ;
      RECT 41.125000 181.015000 41.925000 181.815000 ;
      RECT 41.125000 182.635000 41.925000 183.435000 ;
      RECT 41.125000 184.255000 41.925000 185.055000 ;
      RECT 41.125000 185.875000 41.925000 186.675000 ;
      RECT 41.125000 187.495000 41.925000 188.295000 ;
      RECT 41.125000 189.115000 41.925000 189.915000 ;
      RECT 41.125000 190.735000 41.925000 191.535000 ;
      RECT 41.125000 192.355000 41.925000 193.155000 ;
      RECT 41.125000 193.975000 41.925000 194.775000 ;
      RECT 41.125000 195.595000 41.925000 196.395000 ;
      RECT 41.125000 197.215000 41.925000 198.015000 ;
      RECT 41.125000 198.835000 41.925000 199.635000 ;
      RECT 41.130000   9.295000 41.930000  10.095000 ;
      RECT 41.130000  12.325000 41.930000  13.125000 ;
      RECT 42.725000  20.195000 43.525000  20.995000 ;
      RECT 42.725000  23.225000 43.525000  24.025000 ;
      RECT 42.725000  26.245000 43.525000  27.045000 ;
      RECT 42.725000  29.275000 43.525000  30.075000 ;
      RECT 42.730000   2.450000 43.530000   3.250000 ;
      RECT 42.730000   4.360000 43.530000   5.160000 ;
      RECT 42.730000   6.270000 43.530000   7.070000 ;
      RECT 42.730000  15.345000 43.530000  16.145000 ;
      RECT 42.730000  17.175000 43.530000  17.975000 ;
      RECT 42.730000  32.295000 43.530000  33.095000 ;
      RECT 42.730000  34.125000 43.530000  34.925000 ;
      RECT 42.730000  37.145000 43.530000  37.945000 ;
      RECT 42.730000  38.975000 43.530000  39.775000 ;
      RECT 42.730000  41.995000 43.530000  42.795000 ;
      RECT 42.730000  45.025000 43.530000  45.825000 ;
      RECT 42.730000  51.835000 43.530000  52.635000 ;
      RECT 42.730000  58.645000 43.530000  59.445000 ;
      RECT 42.730000  61.475000 43.530000  62.275000 ;
      RECT 42.730000  64.495000 43.530000  65.295000 ;
      RECT 42.730000  67.325000 43.530000  68.125000 ;
      RECT 42.730000  70.350000 43.530000  71.150000 ;
      RECT 42.730000  72.030000 43.530000  72.830000 ;
      RECT 42.730000  73.710000 43.530000  74.510000 ;
      RECT 42.730000  75.390000 43.530000  76.190000 ;
      RECT 42.730000  77.070000 43.530000  77.870000 ;
      RECT 42.730000  78.750000 43.530000  79.550000 ;
      RECT 42.730000  80.430000 43.530000  81.230000 ;
      RECT 42.730000  82.110000 43.530000  82.910000 ;
      RECT 42.730000  83.790000 43.530000  84.590000 ;
      RECT 42.730000  85.470000 43.530000  86.270000 ;
      RECT 42.730000  87.150000 43.530000  87.950000 ;
      RECT 42.730000  88.830000 43.530000  89.630000 ;
      RECT 42.730000  90.510000 43.530000  91.310000 ;
      RECT 42.730000  92.190000 43.530000  92.990000 ;
      RECT 42.730000  93.870000 43.530000  94.670000 ;
      RECT 42.730000 176.155000 43.530000 176.955000 ;
      RECT 42.730000 177.775000 43.530000 178.575000 ;
      RECT 42.730000 179.395000 43.530000 180.195000 ;
      RECT 42.730000 181.015000 43.530000 181.815000 ;
      RECT 42.730000 182.635000 43.530000 183.435000 ;
      RECT 42.730000 184.255000 43.530000 185.055000 ;
      RECT 42.730000 185.875000 43.530000 186.675000 ;
      RECT 42.730000 187.495000 43.530000 188.295000 ;
      RECT 42.730000 189.115000 43.530000 189.915000 ;
      RECT 42.730000 190.735000 43.530000 191.535000 ;
      RECT 42.730000 192.355000 43.530000 193.155000 ;
      RECT 42.730000 193.975000 43.530000 194.775000 ;
      RECT 42.730000 195.595000 43.530000 196.395000 ;
      RECT 42.730000 197.215000 43.530000 198.015000 ;
      RECT 42.730000 198.835000 43.530000 199.635000 ;
      RECT 42.735000   9.295000 43.535000  10.095000 ;
      RECT 42.735000  12.325000 43.535000  13.125000 ;
      RECT 44.330000  20.195000 45.130000  20.995000 ;
      RECT 44.330000  23.225000 45.130000  24.025000 ;
      RECT 44.330000  26.245000 45.130000  27.045000 ;
      RECT 44.330000  29.275000 45.130000  30.075000 ;
      RECT 44.335000   2.450000 45.135000   3.250000 ;
      RECT 44.335000   4.360000 45.135000   5.160000 ;
      RECT 44.335000   6.270000 45.135000   7.070000 ;
      RECT 44.335000  15.345000 45.135000  16.145000 ;
      RECT 44.335000  17.175000 45.135000  17.975000 ;
      RECT 44.335000  32.295000 45.135000  33.095000 ;
      RECT 44.335000  34.125000 45.135000  34.925000 ;
      RECT 44.335000  37.145000 45.135000  37.945000 ;
      RECT 44.335000  38.975000 45.135000  39.775000 ;
      RECT 44.335000  41.995000 45.135000  42.795000 ;
      RECT 44.335000  45.025000 45.135000  45.825000 ;
      RECT 44.335000  51.835000 45.135000  52.635000 ;
      RECT 44.335000  58.645000 45.135000  59.445000 ;
      RECT 44.335000  61.475000 45.135000  62.275000 ;
      RECT 44.335000  64.495000 45.135000  65.295000 ;
      RECT 44.335000  67.325000 45.135000  68.125000 ;
      RECT 44.335000  70.350000 45.135000  71.150000 ;
      RECT 44.335000  72.030000 45.135000  72.830000 ;
      RECT 44.335000  73.710000 45.135000  74.510000 ;
      RECT 44.335000  75.390000 45.135000  76.190000 ;
      RECT 44.335000  77.070000 45.135000  77.870000 ;
      RECT 44.335000  78.750000 45.135000  79.550000 ;
      RECT 44.335000  80.430000 45.135000  81.230000 ;
      RECT 44.335000  82.110000 45.135000  82.910000 ;
      RECT 44.335000  83.790000 45.135000  84.590000 ;
      RECT 44.335000  85.470000 45.135000  86.270000 ;
      RECT 44.335000  87.150000 45.135000  87.950000 ;
      RECT 44.335000  88.830000 45.135000  89.630000 ;
      RECT 44.335000  90.510000 45.135000  91.310000 ;
      RECT 44.335000  92.190000 45.135000  92.990000 ;
      RECT 44.335000  93.870000 45.135000  94.670000 ;
      RECT 44.335000 176.155000 45.135000 176.955000 ;
      RECT 44.335000 177.775000 45.135000 178.575000 ;
      RECT 44.335000 179.395000 45.135000 180.195000 ;
      RECT 44.335000 181.015000 45.135000 181.815000 ;
      RECT 44.335000 182.635000 45.135000 183.435000 ;
      RECT 44.335000 184.255000 45.135000 185.055000 ;
      RECT 44.335000 185.875000 45.135000 186.675000 ;
      RECT 44.335000 187.495000 45.135000 188.295000 ;
      RECT 44.335000 189.115000 45.135000 189.915000 ;
      RECT 44.335000 190.735000 45.135000 191.535000 ;
      RECT 44.335000 192.355000 45.135000 193.155000 ;
      RECT 44.335000 193.975000 45.135000 194.775000 ;
      RECT 44.335000 195.595000 45.135000 196.395000 ;
      RECT 44.335000 197.215000 45.135000 198.015000 ;
      RECT 44.335000 198.835000 45.135000 199.635000 ;
      RECT 44.340000   9.295000 45.140000  10.095000 ;
      RECT 44.340000  12.325000 45.140000  13.125000 ;
      RECT 45.935000  20.195000 46.735000  20.995000 ;
      RECT 45.935000  23.225000 46.735000  24.025000 ;
      RECT 45.935000  26.245000 46.735000  27.045000 ;
      RECT 45.935000  29.275000 46.735000  30.075000 ;
      RECT 45.940000   2.450000 46.740000   3.250000 ;
      RECT 45.940000   4.360000 46.740000   5.160000 ;
      RECT 45.940000   6.270000 46.740000   7.070000 ;
      RECT 45.940000  15.345000 46.740000  16.145000 ;
      RECT 45.940000  17.175000 46.740000  17.975000 ;
      RECT 45.940000  32.295000 46.740000  33.095000 ;
      RECT 45.940000  34.125000 46.740000  34.925000 ;
      RECT 45.940000  37.145000 46.740000  37.945000 ;
      RECT 45.940000  38.975000 46.740000  39.775000 ;
      RECT 45.940000  41.995000 46.740000  42.795000 ;
      RECT 45.940000  45.025000 46.740000  45.825000 ;
      RECT 45.940000  51.835000 46.740000  52.635000 ;
      RECT 45.940000  58.645000 46.740000  59.445000 ;
      RECT 45.940000  61.475000 46.740000  62.275000 ;
      RECT 45.940000  64.495000 46.740000  65.295000 ;
      RECT 45.940000  67.325000 46.740000  68.125000 ;
      RECT 45.940000  70.350000 46.740000  71.150000 ;
      RECT 45.940000  72.030000 46.740000  72.830000 ;
      RECT 45.940000  73.710000 46.740000  74.510000 ;
      RECT 45.940000  75.390000 46.740000  76.190000 ;
      RECT 45.940000  77.070000 46.740000  77.870000 ;
      RECT 45.940000  78.750000 46.740000  79.550000 ;
      RECT 45.940000  80.430000 46.740000  81.230000 ;
      RECT 45.940000  82.110000 46.740000  82.910000 ;
      RECT 45.940000  83.790000 46.740000  84.590000 ;
      RECT 45.940000  85.470000 46.740000  86.270000 ;
      RECT 45.940000  87.150000 46.740000  87.950000 ;
      RECT 45.940000  88.830000 46.740000  89.630000 ;
      RECT 45.940000  90.510000 46.740000  91.310000 ;
      RECT 45.940000  92.190000 46.740000  92.990000 ;
      RECT 45.940000  93.870000 46.740000  94.670000 ;
      RECT 45.940000 176.155000 46.740000 176.955000 ;
      RECT 45.940000 177.775000 46.740000 178.575000 ;
      RECT 45.940000 179.395000 46.740000 180.195000 ;
      RECT 45.940000 181.015000 46.740000 181.815000 ;
      RECT 45.940000 182.635000 46.740000 183.435000 ;
      RECT 45.940000 184.255000 46.740000 185.055000 ;
      RECT 45.940000 185.875000 46.740000 186.675000 ;
      RECT 45.940000 187.495000 46.740000 188.295000 ;
      RECT 45.940000 189.115000 46.740000 189.915000 ;
      RECT 45.940000 190.735000 46.740000 191.535000 ;
      RECT 45.940000 192.355000 46.740000 193.155000 ;
      RECT 45.940000 193.975000 46.740000 194.775000 ;
      RECT 45.940000 195.595000 46.740000 196.395000 ;
      RECT 45.940000 197.215000 46.740000 198.015000 ;
      RECT 45.940000 198.835000 46.740000 199.635000 ;
      RECT 45.945000   9.295000 46.745000  10.095000 ;
      RECT 45.945000  12.325000 46.745000  13.125000 ;
      RECT 47.540000  20.195000 48.340000  20.995000 ;
      RECT 47.540000  23.225000 48.340000  24.025000 ;
      RECT 47.540000  26.245000 48.340000  27.045000 ;
      RECT 47.540000  29.275000 48.340000  30.075000 ;
      RECT 47.545000   2.450000 48.345000   3.250000 ;
      RECT 47.545000   4.360000 48.345000   5.160000 ;
      RECT 47.545000   6.270000 48.345000   7.070000 ;
      RECT 47.545000  15.345000 48.345000  16.145000 ;
      RECT 47.545000  17.175000 48.345000  17.975000 ;
      RECT 47.545000  32.295000 48.345000  33.095000 ;
      RECT 47.545000  34.125000 48.345000  34.925000 ;
      RECT 47.545000  37.145000 48.345000  37.945000 ;
      RECT 47.545000  38.975000 48.345000  39.775000 ;
      RECT 47.545000  41.995000 48.345000  42.795000 ;
      RECT 47.545000  45.025000 48.345000  45.825000 ;
      RECT 47.545000  51.835000 48.345000  52.635000 ;
      RECT 47.545000  58.645000 48.345000  59.445000 ;
      RECT 47.545000  61.475000 48.345000  62.275000 ;
      RECT 47.545000  64.495000 48.345000  65.295000 ;
      RECT 47.545000  67.325000 48.345000  68.125000 ;
      RECT 47.545000  70.350000 48.345000  71.150000 ;
      RECT 47.545000  72.030000 48.345000  72.830000 ;
      RECT 47.545000  73.710000 48.345000  74.510000 ;
      RECT 47.545000  75.390000 48.345000  76.190000 ;
      RECT 47.545000  77.070000 48.345000  77.870000 ;
      RECT 47.545000  78.750000 48.345000  79.550000 ;
      RECT 47.545000  80.430000 48.345000  81.230000 ;
      RECT 47.545000  82.110000 48.345000  82.910000 ;
      RECT 47.545000  83.790000 48.345000  84.590000 ;
      RECT 47.545000  85.470000 48.345000  86.270000 ;
      RECT 47.545000  87.150000 48.345000  87.950000 ;
      RECT 47.545000  88.830000 48.345000  89.630000 ;
      RECT 47.545000  90.510000 48.345000  91.310000 ;
      RECT 47.545000  92.190000 48.345000  92.990000 ;
      RECT 47.545000  93.870000 48.345000  94.670000 ;
      RECT 47.545000 176.155000 48.345000 176.955000 ;
      RECT 47.545000 177.775000 48.345000 178.575000 ;
      RECT 47.545000 179.395000 48.345000 180.195000 ;
      RECT 47.545000 181.015000 48.345000 181.815000 ;
      RECT 47.545000 182.635000 48.345000 183.435000 ;
      RECT 47.545000 184.255000 48.345000 185.055000 ;
      RECT 47.545000 185.875000 48.345000 186.675000 ;
      RECT 47.545000 187.495000 48.345000 188.295000 ;
      RECT 47.545000 189.115000 48.345000 189.915000 ;
      RECT 47.545000 190.735000 48.345000 191.535000 ;
      RECT 47.545000 192.355000 48.345000 193.155000 ;
      RECT 47.545000 193.975000 48.345000 194.775000 ;
      RECT 47.545000 195.595000 48.345000 196.395000 ;
      RECT 47.545000 197.215000 48.345000 198.015000 ;
      RECT 47.545000 198.835000 48.345000 199.635000 ;
      RECT 47.550000   9.295000 48.350000  10.095000 ;
      RECT 47.550000  12.325000 48.350000  13.125000 ;
      RECT 49.145000  20.195000 49.945000  20.995000 ;
      RECT 49.145000  23.225000 49.945000  24.025000 ;
      RECT 49.145000  26.245000 49.945000  27.045000 ;
      RECT 49.145000  29.275000 49.945000  30.075000 ;
      RECT 49.150000   2.450000 49.950000   3.250000 ;
      RECT 49.150000   4.360000 49.950000   5.160000 ;
      RECT 49.150000   6.270000 49.950000   7.070000 ;
      RECT 49.150000  15.345000 49.950000  16.145000 ;
      RECT 49.150000  17.175000 49.950000  17.975000 ;
      RECT 49.150000  32.295000 49.950000  33.095000 ;
      RECT 49.150000  34.125000 49.950000  34.925000 ;
      RECT 49.150000  37.145000 49.950000  37.945000 ;
      RECT 49.150000  38.975000 49.950000  39.775000 ;
      RECT 49.150000  41.995000 49.950000  42.795000 ;
      RECT 49.150000  45.025000 49.950000  45.825000 ;
      RECT 49.150000  51.835000 49.950000  52.635000 ;
      RECT 49.150000  58.645000 49.950000  59.445000 ;
      RECT 49.150000  61.475000 49.950000  62.275000 ;
      RECT 49.150000  64.495000 49.950000  65.295000 ;
      RECT 49.150000  67.325000 49.950000  68.125000 ;
      RECT 49.150000  70.350000 49.950000  71.150000 ;
      RECT 49.150000  72.030000 49.950000  72.830000 ;
      RECT 49.150000  73.710000 49.950000  74.510000 ;
      RECT 49.150000  75.390000 49.950000  76.190000 ;
      RECT 49.150000  77.070000 49.950000  77.870000 ;
      RECT 49.150000  78.750000 49.950000  79.550000 ;
      RECT 49.150000  80.430000 49.950000  81.230000 ;
      RECT 49.150000  82.110000 49.950000  82.910000 ;
      RECT 49.150000  83.790000 49.950000  84.590000 ;
      RECT 49.150000  85.470000 49.950000  86.270000 ;
      RECT 49.150000  87.150000 49.950000  87.950000 ;
      RECT 49.150000  88.830000 49.950000  89.630000 ;
      RECT 49.150000  90.510000 49.950000  91.310000 ;
      RECT 49.150000  92.190000 49.950000  92.990000 ;
      RECT 49.150000  93.870000 49.950000  94.670000 ;
      RECT 49.150000 176.155000 49.950000 176.955000 ;
      RECT 49.150000 177.775000 49.950000 178.575000 ;
      RECT 49.150000 179.395000 49.950000 180.195000 ;
      RECT 49.150000 181.015000 49.950000 181.815000 ;
      RECT 49.150000 182.635000 49.950000 183.435000 ;
      RECT 49.150000 184.255000 49.950000 185.055000 ;
      RECT 49.150000 185.875000 49.950000 186.675000 ;
      RECT 49.150000 187.495000 49.950000 188.295000 ;
      RECT 49.150000 189.115000 49.950000 189.915000 ;
      RECT 49.150000 190.735000 49.950000 191.535000 ;
      RECT 49.150000 192.355000 49.950000 193.155000 ;
      RECT 49.150000 193.975000 49.950000 194.775000 ;
      RECT 49.150000 195.595000 49.950000 196.395000 ;
      RECT 49.150000 197.215000 49.950000 198.015000 ;
      RECT 49.150000 198.835000 49.950000 199.635000 ;
      RECT 49.155000   9.295000 49.955000  10.095000 ;
      RECT 49.155000  12.325000 49.955000  13.125000 ;
      RECT 50.750000  20.195000 51.550000  20.995000 ;
      RECT 50.750000  23.225000 51.550000  24.025000 ;
      RECT 50.750000  26.245000 51.550000  27.045000 ;
      RECT 50.750000  29.275000 51.550000  30.075000 ;
      RECT 50.755000   2.450000 51.555000   3.250000 ;
      RECT 50.755000   4.360000 51.555000   5.160000 ;
      RECT 50.755000   6.270000 51.555000   7.070000 ;
      RECT 50.755000  15.345000 51.555000  16.145000 ;
      RECT 50.755000  17.175000 51.555000  17.975000 ;
      RECT 50.755000  32.295000 51.555000  33.095000 ;
      RECT 50.755000  34.125000 51.555000  34.925000 ;
      RECT 50.755000  37.145000 51.555000  37.945000 ;
      RECT 50.755000  38.975000 51.555000  39.775000 ;
      RECT 50.755000  41.995000 51.555000  42.795000 ;
      RECT 50.755000  45.025000 51.555000  45.825000 ;
      RECT 50.755000  51.835000 51.555000  52.635000 ;
      RECT 50.755000  58.645000 51.555000  59.445000 ;
      RECT 50.755000  61.475000 51.555000  62.275000 ;
      RECT 50.755000  64.495000 51.555000  65.295000 ;
      RECT 50.755000  67.325000 51.555000  68.125000 ;
      RECT 50.755000  70.350000 51.555000  71.150000 ;
      RECT 50.755000  72.030000 51.555000  72.830000 ;
      RECT 50.755000  73.710000 51.555000  74.510000 ;
      RECT 50.755000  75.390000 51.555000  76.190000 ;
      RECT 50.755000  77.070000 51.555000  77.870000 ;
      RECT 50.755000  78.750000 51.555000  79.550000 ;
      RECT 50.755000  80.430000 51.555000  81.230000 ;
      RECT 50.755000  82.110000 51.555000  82.910000 ;
      RECT 50.755000  83.790000 51.555000  84.590000 ;
      RECT 50.755000  85.470000 51.555000  86.270000 ;
      RECT 50.755000  87.150000 51.555000  87.950000 ;
      RECT 50.755000  88.830000 51.555000  89.630000 ;
      RECT 50.755000  90.510000 51.555000  91.310000 ;
      RECT 50.755000  92.190000 51.555000  92.990000 ;
      RECT 50.755000  93.870000 51.555000  94.670000 ;
      RECT 50.755000 176.155000 51.555000 176.955000 ;
      RECT 50.755000 177.775000 51.555000 178.575000 ;
      RECT 50.755000 179.395000 51.555000 180.195000 ;
      RECT 50.755000 181.015000 51.555000 181.815000 ;
      RECT 50.755000 182.635000 51.555000 183.435000 ;
      RECT 50.755000 184.255000 51.555000 185.055000 ;
      RECT 50.755000 185.875000 51.555000 186.675000 ;
      RECT 50.755000 187.495000 51.555000 188.295000 ;
      RECT 50.755000 189.115000 51.555000 189.915000 ;
      RECT 50.755000 190.735000 51.555000 191.535000 ;
      RECT 50.755000 192.355000 51.555000 193.155000 ;
      RECT 50.755000 193.975000 51.555000 194.775000 ;
      RECT 50.755000 195.595000 51.555000 196.395000 ;
      RECT 50.755000 197.215000 51.555000 198.015000 ;
      RECT 50.755000 198.835000 51.555000 199.635000 ;
      RECT 50.760000   9.295000 51.560000  10.095000 ;
      RECT 50.760000  12.325000 51.560000  13.125000 ;
      RECT 52.355000  20.195000 53.155000  20.995000 ;
      RECT 52.355000  23.225000 53.155000  24.025000 ;
      RECT 52.355000  26.245000 53.155000  27.045000 ;
      RECT 52.355000  29.275000 53.155000  30.075000 ;
      RECT 52.360000   2.450000 53.160000   3.250000 ;
      RECT 52.360000   4.360000 53.160000   5.160000 ;
      RECT 52.360000   6.270000 53.160000   7.070000 ;
      RECT 52.360000  15.345000 53.160000  16.145000 ;
      RECT 52.360000  17.175000 53.160000  17.975000 ;
      RECT 52.360000  32.295000 53.160000  33.095000 ;
      RECT 52.360000  34.125000 53.160000  34.925000 ;
      RECT 52.360000  37.145000 53.160000  37.945000 ;
      RECT 52.360000  38.975000 53.160000  39.775000 ;
      RECT 52.360000  41.995000 53.160000  42.795000 ;
      RECT 52.360000  45.025000 53.160000  45.825000 ;
      RECT 52.360000  51.835000 53.160000  52.635000 ;
      RECT 52.360000  58.645000 53.160000  59.445000 ;
      RECT 52.360000  61.475000 53.160000  62.275000 ;
      RECT 52.360000  64.495000 53.160000  65.295000 ;
      RECT 52.360000  67.325000 53.160000  68.125000 ;
      RECT 52.360000  70.350000 53.160000  71.150000 ;
      RECT 52.360000  72.030000 53.160000  72.830000 ;
      RECT 52.360000  73.710000 53.160000  74.510000 ;
      RECT 52.360000  75.390000 53.160000  76.190000 ;
      RECT 52.360000  77.070000 53.160000  77.870000 ;
      RECT 52.360000  78.750000 53.160000  79.550000 ;
      RECT 52.360000  80.430000 53.160000  81.230000 ;
      RECT 52.360000  82.110000 53.160000  82.910000 ;
      RECT 52.360000  83.790000 53.160000  84.590000 ;
      RECT 52.360000  85.470000 53.160000  86.270000 ;
      RECT 52.360000  87.150000 53.160000  87.950000 ;
      RECT 52.360000  88.830000 53.160000  89.630000 ;
      RECT 52.360000  90.510000 53.160000  91.310000 ;
      RECT 52.360000  92.190000 53.160000  92.990000 ;
      RECT 52.360000  93.870000 53.160000  94.670000 ;
      RECT 52.360000 176.155000 53.160000 176.955000 ;
      RECT 52.360000 177.775000 53.160000 178.575000 ;
      RECT 52.360000 179.395000 53.160000 180.195000 ;
      RECT 52.360000 181.015000 53.160000 181.815000 ;
      RECT 52.360000 182.635000 53.160000 183.435000 ;
      RECT 52.360000 184.255000 53.160000 185.055000 ;
      RECT 52.360000 185.875000 53.160000 186.675000 ;
      RECT 52.360000 187.495000 53.160000 188.295000 ;
      RECT 52.360000 189.115000 53.160000 189.915000 ;
      RECT 52.360000 190.735000 53.160000 191.535000 ;
      RECT 52.360000 192.355000 53.160000 193.155000 ;
      RECT 52.360000 193.975000 53.160000 194.775000 ;
      RECT 52.360000 195.595000 53.160000 196.395000 ;
      RECT 52.360000 197.215000 53.160000 198.015000 ;
      RECT 52.360000 198.835000 53.160000 199.635000 ;
      RECT 52.365000   9.295000 53.165000  10.095000 ;
      RECT 52.365000  12.325000 53.165000  13.125000 ;
      RECT 53.960000  20.195000 54.760000  20.995000 ;
      RECT 53.960000  23.225000 54.760000  24.025000 ;
      RECT 53.960000  26.245000 54.760000  27.045000 ;
      RECT 53.960000  29.275000 54.760000  30.075000 ;
      RECT 53.965000   2.450000 54.765000   3.250000 ;
      RECT 53.965000   4.360000 54.765000   5.160000 ;
      RECT 53.965000   6.270000 54.765000   7.070000 ;
      RECT 53.965000  15.345000 54.765000  16.145000 ;
      RECT 53.965000  17.175000 54.765000  17.975000 ;
      RECT 53.965000  32.295000 54.765000  33.095000 ;
      RECT 53.965000  34.125000 54.765000  34.925000 ;
      RECT 53.965000  37.145000 54.765000  37.945000 ;
      RECT 53.965000  38.975000 54.765000  39.775000 ;
      RECT 53.965000  41.995000 54.765000  42.795000 ;
      RECT 53.965000  45.025000 54.765000  45.825000 ;
      RECT 53.965000  51.835000 54.765000  52.635000 ;
      RECT 53.965000  58.645000 54.765000  59.445000 ;
      RECT 53.965000  61.475000 54.765000  62.275000 ;
      RECT 53.965000  64.495000 54.765000  65.295000 ;
      RECT 53.965000  67.325000 54.765000  68.125000 ;
      RECT 53.965000  70.350000 54.765000  71.150000 ;
      RECT 53.965000  72.030000 54.765000  72.830000 ;
      RECT 53.965000  73.710000 54.765000  74.510000 ;
      RECT 53.965000  75.390000 54.765000  76.190000 ;
      RECT 53.965000  77.070000 54.765000  77.870000 ;
      RECT 53.965000  78.750000 54.765000  79.550000 ;
      RECT 53.965000  80.430000 54.765000  81.230000 ;
      RECT 53.965000  82.110000 54.765000  82.910000 ;
      RECT 53.965000  83.790000 54.765000  84.590000 ;
      RECT 53.965000  85.470000 54.765000  86.270000 ;
      RECT 53.965000  87.150000 54.765000  87.950000 ;
      RECT 53.965000  88.830000 54.765000  89.630000 ;
      RECT 53.965000  90.510000 54.765000  91.310000 ;
      RECT 53.965000  92.190000 54.765000  92.990000 ;
      RECT 53.965000  93.870000 54.765000  94.670000 ;
      RECT 53.965000 176.155000 54.765000 176.955000 ;
      RECT 53.965000 177.775000 54.765000 178.575000 ;
      RECT 53.965000 179.395000 54.765000 180.195000 ;
      RECT 53.965000 181.015000 54.765000 181.815000 ;
      RECT 53.965000 182.635000 54.765000 183.435000 ;
      RECT 53.965000 184.255000 54.765000 185.055000 ;
      RECT 53.965000 185.875000 54.765000 186.675000 ;
      RECT 53.965000 187.495000 54.765000 188.295000 ;
      RECT 53.965000 189.115000 54.765000 189.915000 ;
      RECT 53.965000 190.735000 54.765000 191.535000 ;
      RECT 53.965000 192.355000 54.765000 193.155000 ;
      RECT 53.965000 193.975000 54.765000 194.775000 ;
      RECT 53.965000 195.595000 54.765000 196.395000 ;
      RECT 53.965000 197.215000 54.765000 198.015000 ;
      RECT 53.965000 198.835000 54.765000 199.635000 ;
      RECT 53.970000   9.295000 54.770000  10.095000 ;
      RECT 53.970000  12.325000 54.770000  13.125000 ;
      RECT 55.565000  20.195000 56.365000  20.995000 ;
      RECT 55.565000  23.225000 56.365000  24.025000 ;
      RECT 55.565000  26.245000 56.365000  27.045000 ;
      RECT 55.565000  29.275000 56.365000  30.075000 ;
      RECT 55.570000   2.450000 56.370000   3.250000 ;
      RECT 55.570000   4.360000 56.370000   5.160000 ;
      RECT 55.570000   6.270000 56.370000   7.070000 ;
      RECT 55.570000  15.345000 56.370000  16.145000 ;
      RECT 55.570000  17.175000 56.370000  17.975000 ;
      RECT 55.570000  32.295000 56.370000  33.095000 ;
      RECT 55.570000  34.125000 56.370000  34.925000 ;
      RECT 55.570000  37.145000 56.370000  37.945000 ;
      RECT 55.570000  38.975000 56.370000  39.775000 ;
      RECT 55.570000  41.995000 56.370000  42.795000 ;
      RECT 55.570000  45.025000 56.370000  45.825000 ;
      RECT 55.570000  51.835000 56.370000  52.635000 ;
      RECT 55.570000  58.645000 56.370000  59.445000 ;
      RECT 55.570000  61.475000 56.370000  62.275000 ;
      RECT 55.570000  64.495000 56.370000  65.295000 ;
      RECT 55.570000  67.325000 56.370000  68.125000 ;
      RECT 55.570000  70.350000 56.370000  71.150000 ;
      RECT 55.570000  72.030000 56.370000  72.830000 ;
      RECT 55.570000  73.710000 56.370000  74.510000 ;
      RECT 55.570000  75.390000 56.370000  76.190000 ;
      RECT 55.570000  77.070000 56.370000  77.870000 ;
      RECT 55.570000  78.750000 56.370000  79.550000 ;
      RECT 55.570000  80.430000 56.370000  81.230000 ;
      RECT 55.570000  82.110000 56.370000  82.910000 ;
      RECT 55.570000  83.790000 56.370000  84.590000 ;
      RECT 55.570000  85.470000 56.370000  86.270000 ;
      RECT 55.570000  87.150000 56.370000  87.950000 ;
      RECT 55.570000  88.830000 56.370000  89.630000 ;
      RECT 55.570000  90.510000 56.370000  91.310000 ;
      RECT 55.570000  92.190000 56.370000  92.990000 ;
      RECT 55.570000  93.870000 56.370000  94.670000 ;
      RECT 55.570000 176.155000 56.370000 176.955000 ;
      RECT 55.570000 177.775000 56.370000 178.575000 ;
      RECT 55.570000 179.395000 56.370000 180.195000 ;
      RECT 55.570000 181.015000 56.370000 181.815000 ;
      RECT 55.570000 182.635000 56.370000 183.435000 ;
      RECT 55.570000 184.255000 56.370000 185.055000 ;
      RECT 55.570000 185.875000 56.370000 186.675000 ;
      RECT 55.570000 187.495000 56.370000 188.295000 ;
      RECT 55.570000 189.115000 56.370000 189.915000 ;
      RECT 55.570000 190.735000 56.370000 191.535000 ;
      RECT 55.570000 192.355000 56.370000 193.155000 ;
      RECT 55.570000 193.975000 56.370000 194.775000 ;
      RECT 55.570000 195.595000 56.370000 196.395000 ;
      RECT 55.570000 197.215000 56.370000 198.015000 ;
      RECT 55.570000 198.835000 56.370000 199.635000 ;
      RECT 55.575000   9.295000 56.375000  10.095000 ;
      RECT 55.575000  12.325000 56.375000  13.125000 ;
      RECT 57.170000  20.195000 57.970000  20.995000 ;
      RECT 57.170000  23.225000 57.970000  24.025000 ;
      RECT 57.170000  26.245000 57.970000  27.045000 ;
      RECT 57.170000  29.275000 57.970000  30.075000 ;
      RECT 57.175000   2.450000 57.975000   3.250000 ;
      RECT 57.175000   4.360000 57.975000   5.160000 ;
      RECT 57.175000   6.270000 57.975000   7.070000 ;
      RECT 57.175000   9.295000 57.975000  10.095000 ;
      RECT 57.175000  12.325000 57.975000  13.125000 ;
      RECT 57.175000  15.345000 57.975000  16.145000 ;
      RECT 57.175000  17.175000 57.975000  17.975000 ;
      RECT 57.175000  32.295000 57.975000  33.095000 ;
      RECT 57.175000  34.125000 57.975000  34.925000 ;
      RECT 57.175000  37.145000 57.975000  37.945000 ;
      RECT 57.175000  38.975000 57.975000  39.775000 ;
      RECT 57.175000  41.995000 57.975000  42.795000 ;
      RECT 57.175000  45.025000 57.975000  45.825000 ;
      RECT 57.175000  51.835000 57.975000  52.635000 ;
      RECT 57.175000  58.645000 57.975000  59.445000 ;
      RECT 57.175000  61.475000 57.975000  62.275000 ;
      RECT 57.175000  64.495000 57.975000  65.295000 ;
      RECT 57.175000  67.325000 57.975000  68.125000 ;
      RECT 57.175000  70.350000 57.975000  71.150000 ;
      RECT 57.175000  72.030000 57.975000  72.830000 ;
      RECT 57.175000  73.710000 57.975000  74.510000 ;
      RECT 57.175000  75.390000 57.975000  76.190000 ;
      RECT 57.175000  77.070000 57.975000  77.870000 ;
      RECT 57.175000  78.750000 57.975000  79.550000 ;
      RECT 57.175000  80.430000 57.975000  81.230000 ;
      RECT 57.175000  82.110000 57.975000  82.910000 ;
      RECT 57.175000  83.790000 57.975000  84.590000 ;
      RECT 57.175000  85.470000 57.975000  86.270000 ;
      RECT 57.175000  87.150000 57.975000  87.950000 ;
      RECT 57.175000  88.830000 57.975000  89.630000 ;
      RECT 57.175000  90.510000 57.975000  91.310000 ;
      RECT 57.175000  92.190000 57.975000  92.990000 ;
      RECT 57.175000  93.870000 57.975000  94.670000 ;
      RECT 57.175000 176.155000 57.975000 176.955000 ;
      RECT 57.175000 177.775000 57.975000 178.575000 ;
      RECT 57.175000 179.395000 57.975000 180.195000 ;
      RECT 57.175000 181.015000 57.975000 181.815000 ;
      RECT 57.175000 182.635000 57.975000 183.435000 ;
      RECT 57.175000 184.255000 57.975000 185.055000 ;
      RECT 57.175000 185.875000 57.975000 186.675000 ;
      RECT 57.175000 187.495000 57.975000 188.295000 ;
      RECT 57.175000 189.115000 57.975000 189.915000 ;
      RECT 57.175000 190.735000 57.975000 191.535000 ;
      RECT 57.175000 192.355000 57.975000 193.155000 ;
      RECT 57.175000 193.975000 57.975000 194.775000 ;
      RECT 57.175000 195.595000 57.975000 196.395000 ;
      RECT 57.175000 197.215000 57.975000 198.015000 ;
      RECT 57.175000 198.835000 57.975000 199.635000 ;
      RECT 58.775000   9.295000 59.575000  10.095000 ;
      RECT 58.775000  12.325000 59.575000  13.125000 ;
      RECT 58.775000  20.195000 59.575000  20.995000 ;
      RECT 58.775000  23.225000 59.575000  24.025000 ;
      RECT 58.775000  26.245000 59.575000  27.045000 ;
      RECT 58.775000  29.275000 59.575000  30.075000 ;
      RECT 58.775000  41.995000 59.575000  42.795000 ;
      RECT 58.775000  45.025000 59.575000  45.825000 ;
      RECT 58.780000   2.450000 59.580000   3.250000 ;
      RECT 58.780000   4.360000 59.580000   5.160000 ;
      RECT 58.780000   6.270000 59.580000   7.070000 ;
      RECT 58.780000  15.345000 59.580000  16.145000 ;
      RECT 58.780000  17.175000 59.580000  17.975000 ;
      RECT 58.780000  32.295000 59.580000  33.095000 ;
      RECT 58.780000  34.125000 59.580000  34.925000 ;
      RECT 58.780000  37.145000 59.580000  37.945000 ;
      RECT 58.780000  38.975000 59.580000  39.775000 ;
      RECT 58.780000  51.835000 59.580000  52.635000 ;
      RECT 58.780000  58.645000 59.580000  59.445000 ;
      RECT 58.780000  61.475000 59.580000  62.275000 ;
      RECT 58.780000  64.495000 59.580000  65.295000 ;
      RECT 58.780000  67.325000 59.580000  68.125000 ;
      RECT 58.780000  70.350000 59.580000  71.150000 ;
      RECT 58.780000  72.030000 59.580000  72.830000 ;
      RECT 58.780000  73.710000 59.580000  74.510000 ;
      RECT 58.780000  75.390000 59.580000  76.190000 ;
      RECT 58.780000  77.070000 59.580000  77.870000 ;
      RECT 58.780000  78.750000 59.580000  79.550000 ;
      RECT 58.780000  80.430000 59.580000  81.230000 ;
      RECT 58.780000  82.110000 59.580000  82.910000 ;
      RECT 58.780000  83.790000 59.580000  84.590000 ;
      RECT 58.780000  85.470000 59.580000  86.270000 ;
      RECT 58.780000  87.150000 59.580000  87.950000 ;
      RECT 58.780000  88.830000 59.580000  89.630000 ;
      RECT 58.780000  90.510000 59.580000  91.310000 ;
      RECT 58.780000  92.190000 59.580000  92.990000 ;
      RECT 58.780000  93.870000 59.580000  94.670000 ;
      RECT 58.780000 176.155000 59.580000 176.955000 ;
      RECT 58.780000 177.775000 59.580000 178.575000 ;
      RECT 58.780000 179.395000 59.580000 180.195000 ;
      RECT 58.780000 181.015000 59.580000 181.815000 ;
      RECT 58.780000 182.635000 59.580000 183.435000 ;
      RECT 58.780000 184.255000 59.580000 185.055000 ;
      RECT 58.780000 185.875000 59.580000 186.675000 ;
      RECT 58.780000 187.495000 59.580000 188.295000 ;
      RECT 58.780000 189.115000 59.580000 189.915000 ;
      RECT 58.780000 190.735000 59.580000 191.535000 ;
      RECT 58.780000 192.355000 59.580000 193.155000 ;
      RECT 58.780000 193.975000 59.580000 194.775000 ;
      RECT 58.780000 195.595000 59.580000 196.395000 ;
      RECT 58.780000 197.215000 59.580000 198.015000 ;
      RECT 58.780000 198.835000 59.580000 199.635000 ;
      RECT 60.375000   9.295000 61.175000  10.095000 ;
      RECT 60.375000  12.325000 61.175000  13.125000 ;
      RECT 60.375000  20.195000 61.175000  20.995000 ;
      RECT 60.375000  23.225000 61.175000  24.025000 ;
      RECT 60.375000  41.995000 61.175000  42.795000 ;
      RECT 60.375000  45.025000 61.175000  45.825000 ;
      RECT 60.380000   2.450000 61.180000   3.250000 ;
      RECT 60.380000   4.360000 61.180000   5.160000 ;
      RECT 60.380000   6.270000 61.180000   7.070000 ;
      RECT 60.380000  15.345000 61.180000  16.145000 ;
      RECT 60.380000  17.175000 61.180000  17.975000 ;
      RECT 60.380000  26.245000 61.180000  27.045000 ;
      RECT 60.380000  29.275000 61.180000  30.075000 ;
      RECT 60.380000  32.295000 61.180000  33.095000 ;
      RECT 60.380000  34.125000 61.180000  34.925000 ;
      RECT 60.380000  51.835000 61.180000  52.635000 ;
      RECT 60.380000  64.495000 61.180000  65.295000 ;
      RECT 60.380000  67.325000 61.180000  68.125000 ;
      RECT 60.380000  70.350000 61.180000  71.150000 ;
      RECT 60.380000  72.030000 61.180000  72.830000 ;
      RECT 60.380000  73.710000 61.180000  74.510000 ;
      RECT 60.380000  75.390000 61.180000  76.190000 ;
      RECT 60.380000  77.070000 61.180000  77.870000 ;
      RECT 60.380000  78.750000 61.180000  79.550000 ;
      RECT 60.380000  80.430000 61.180000  81.230000 ;
      RECT 60.380000  82.110000 61.180000  82.910000 ;
      RECT 60.380000  83.790000 61.180000  84.590000 ;
      RECT 60.380000  85.470000 61.180000  86.270000 ;
      RECT 60.380000  87.150000 61.180000  87.950000 ;
      RECT 60.380000  88.830000 61.180000  89.630000 ;
      RECT 60.380000  90.510000 61.180000  91.310000 ;
      RECT 60.380000  92.190000 61.180000  92.990000 ;
      RECT 60.380000  93.870000 61.180000  94.670000 ;
      RECT 60.380000 176.155000 61.180000 176.955000 ;
      RECT 60.380000 177.775000 61.180000 178.575000 ;
      RECT 60.380000 179.395000 61.180000 180.195000 ;
      RECT 60.380000 181.015000 61.180000 181.815000 ;
      RECT 60.380000 182.635000 61.180000 183.435000 ;
      RECT 60.380000 184.255000 61.180000 185.055000 ;
      RECT 60.380000 185.875000 61.180000 186.675000 ;
      RECT 60.380000 187.495000 61.180000 188.295000 ;
      RECT 60.380000 189.115000 61.180000 189.915000 ;
      RECT 60.380000 190.735000 61.180000 191.535000 ;
      RECT 60.380000 192.355000 61.180000 193.155000 ;
      RECT 60.380000 193.975000 61.180000 194.775000 ;
      RECT 60.380000 195.595000 61.180000 196.395000 ;
      RECT 60.380000 197.215000 61.180000 198.015000 ;
      RECT 60.380000 198.835000 61.180000 199.635000 ;
      RECT 60.385000  37.145000 61.185000  37.945000 ;
      RECT 60.385000  38.975000 61.185000  39.775000 ;
      RECT 60.385000  58.645000 61.185000  59.445000 ;
      RECT 60.385000  61.475000 61.185000  62.275000 ;
      RECT 61.975000   9.295000 62.775000  10.095000 ;
      RECT 61.975000  12.325000 62.775000  13.125000 ;
      RECT 61.975000  20.195000 62.775000  20.995000 ;
      RECT 61.975000  23.225000 62.775000  24.025000 ;
      RECT 61.975000  41.995000 62.775000  42.795000 ;
      RECT 61.975000  45.025000 62.775000  45.825000 ;
      RECT 61.980000   2.450000 62.780000   3.250000 ;
      RECT 61.980000   4.360000 62.780000   5.160000 ;
      RECT 61.980000   6.270000 62.780000   7.070000 ;
      RECT 61.980000  15.345000 62.780000  16.145000 ;
      RECT 61.980000  17.175000 62.780000  17.975000 ;
      RECT 61.980000  26.245000 62.780000  27.045000 ;
      RECT 61.980000  29.275000 62.780000  30.075000 ;
      RECT 61.980000  32.295000 62.780000  33.095000 ;
      RECT 61.980000  34.125000 62.780000  34.925000 ;
      RECT 61.980000  51.835000 62.780000  52.635000 ;
      RECT 61.980000  64.495000 62.780000  65.295000 ;
      RECT 61.980000  67.325000 62.780000  68.125000 ;
      RECT 61.980000  70.350000 62.780000  71.150000 ;
      RECT 61.980000  72.030000 62.780000  72.830000 ;
      RECT 61.980000  73.710000 62.780000  74.510000 ;
      RECT 61.980000  75.390000 62.780000  76.190000 ;
      RECT 61.980000  77.070000 62.780000  77.870000 ;
      RECT 61.980000  78.750000 62.780000  79.550000 ;
      RECT 61.980000  80.430000 62.780000  81.230000 ;
      RECT 61.980000  82.110000 62.780000  82.910000 ;
      RECT 61.980000  83.790000 62.780000  84.590000 ;
      RECT 61.980000  85.470000 62.780000  86.270000 ;
      RECT 61.980000  87.150000 62.780000  87.950000 ;
      RECT 61.980000  88.830000 62.780000  89.630000 ;
      RECT 61.980000  90.510000 62.780000  91.310000 ;
      RECT 61.980000  92.190000 62.780000  92.990000 ;
      RECT 61.980000  93.870000 62.780000  94.670000 ;
      RECT 61.980000 176.155000 62.780000 176.955000 ;
      RECT 61.980000 177.775000 62.780000 178.575000 ;
      RECT 61.980000 179.395000 62.780000 180.195000 ;
      RECT 61.980000 181.015000 62.780000 181.815000 ;
      RECT 61.980000 182.635000 62.780000 183.435000 ;
      RECT 61.980000 184.255000 62.780000 185.055000 ;
      RECT 61.980000 185.875000 62.780000 186.675000 ;
      RECT 61.980000 187.495000 62.780000 188.295000 ;
      RECT 61.980000 189.115000 62.780000 189.915000 ;
      RECT 61.980000 190.735000 62.780000 191.535000 ;
      RECT 61.980000 192.355000 62.780000 193.155000 ;
      RECT 61.980000 193.975000 62.780000 194.775000 ;
      RECT 61.980000 195.595000 62.780000 196.395000 ;
      RECT 61.980000 197.215000 62.780000 198.015000 ;
      RECT 61.980000 198.835000 62.780000 199.635000 ;
      RECT 61.985000  37.145000 62.785000  37.945000 ;
      RECT 61.985000  38.975000 62.785000  39.775000 ;
      RECT 61.985000  58.645000 62.785000  59.445000 ;
      RECT 61.985000  61.475000 62.785000  62.275000 ;
      RECT 63.575000   9.295000 64.375000  10.095000 ;
      RECT 63.575000  12.325000 64.375000  13.125000 ;
      RECT 63.575000  20.195000 64.375000  20.995000 ;
      RECT 63.575000  23.225000 64.375000  24.025000 ;
      RECT 63.575000  41.995000 64.375000  42.795000 ;
      RECT 63.575000  45.025000 64.375000  45.825000 ;
      RECT 63.580000   2.450000 64.380000   3.250000 ;
      RECT 63.580000   4.360000 64.380000   5.160000 ;
      RECT 63.580000   6.270000 64.380000   7.070000 ;
      RECT 63.580000  15.345000 64.380000  16.145000 ;
      RECT 63.580000  17.175000 64.380000  17.975000 ;
      RECT 63.580000  26.245000 64.380000  27.045000 ;
      RECT 63.580000  29.275000 64.380000  30.075000 ;
      RECT 63.580000  32.295000 64.380000  33.095000 ;
      RECT 63.580000  34.125000 64.380000  34.925000 ;
      RECT 63.580000  51.835000 64.380000  52.635000 ;
      RECT 63.580000  64.495000 64.380000  65.295000 ;
      RECT 63.580000  67.325000 64.380000  68.125000 ;
      RECT 63.580000  70.350000 64.380000  71.150000 ;
      RECT 63.580000  72.030000 64.380000  72.830000 ;
      RECT 63.580000  73.710000 64.380000  74.510000 ;
      RECT 63.580000  75.390000 64.380000  76.190000 ;
      RECT 63.580000  77.070000 64.380000  77.870000 ;
      RECT 63.580000  78.750000 64.380000  79.550000 ;
      RECT 63.580000  80.430000 64.380000  81.230000 ;
      RECT 63.580000  82.110000 64.380000  82.910000 ;
      RECT 63.580000  83.790000 64.380000  84.590000 ;
      RECT 63.580000  85.470000 64.380000  86.270000 ;
      RECT 63.580000  87.150000 64.380000  87.950000 ;
      RECT 63.580000  88.830000 64.380000  89.630000 ;
      RECT 63.580000  90.510000 64.380000  91.310000 ;
      RECT 63.580000  92.190000 64.380000  92.990000 ;
      RECT 63.580000  93.870000 64.380000  94.670000 ;
      RECT 63.580000 176.155000 64.380000 176.955000 ;
      RECT 63.580000 177.775000 64.380000 178.575000 ;
      RECT 63.580000 179.395000 64.380000 180.195000 ;
      RECT 63.580000 181.015000 64.380000 181.815000 ;
      RECT 63.580000 182.635000 64.380000 183.435000 ;
      RECT 63.580000 184.255000 64.380000 185.055000 ;
      RECT 63.580000 185.875000 64.380000 186.675000 ;
      RECT 63.580000 187.495000 64.380000 188.295000 ;
      RECT 63.580000 189.115000 64.380000 189.915000 ;
      RECT 63.580000 190.735000 64.380000 191.535000 ;
      RECT 63.580000 192.355000 64.380000 193.155000 ;
      RECT 63.580000 193.975000 64.380000 194.775000 ;
      RECT 63.580000 195.595000 64.380000 196.395000 ;
      RECT 63.580000 197.215000 64.380000 198.015000 ;
      RECT 63.580000 198.835000 64.380000 199.635000 ;
      RECT 63.585000  37.145000 64.385000  37.945000 ;
      RECT 63.585000  38.975000 64.385000  39.775000 ;
      RECT 63.585000  58.645000 64.385000  59.445000 ;
      RECT 63.585000  61.475000 64.385000  62.275000 ;
      RECT 65.175000   9.295000 65.975000  10.095000 ;
      RECT 65.175000  12.325000 65.975000  13.125000 ;
      RECT 65.175000  20.195000 65.975000  20.995000 ;
      RECT 65.175000  23.225000 65.975000  24.025000 ;
      RECT 65.175000  41.995000 65.975000  42.795000 ;
      RECT 65.175000  45.025000 65.975000  45.825000 ;
      RECT 65.180000   2.450000 65.980000   3.250000 ;
      RECT 65.180000   4.360000 65.980000   5.160000 ;
      RECT 65.180000   6.270000 65.980000   7.070000 ;
      RECT 65.180000  15.345000 65.980000  16.145000 ;
      RECT 65.180000  17.175000 65.980000  17.975000 ;
      RECT 65.180000  26.245000 65.980000  27.045000 ;
      RECT 65.180000  29.275000 65.980000  30.075000 ;
      RECT 65.180000  32.295000 65.980000  33.095000 ;
      RECT 65.180000  34.125000 65.980000  34.925000 ;
      RECT 65.180000  51.835000 65.980000  52.635000 ;
      RECT 65.180000  64.495000 65.980000  65.295000 ;
      RECT 65.180000  67.325000 65.980000  68.125000 ;
      RECT 65.180000  70.350000 65.980000  71.150000 ;
      RECT 65.180000  72.030000 65.980000  72.830000 ;
      RECT 65.180000  73.710000 65.980000  74.510000 ;
      RECT 65.180000  75.390000 65.980000  76.190000 ;
      RECT 65.180000  77.070000 65.980000  77.870000 ;
      RECT 65.180000  78.750000 65.980000  79.550000 ;
      RECT 65.180000  80.430000 65.980000  81.230000 ;
      RECT 65.180000  82.110000 65.980000  82.910000 ;
      RECT 65.180000  83.790000 65.980000  84.590000 ;
      RECT 65.180000  85.470000 65.980000  86.270000 ;
      RECT 65.180000  87.150000 65.980000  87.950000 ;
      RECT 65.180000  88.830000 65.980000  89.630000 ;
      RECT 65.180000  90.510000 65.980000  91.310000 ;
      RECT 65.180000  92.190000 65.980000  92.990000 ;
      RECT 65.180000  93.870000 65.980000  94.670000 ;
      RECT 65.180000 176.155000 65.980000 176.955000 ;
      RECT 65.180000 177.775000 65.980000 178.575000 ;
      RECT 65.180000 179.395000 65.980000 180.195000 ;
      RECT 65.180000 181.015000 65.980000 181.815000 ;
      RECT 65.180000 182.635000 65.980000 183.435000 ;
      RECT 65.180000 184.255000 65.980000 185.055000 ;
      RECT 65.180000 185.875000 65.980000 186.675000 ;
      RECT 65.180000 187.495000 65.980000 188.295000 ;
      RECT 65.180000 189.115000 65.980000 189.915000 ;
      RECT 65.180000 190.735000 65.980000 191.535000 ;
      RECT 65.180000 192.355000 65.980000 193.155000 ;
      RECT 65.180000 193.975000 65.980000 194.775000 ;
      RECT 65.180000 195.595000 65.980000 196.395000 ;
      RECT 65.180000 197.215000 65.980000 198.015000 ;
      RECT 65.180000 198.835000 65.980000 199.635000 ;
      RECT 65.185000  37.145000 65.985000  37.945000 ;
      RECT 65.185000  38.975000 65.985000  39.775000 ;
      RECT 65.185000  58.645000 65.985000  59.445000 ;
      RECT 65.185000  61.475000 65.985000  62.275000 ;
      RECT 66.775000   9.295000 67.575000  10.095000 ;
      RECT 66.775000  12.325000 67.575000  13.125000 ;
      RECT 66.775000  20.195000 67.575000  20.995000 ;
      RECT 66.775000  23.225000 67.575000  24.025000 ;
      RECT 66.775000  41.995000 67.575000  42.795000 ;
      RECT 66.775000  45.025000 67.575000  45.825000 ;
      RECT 66.780000   2.450000 67.580000   3.250000 ;
      RECT 66.780000   4.360000 67.580000   5.160000 ;
      RECT 66.780000   6.270000 67.580000   7.070000 ;
      RECT 66.780000  15.345000 67.580000  16.145000 ;
      RECT 66.780000  17.175000 67.580000  17.975000 ;
      RECT 66.780000  26.245000 67.580000  27.045000 ;
      RECT 66.780000  29.275000 67.580000  30.075000 ;
      RECT 66.780000  32.295000 67.580000  33.095000 ;
      RECT 66.780000  34.125000 67.580000  34.925000 ;
      RECT 66.780000  51.835000 67.580000  52.635000 ;
      RECT 66.780000  64.495000 67.580000  65.295000 ;
      RECT 66.780000  67.325000 67.580000  68.125000 ;
      RECT 66.780000  70.350000 67.580000  71.150000 ;
      RECT 66.780000  72.030000 67.580000  72.830000 ;
      RECT 66.780000  73.710000 67.580000  74.510000 ;
      RECT 66.780000  75.390000 67.580000  76.190000 ;
      RECT 66.780000  77.070000 67.580000  77.870000 ;
      RECT 66.780000  78.750000 67.580000  79.550000 ;
      RECT 66.780000  80.430000 67.580000  81.230000 ;
      RECT 66.780000  82.110000 67.580000  82.910000 ;
      RECT 66.780000  83.790000 67.580000  84.590000 ;
      RECT 66.780000  85.470000 67.580000  86.270000 ;
      RECT 66.780000  87.150000 67.580000  87.950000 ;
      RECT 66.780000  88.830000 67.580000  89.630000 ;
      RECT 66.780000  90.510000 67.580000  91.310000 ;
      RECT 66.780000  92.190000 67.580000  92.990000 ;
      RECT 66.780000  93.870000 67.580000  94.670000 ;
      RECT 66.780000 176.155000 67.580000 176.955000 ;
      RECT 66.780000 177.775000 67.580000 178.575000 ;
      RECT 66.780000 179.395000 67.580000 180.195000 ;
      RECT 66.780000 181.015000 67.580000 181.815000 ;
      RECT 66.780000 182.635000 67.580000 183.435000 ;
      RECT 66.780000 184.255000 67.580000 185.055000 ;
      RECT 66.780000 185.875000 67.580000 186.675000 ;
      RECT 66.780000 187.495000 67.580000 188.295000 ;
      RECT 66.780000 189.115000 67.580000 189.915000 ;
      RECT 66.780000 190.735000 67.580000 191.535000 ;
      RECT 66.780000 192.355000 67.580000 193.155000 ;
      RECT 66.780000 193.975000 67.580000 194.775000 ;
      RECT 66.780000 195.595000 67.580000 196.395000 ;
      RECT 66.780000 197.215000 67.580000 198.015000 ;
      RECT 66.780000 198.835000 67.580000 199.635000 ;
      RECT 66.785000  37.145000 67.585000  37.945000 ;
      RECT 66.785000  38.975000 67.585000  39.775000 ;
      RECT 66.785000  58.645000 67.585000  59.445000 ;
      RECT 66.785000  61.475000 67.585000  62.275000 ;
      RECT 68.375000   9.295000 69.175000  10.095000 ;
      RECT 68.375000  12.325000 69.175000  13.125000 ;
      RECT 68.375000  20.195000 69.175000  20.995000 ;
      RECT 68.375000  23.225000 69.175000  24.025000 ;
      RECT 68.375000  41.995000 69.175000  42.795000 ;
      RECT 68.375000  45.025000 69.175000  45.825000 ;
      RECT 68.380000   2.450000 69.180000   3.250000 ;
      RECT 68.380000   4.360000 69.180000   5.160000 ;
      RECT 68.380000   6.270000 69.180000   7.070000 ;
      RECT 68.380000  15.345000 69.180000  16.145000 ;
      RECT 68.380000  17.175000 69.180000  17.975000 ;
      RECT 68.380000  26.245000 69.180000  27.045000 ;
      RECT 68.380000  29.275000 69.180000  30.075000 ;
      RECT 68.380000  32.295000 69.180000  33.095000 ;
      RECT 68.380000  34.125000 69.180000  34.925000 ;
      RECT 68.380000  51.835000 69.180000  52.635000 ;
      RECT 68.380000  64.495000 69.180000  65.295000 ;
      RECT 68.380000  67.325000 69.180000  68.125000 ;
      RECT 68.380000  70.350000 69.180000  71.150000 ;
      RECT 68.380000  72.030000 69.180000  72.830000 ;
      RECT 68.380000  73.710000 69.180000  74.510000 ;
      RECT 68.380000  75.390000 69.180000  76.190000 ;
      RECT 68.380000  77.070000 69.180000  77.870000 ;
      RECT 68.380000  78.750000 69.180000  79.550000 ;
      RECT 68.380000  80.430000 69.180000  81.230000 ;
      RECT 68.380000  82.110000 69.180000  82.910000 ;
      RECT 68.380000  83.790000 69.180000  84.590000 ;
      RECT 68.380000  85.470000 69.180000  86.270000 ;
      RECT 68.380000  87.150000 69.180000  87.950000 ;
      RECT 68.380000  88.830000 69.180000  89.630000 ;
      RECT 68.380000  90.510000 69.180000  91.310000 ;
      RECT 68.380000  92.190000 69.180000  92.990000 ;
      RECT 68.380000  93.870000 69.180000  94.670000 ;
      RECT 68.380000 176.155000 69.180000 176.955000 ;
      RECT 68.380000 177.775000 69.180000 178.575000 ;
      RECT 68.380000 179.395000 69.180000 180.195000 ;
      RECT 68.380000 181.015000 69.180000 181.815000 ;
      RECT 68.380000 182.635000 69.180000 183.435000 ;
      RECT 68.380000 184.255000 69.180000 185.055000 ;
      RECT 68.380000 185.875000 69.180000 186.675000 ;
      RECT 68.380000 187.495000 69.180000 188.295000 ;
      RECT 68.380000 189.115000 69.180000 189.915000 ;
      RECT 68.380000 190.735000 69.180000 191.535000 ;
      RECT 68.380000 192.355000 69.180000 193.155000 ;
      RECT 68.380000 193.975000 69.180000 194.775000 ;
      RECT 68.380000 195.595000 69.180000 196.395000 ;
      RECT 68.380000 197.215000 69.180000 198.015000 ;
      RECT 68.380000 198.835000 69.180000 199.635000 ;
      RECT 68.385000  37.145000 69.185000  37.945000 ;
      RECT 68.385000  38.975000 69.185000  39.775000 ;
      RECT 68.385000  58.645000 69.185000  59.445000 ;
      RECT 68.385000  61.475000 69.185000  62.275000 ;
      RECT 69.975000   9.295000 70.775000  10.095000 ;
      RECT 69.975000  12.325000 70.775000  13.125000 ;
      RECT 69.975000  20.195000 70.775000  20.995000 ;
      RECT 69.975000  23.225000 70.775000  24.025000 ;
      RECT 69.975000  41.995000 70.775000  42.795000 ;
      RECT 69.975000  45.025000 70.775000  45.825000 ;
      RECT 69.980000   2.450000 70.780000   3.250000 ;
      RECT 69.980000   4.360000 70.780000   5.160000 ;
      RECT 69.980000   6.270000 70.780000   7.070000 ;
      RECT 69.980000  15.345000 70.780000  16.145000 ;
      RECT 69.980000  17.175000 70.780000  17.975000 ;
      RECT 69.980000  26.245000 70.780000  27.045000 ;
      RECT 69.980000  29.275000 70.780000  30.075000 ;
      RECT 69.980000  32.295000 70.780000  33.095000 ;
      RECT 69.980000  34.125000 70.780000  34.925000 ;
      RECT 69.980000  51.835000 70.780000  52.635000 ;
      RECT 69.980000  64.495000 70.780000  65.295000 ;
      RECT 69.980000  67.325000 70.780000  68.125000 ;
      RECT 69.980000  70.350000 70.780000  71.150000 ;
      RECT 69.980000  72.030000 70.780000  72.830000 ;
      RECT 69.980000  73.710000 70.780000  74.510000 ;
      RECT 69.980000  75.390000 70.780000  76.190000 ;
      RECT 69.980000  77.070000 70.780000  77.870000 ;
      RECT 69.980000  78.750000 70.780000  79.550000 ;
      RECT 69.980000  80.430000 70.780000  81.230000 ;
      RECT 69.980000  82.110000 70.780000  82.910000 ;
      RECT 69.980000  83.790000 70.780000  84.590000 ;
      RECT 69.980000  85.470000 70.780000  86.270000 ;
      RECT 69.980000  87.150000 70.780000  87.950000 ;
      RECT 69.980000  88.830000 70.780000  89.630000 ;
      RECT 69.980000  90.510000 70.780000  91.310000 ;
      RECT 69.980000  92.190000 70.780000  92.990000 ;
      RECT 69.980000  93.870000 70.780000  94.670000 ;
      RECT 69.980000 176.155000 70.780000 176.955000 ;
      RECT 69.980000 177.775000 70.780000 178.575000 ;
      RECT 69.980000 179.395000 70.780000 180.195000 ;
      RECT 69.980000 181.015000 70.780000 181.815000 ;
      RECT 69.980000 182.635000 70.780000 183.435000 ;
      RECT 69.980000 184.255000 70.780000 185.055000 ;
      RECT 69.980000 185.875000 70.780000 186.675000 ;
      RECT 69.980000 187.495000 70.780000 188.295000 ;
      RECT 69.980000 189.115000 70.780000 189.915000 ;
      RECT 69.980000 190.735000 70.780000 191.535000 ;
      RECT 69.980000 192.355000 70.780000 193.155000 ;
      RECT 69.980000 193.975000 70.780000 194.775000 ;
      RECT 69.980000 195.595000 70.780000 196.395000 ;
      RECT 69.980000 197.215000 70.780000 198.015000 ;
      RECT 69.980000 198.835000 70.780000 199.635000 ;
      RECT 69.985000  37.145000 70.785000  37.945000 ;
      RECT 69.985000  38.975000 70.785000  39.775000 ;
      RECT 69.985000  58.645000 70.785000  59.445000 ;
      RECT 69.985000  61.475000 70.785000  62.275000 ;
      RECT 71.575000   9.295000 72.375000  10.095000 ;
      RECT 71.575000  12.325000 72.375000  13.125000 ;
      RECT 71.575000  20.195000 72.375000  20.995000 ;
      RECT 71.575000  23.225000 72.375000  24.025000 ;
      RECT 71.575000  41.995000 72.375000  42.795000 ;
      RECT 71.575000  45.025000 72.375000  45.825000 ;
      RECT 71.580000   2.450000 72.380000   3.250000 ;
      RECT 71.580000   4.360000 72.380000   5.160000 ;
      RECT 71.580000   6.270000 72.380000   7.070000 ;
      RECT 71.580000  15.345000 72.380000  16.145000 ;
      RECT 71.580000  17.175000 72.380000  17.975000 ;
      RECT 71.580000  26.245000 72.380000  27.045000 ;
      RECT 71.580000  29.275000 72.380000  30.075000 ;
      RECT 71.580000  32.295000 72.380000  33.095000 ;
      RECT 71.580000  34.125000 72.380000  34.925000 ;
      RECT 71.580000  51.835000 72.380000  52.635000 ;
      RECT 71.580000  64.495000 72.380000  65.295000 ;
      RECT 71.580000  67.325000 72.380000  68.125000 ;
      RECT 71.580000  70.350000 72.380000  71.150000 ;
      RECT 71.580000  72.030000 72.380000  72.830000 ;
      RECT 71.580000  73.710000 72.380000  74.510000 ;
      RECT 71.580000  75.390000 72.380000  76.190000 ;
      RECT 71.580000  77.070000 72.380000  77.870000 ;
      RECT 71.580000  78.750000 72.380000  79.550000 ;
      RECT 71.580000  80.430000 72.380000  81.230000 ;
      RECT 71.580000  82.110000 72.380000  82.910000 ;
      RECT 71.580000  83.790000 72.380000  84.590000 ;
      RECT 71.580000  85.470000 72.380000  86.270000 ;
      RECT 71.580000  87.150000 72.380000  87.950000 ;
      RECT 71.580000  88.830000 72.380000  89.630000 ;
      RECT 71.580000  90.510000 72.380000  91.310000 ;
      RECT 71.580000  92.190000 72.380000  92.990000 ;
      RECT 71.580000  93.870000 72.380000  94.670000 ;
      RECT 71.580000 176.155000 72.380000 176.955000 ;
      RECT 71.580000 177.775000 72.380000 178.575000 ;
      RECT 71.580000 179.395000 72.380000 180.195000 ;
      RECT 71.580000 181.015000 72.380000 181.815000 ;
      RECT 71.580000 182.635000 72.380000 183.435000 ;
      RECT 71.580000 184.255000 72.380000 185.055000 ;
      RECT 71.580000 185.875000 72.380000 186.675000 ;
      RECT 71.580000 187.495000 72.380000 188.295000 ;
      RECT 71.580000 189.115000 72.380000 189.915000 ;
      RECT 71.580000 190.735000 72.380000 191.535000 ;
      RECT 71.580000 192.355000 72.380000 193.155000 ;
      RECT 71.580000 193.975000 72.380000 194.775000 ;
      RECT 71.580000 195.595000 72.380000 196.395000 ;
      RECT 71.580000 197.215000 72.380000 198.015000 ;
      RECT 71.580000 198.835000 72.380000 199.635000 ;
      RECT 71.585000  37.145000 72.385000  37.945000 ;
      RECT 71.585000  38.975000 72.385000  39.775000 ;
      RECT 71.585000  58.645000 72.385000  59.445000 ;
      RECT 71.585000  61.475000 72.385000  62.275000 ;
      RECT 73.175000   9.295000 73.975000  10.095000 ;
      RECT 73.175000  12.325000 73.975000  13.125000 ;
      RECT 73.175000  20.195000 73.975000  20.995000 ;
      RECT 73.175000  23.225000 73.975000  24.025000 ;
      RECT 73.175000  41.995000 73.975000  42.795000 ;
      RECT 73.175000  45.025000 73.975000  45.825000 ;
      RECT 73.180000   2.450000 73.980000   3.250000 ;
      RECT 73.180000   4.360000 73.980000   5.160000 ;
      RECT 73.180000   6.270000 73.980000   7.070000 ;
      RECT 73.180000  15.345000 73.980000  16.145000 ;
      RECT 73.180000  17.175000 73.980000  17.975000 ;
      RECT 73.180000  26.245000 73.980000  27.045000 ;
      RECT 73.180000  29.275000 73.980000  30.075000 ;
      RECT 73.180000  32.295000 73.980000  33.095000 ;
      RECT 73.180000  34.125000 73.980000  34.925000 ;
      RECT 73.180000  51.835000 73.980000  52.635000 ;
      RECT 73.180000  64.495000 73.980000  65.295000 ;
      RECT 73.180000  67.325000 73.980000  68.125000 ;
      RECT 73.180000  70.350000 73.980000  71.150000 ;
      RECT 73.180000  72.030000 73.980000  72.830000 ;
      RECT 73.180000  73.710000 73.980000  74.510000 ;
      RECT 73.180000  75.390000 73.980000  76.190000 ;
      RECT 73.180000  77.070000 73.980000  77.870000 ;
      RECT 73.180000  78.750000 73.980000  79.550000 ;
      RECT 73.180000  80.430000 73.980000  81.230000 ;
      RECT 73.180000  82.110000 73.980000  82.910000 ;
      RECT 73.180000  83.790000 73.980000  84.590000 ;
      RECT 73.180000  85.470000 73.980000  86.270000 ;
      RECT 73.180000  87.150000 73.980000  87.950000 ;
      RECT 73.180000  88.830000 73.980000  89.630000 ;
      RECT 73.180000  90.510000 73.980000  91.310000 ;
      RECT 73.180000  92.190000 73.980000  92.990000 ;
      RECT 73.180000  93.870000 73.980000  94.670000 ;
      RECT 73.180000 176.155000 73.980000 176.955000 ;
      RECT 73.180000 177.775000 73.980000 178.575000 ;
      RECT 73.180000 179.395000 73.980000 180.195000 ;
      RECT 73.180000 181.015000 73.980000 181.815000 ;
      RECT 73.180000 182.635000 73.980000 183.435000 ;
      RECT 73.180000 184.255000 73.980000 185.055000 ;
      RECT 73.180000 185.875000 73.980000 186.675000 ;
      RECT 73.180000 187.495000 73.980000 188.295000 ;
      RECT 73.180000 189.115000 73.980000 189.915000 ;
      RECT 73.180000 190.735000 73.980000 191.535000 ;
      RECT 73.180000 192.355000 73.980000 193.155000 ;
      RECT 73.180000 193.975000 73.980000 194.775000 ;
      RECT 73.180000 195.595000 73.980000 196.395000 ;
      RECT 73.180000 197.215000 73.980000 198.015000 ;
      RECT 73.180000 198.835000 73.980000 199.635000 ;
      RECT 73.185000  37.145000 73.985000  37.945000 ;
      RECT 73.185000  38.975000 73.985000  39.775000 ;
      RECT 73.185000  58.645000 73.985000  59.445000 ;
      RECT 73.185000  61.475000 73.985000  62.275000 ;
      RECT 74.775000   9.295000 75.575000  10.095000 ;
      RECT 74.775000  12.325000 75.575000  13.125000 ;
      RECT 74.775000  20.195000 75.575000  20.995000 ;
      RECT 74.775000  23.225000 75.575000  24.025000 ;
      RECT 74.775000  41.995000 75.575000  42.795000 ;
      RECT 74.775000  45.025000 75.575000  45.825000 ;
      RECT 74.780000   2.450000 75.580000   3.250000 ;
      RECT 74.780000   4.360000 75.580000   5.160000 ;
      RECT 74.780000   6.270000 75.580000   7.070000 ;
      RECT 74.780000  15.345000 75.580000  16.145000 ;
      RECT 74.780000  17.175000 75.580000  17.975000 ;
      RECT 74.780000  26.245000 75.580000  27.045000 ;
      RECT 74.780000  29.275000 75.580000  30.075000 ;
      RECT 74.780000  32.295000 75.580000  33.095000 ;
      RECT 74.780000  34.125000 75.580000  34.925000 ;
      RECT 74.780000  51.835000 75.580000  52.635000 ;
      RECT 74.780000  64.495000 75.580000  65.295000 ;
      RECT 74.780000  67.325000 75.580000  68.125000 ;
      RECT 74.780000  70.350000 75.580000  71.150000 ;
      RECT 74.780000  72.030000 75.580000  72.830000 ;
      RECT 74.780000  73.710000 75.580000  74.510000 ;
      RECT 74.780000  75.390000 75.580000  76.190000 ;
      RECT 74.780000  77.070000 75.580000  77.870000 ;
      RECT 74.780000  78.750000 75.580000  79.550000 ;
      RECT 74.780000  80.430000 75.580000  81.230000 ;
      RECT 74.780000  82.110000 75.580000  82.910000 ;
      RECT 74.780000  83.790000 75.580000  84.590000 ;
      RECT 74.780000  85.470000 75.580000  86.270000 ;
      RECT 74.780000  87.150000 75.580000  87.950000 ;
      RECT 74.780000  88.830000 75.580000  89.630000 ;
      RECT 74.780000  90.510000 75.580000  91.310000 ;
      RECT 74.780000  92.190000 75.580000  92.990000 ;
      RECT 74.780000  93.870000 75.580000  94.670000 ;
      RECT 74.780000 176.155000 75.580000 176.955000 ;
      RECT 74.780000 177.775000 75.580000 178.575000 ;
      RECT 74.780000 179.395000 75.580000 180.195000 ;
      RECT 74.780000 181.015000 75.580000 181.815000 ;
      RECT 74.780000 182.635000 75.580000 183.435000 ;
      RECT 74.780000 184.255000 75.580000 185.055000 ;
      RECT 74.780000 185.875000 75.580000 186.675000 ;
      RECT 74.780000 187.495000 75.580000 188.295000 ;
      RECT 74.780000 189.115000 75.580000 189.915000 ;
      RECT 74.780000 190.735000 75.580000 191.535000 ;
      RECT 74.780000 192.355000 75.580000 193.155000 ;
      RECT 74.780000 193.975000 75.580000 194.775000 ;
      RECT 74.780000 195.595000 75.580000 196.395000 ;
      RECT 74.780000 197.215000 75.580000 198.015000 ;
      RECT 74.780000 198.835000 75.580000 199.635000 ;
      RECT 74.785000  37.145000 75.585000  37.945000 ;
      RECT 74.785000  38.975000 75.585000  39.775000 ;
      RECT 74.785000  58.645000 75.585000  59.445000 ;
      RECT 74.785000  61.475000 75.585000  62.275000 ;
      RECT 76.375000   9.295000 77.175000  10.095000 ;
      RECT 76.375000  12.325000 77.175000  13.125000 ;
      RECT 76.375000  20.195000 77.175000  20.995000 ;
      RECT 76.375000  23.225000 77.175000  24.025000 ;
      RECT 76.375000  41.995000 77.175000  42.795000 ;
      RECT 76.375000  45.025000 77.175000  45.825000 ;
      RECT 76.380000   2.450000 77.180000   3.250000 ;
      RECT 76.380000   4.360000 77.180000   5.160000 ;
      RECT 76.380000   6.270000 77.180000   7.070000 ;
      RECT 76.380000  15.345000 77.180000  16.145000 ;
      RECT 76.380000  17.175000 77.180000  17.975000 ;
      RECT 76.380000  26.245000 77.180000  27.045000 ;
      RECT 76.380000  29.275000 77.180000  30.075000 ;
      RECT 76.380000  32.295000 77.180000  33.095000 ;
      RECT 76.380000  34.125000 77.180000  34.925000 ;
      RECT 76.380000  51.835000 77.180000  52.635000 ;
      RECT 76.380000  64.495000 77.180000  65.295000 ;
      RECT 76.380000  67.325000 77.180000  68.125000 ;
      RECT 76.380000  70.350000 77.180000  71.150000 ;
      RECT 76.380000  72.030000 77.180000  72.830000 ;
      RECT 76.380000  73.710000 77.180000  74.510000 ;
      RECT 76.380000  75.390000 77.180000  76.190000 ;
      RECT 76.380000  77.070000 77.180000  77.870000 ;
      RECT 76.380000  78.750000 77.180000  79.550000 ;
      RECT 76.380000  80.430000 77.180000  81.230000 ;
      RECT 76.380000  82.110000 77.180000  82.910000 ;
      RECT 76.380000  83.790000 77.180000  84.590000 ;
      RECT 76.380000  85.470000 77.180000  86.270000 ;
      RECT 76.380000  87.150000 77.180000  87.950000 ;
      RECT 76.380000  88.830000 77.180000  89.630000 ;
      RECT 76.380000  90.510000 77.180000  91.310000 ;
      RECT 76.380000  92.190000 77.180000  92.990000 ;
      RECT 76.380000  93.870000 77.180000  94.670000 ;
      RECT 76.380000 176.155000 77.180000 176.955000 ;
      RECT 76.380000 177.775000 77.180000 178.575000 ;
      RECT 76.380000 179.395000 77.180000 180.195000 ;
      RECT 76.380000 181.015000 77.180000 181.815000 ;
      RECT 76.380000 182.635000 77.180000 183.435000 ;
      RECT 76.380000 184.255000 77.180000 185.055000 ;
      RECT 76.380000 185.875000 77.180000 186.675000 ;
      RECT 76.380000 187.495000 77.180000 188.295000 ;
      RECT 76.380000 189.115000 77.180000 189.915000 ;
      RECT 76.380000 190.735000 77.180000 191.535000 ;
      RECT 76.380000 192.355000 77.180000 193.155000 ;
      RECT 76.380000 193.975000 77.180000 194.775000 ;
      RECT 76.380000 195.595000 77.180000 196.395000 ;
      RECT 76.380000 197.215000 77.180000 198.015000 ;
      RECT 76.380000 198.835000 77.180000 199.635000 ;
      RECT 76.385000  37.145000 77.185000  37.945000 ;
      RECT 76.385000  38.975000 77.185000  39.775000 ;
      RECT 76.385000  58.645000 77.185000  59.445000 ;
      RECT 76.385000  61.475000 77.185000  62.275000 ;
      RECT 77.975000   9.295000 78.775000  10.095000 ;
      RECT 77.975000  12.325000 78.775000  13.125000 ;
      RECT 77.975000  20.195000 78.775000  20.995000 ;
      RECT 77.975000  23.225000 78.775000  24.025000 ;
      RECT 77.975000  41.995000 78.775000  42.795000 ;
      RECT 77.975000  45.025000 78.775000  45.825000 ;
      RECT 77.980000   2.450000 78.780000   3.250000 ;
      RECT 77.980000   4.360000 78.780000   5.160000 ;
      RECT 77.980000   6.270000 78.780000   7.070000 ;
      RECT 77.980000  15.345000 78.780000  16.145000 ;
      RECT 77.980000  17.175000 78.780000  17.975000 ;
      RECT 77.980000  26.245000 78.780000  27.045000 ;
      RECT 77.980000  29.275000 78.780000  30.075000 ;
      RECT 77.980000  32.295000 78.780000  33.095000 ;
      RECT 77.980000  34.125000 78.780000  34.925000 ;
      RECT 77.980000  51.835000 78.780000  52.635000 ;
      RECT 77.980000  64.495000 78.780000  65.295000 ;
      RECT 77.980000  67.325000 78.780000  68.125000 ;
      RECT 77.980000  70.350000 78.780000  71.150000 ;
      RECT 77.980000  72.030000 78.780000  72.830000 ;
      RECT 77.980000  73.710000 78.780000  74.510000 ;
      RECT 77.980000  75.390000 78.780000  76.190000 ;
      RECT 77.980000  77.070000 78.780000  77.870000 ;
      RECT 77.980000  78.750000 78.780000  79.550000 ;
      RECT 77.980000  80.430000 78.780000  81.230000 ;
      RECT 77.980000  82.110000 78.780000  82.910000 ;
      RECT 77.980000  83.790000 78.780000  84.590000 ;
      RECT 77.980000  85.470000 78.780000  86.270000 ;
      RECT 77.980000  87.150000 78.780000  87.950000 ;
      RECT 77.980000  88.830000 78.780000  89.630000 ;
      RECT 77.980000  90.510000 78.780000  91.310000 ;
      RECT 77.980000  92.190000 78.780000  92.990000 ;
      RECT 77.980000  93.870000 78.780000  94.670000 ;
      RECT 77.980000 176.155000 78.780000 176.955000 ;
      RECT 77.980000 177.775000 78.780000 178.575000 ;
      RECT 77.980000 179.395000 78.780000 180.195000 ;
      RECT 77.980000 181.015000 78.780000 181.815000 ;
      RECT 77.980000 182.635000 78.780000 183.435000 ;
      RECT 77.980000 184.255000 78.780000 185.055000 ;
      RECT 77.980000 185.875000 78.780000 186.675000 ;
      RECT 77.980000 187.495000 78.780000 188.295000 ;
      RECT 77.980000 189.115000 78.780000 189.915000 ;
      RECT 77.980000 190.735000 78.780000 191.535000 ;
      RECT 77.980000 192.355000 78.780000 193.155000 ;
      RECT 77.980000 193.975000 78.780000 194.775000 ;
      RECT 77.980000 195.595000 78.780000 196.395000 ;
      RECT 77.980000 197.215000 78.780000 198.015000 ;
      RECT 77.980000 198.835000 78.780000 199.635000 ;
      RECT 77.985000  37.145000 78.785000  37.945000 ;
      RECT 77.985000  38.975000 78.785000  39.775000 ;
      RECT 77.985000  58.645000 78.785000  59.445000 ;
      RECT 77.985000  61.475000 78.785000  62.275000 ;
  END
END sky130_fd_io__overlay_gpiov2


MACRO sky130_fd_io__top_xres4v2
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN DISABLE_PULLUP_H
    ANTENNAPARTIALCUTAREA  0.045000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 28.635000 28.540000 33.025000 28.580000 ;
        RECT 28.635000 28.580000 28.950000 28.650000 ;
        RECT 28.635000 28.650000 28.880000 28.720000 ;
        RECT 28.635000 28.720000 28.865000 28.735000 ;
        RECT 28.635000 28.735000 28.865000 32.435000 ;
        RECT 28.685000 28.490000 33.025000 28.540000 ;
        RECT 28.755000 28.420000 33.025000 28.490000 ;
        RECT 28.825000 28.350000 33.025000 28.420000 ;
        RECT 32.555000 28.340000 33.025000 28.350000 ;
        RECT 32.625000 28.270000 33.025000 28.340000 ;
        RECT 32.695000 28.200000 33.025000 28.270000 ;
        RECT 32.760000  0.000000 33.020000  8.720000 ;
        RECT 32.760000  8.720000 33.020000  8.725000 ;
        RECT 32.760000  8.725000 33.025000  8.830000 ;
        RECT 32.765000  8.830000 33.025000  8.835000 ;
        RECT 32.765000  8.835000 33.025000 28.130000 ;
        RECT 32.765000 28.130000 33.025000 28.200000 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.760000 0.000000 33.020000 0.640000 ;
    END
  END DISABLE_PULLUP_H
  PIN ENABLE_H
    ANTENNAPARTIALCUTAREA  0.180000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 12.145000  6.635000 12.545000  6.665000 ;
        RECT 12.215000  6.565000 12.545000  6.635000 ;
        RECT 12.285000  0.000000 12.545000  6.495000 ;
        RECT 12.285000  6.495000 12.545000  6.565000 ;
        RECT 12.370000  6.665000 12.545000  6.775000 ;
        RECT 12.370000  6.775000 12.545000  6.845000 ;
        RECT 12.370000  6.845000 12.615000  6.915000 ;
        RECT 12.370000  6.915000 12.685000  6.925000 ;
        RECT 12.440000  6.925000 12.695000  6.995000 ;
        RECT 12.510000  6.995000 12.765000  7.065000 ;
        RECT 12.575000  7.065000 12.835000  7.130000 ;
        RECT 12.635000  7.130000 12.900000  7.190000 ;
        RECT 12.695000  7.190000 12.900000  7.250000 ;
        RECT 12.695000  7.250000 12.900000 10.230000 ;
        RECT 12.800000 10.230000 12.865000 10.265000 ;
        RECT 12.800000 10.265000 12.830000 10.300000 ;
        RECT 12.800000 10.300000 12.825000 10.305000 ;
    END
    PORT
      LAYER met2 ;
        RECT 12.285000 0.000000 12.545000 1.470000 ;
    END
  END ENABLE_H
  PIN ENABLE_VDDIO
    ANTENNAPARTIALCUTAREA  0.200000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.425000 0.000000 8.895000 1.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775000 17.410000  7.400000 17.515000 ;
        RECT 6.775000 17.515000  7.295000 17.620000 ;
        RECT 6.775000 17.620000  7.295000 31.295000 ;
        RECT 6.775000 31.295000  7.295000 31.400000 ;
        RECT 6.775000 31.400000  7.400000 31.505000 ;
        RECT 6.840000 17.345000  7.505000 17.410000 ;
        RECT 6.925000 31.505000  7.505000 31.655000 ;
        RECT 6.990000 17.195000  7.570000 17.345000 ;
        RECT 7.075000 31.655000  7.655000 31.805000 ;
        RECT 7.140000 17.045000  7.720000 17.195000 ;
        RECT 7.225000 31.805000  7.805000 31.955000 ;
        RECT 7.290000 16.895000  7.870000 17.045000 ;
        RECT 7.375000 31.955000  7.955000 32.105000 ;
        RECT 7.440000 16.745000  8.020000 16.895000 ;
        RECT 7.525000 32.105000  8.105000 32.255000 ;
        RECT 7.590000 16.595000  8.170000 16.745000 ;
        RECT 7.675000 32.255000  8.255000 32.405000 ;
        RECT 7.740000 16.445000  8.320000 16.595000 ;
        RECT 7.825000 32.405000  8.405000 32.555000 ;
        RECT 7.890000 16.295000  8.470000 16.445000 ;
        RECT 7.975000 32.555000  8.555000 32.705000 ;
        RECT 8.040000 16.145000  8.620000 16.295000 ;
        RECT 8.125000 32.705000  8.705000 32.855000 ;
        RECT 8.190000 15.995000  8.770000 16.145000 ;
        RECT 8.275000 32.855000  8.855000 33.005000 ;
        RECT 8.295000 15.890000  8.920000 15.995000 ;
        RECT 8.400000  0.000000  8.920000 15.785000 ;
        RECT 8.400000 15.785000  8.920000 15.890000 ;
        RECT 8.425000 33.005000  9.005000 33.155000 ;
        RECT 8.575000 33.155000  9.155000 33.305000 ;
        RECT 8.665000 33.305000  9.305000 33.395000 ;
        RECT 8.815000 33.395000 22.275000 33.545000 ;
        RECT 8.965000 33.545000 22.275000 33.695000 ;
        RECT 9.115000 33.695000 22.275000 33.845000 ;
        RECT 9.265000 33.845000 22.275000 33.995000 ;
        RECT 9.395000 33.995000 22.275000 34.125000 ;
    END
  END ENABLE_VDDIO
  PIN EN_VDDIO_SIG_H
    ANTENNAPARTIALCUTAREA  0.157500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 22.360000 0.000000 22.660000 1.205000 ;
    END
    PORT
      LAYER met2 ;
        RECT  9.735000  4.520000 10.050000  4.575000 ;
        RECT  9.735000  4.575000  9.995000  4.630000 ;
        RECT  9.735000  4.630000  9.995000  8.860000 ;
        RECT  9.735000  8.860000  9.995000  8.915000 ;
        RECT  9.735000  8.915000 10.050000  8.970000 ;
        RECT  9.790000  4.465000 10.105000  4.520000 ;
        RECT  9.805000  8.970000 10.105000  9.040000 ;
        RECT  9.860000  4.395000 10.160000  4.465000 ;
        RECT  9.875000  9.040000 10.175000  9.110000 ;
        RECT  9.930000  4.325000 10.230000  4.395000 ;
        RECT  9.945000  9.110000 10.245000  9.180000 ;
        RECT 10.000000  4.255000 10.300000  4.325000 ;
        RECT 10.015000  9.180000 10.315000  9.250000 ;
        RECT 10.070000  4.185000 10.370000  4.255000 ;
        RECT 10.085000  9.250000 10.385000  9.320000 ;
        RECT 10.140000  4.115000 10.440000  4.185000 ;
        RECT 10.155000  9.320000 10.455000  9.390000 ;
        RECT 10.210000  4.045000 10.510000  4.115000 ;
        RECT 10.225000  9.390000 10.525000  9.460000 ;
        RECT 10.280000  3.975000 10.580000  4.045000 ;
        RECT 10.295000  9.460000 10.595000  9.530000 ;
        RECT 10.350000  3.905000 10.650000  3.975000 ;
        RECT 10.365000  9.530000 10.665000  9.600000 ;
        RECT 10.420000  3.835000 10.720000  3.905000 ;
        RECT 10.435000  9.600000 10.735000  9.670000 ;
        RECT 10.490000  3.765000 10.790000  3.835000 ;
        RECT 10.505000  9.670000 10.805000  9.740000 ;
        RECT 10.560000  3.695000 10.860000  3.765000 ;
        RECT 10.575000  9.740000 10.875000  9.810000 ;
        RECT 10.610000  3.645000 15.095000  3.695000 ;
        RECT 10.645000  9.810000 10.945000  9.880000 ;
        RECT 10.650000 26.825000 11.125000 27.085000 ;
        RECT 10.650000 27.085000 11.055000 27.155000 ;
        RECT 10.650000 27.155000 10.985000 27.225000 ;
        RECT 10.650000 27.225000 10.915000 27.295000 ;
        RECT 10.650000 27.295000 10.910000 27.300000 ;
        RECT 10.650000 27.300000 10.910000 27.935000 ;
        RECT 10.650000 27.935000 10.910000 28.005000 ;
        RECT 10.650000 28.005000 10.980000 28.075000 ;
        RECT 10.650000 28.075000 11.050000 28.145000 ;
        RECT 10.650000 28.145000 11.120000 28.150000 ;
        RECT 10.650000 28.150000 11.125000 28.410000 ;
        RECT 10.655000 26.820000 11.125000 26.825000 ;
        RECT 10.680000  3.575000 15.025000  3.645000 ;
        RECT 10.715000  9.880000 11.015000  9.950000 ;
        RECT 10.720000 28.410000 11.125000 28.480000 ;
        RECT 10.725000 26.750000 11.125000 26.820000 ;
        RECT 10.750000  3.505000 14.955000  3.575000 ;
        RECT 10.755000  9.950000 11.085000  9.990000 ;
        RECT 10.790000 28.480000 11.125000 28.550000 ;
        RECT 10.795000 26.680000 11.125000 26.750000 ;
        RECT 10.810000  9.990000 11.125000 10.045000 ;
        RECT 10.820000  3.435000 14.885000  3.505000 ;
        RECT 10.860000 28.550000 11.125000 28.620000 ;
        RECT 10.865000 10.045000 11.125000 10.100000 ;
        RECT 10.865000 10.100000 11.125000 26.610000 ;
        RECT 10.865000 26.610000 11.125000 26.680000 ;
        RECT 10.865000 28.620000 11.125000 28.625000 ;
        RECT 10.865000 28.625000 11.125000 31.085000 ;
        RECT 10.865000 31.085000 11.125000 31.140000 ;
        RECT 10.865000 31.140000 11.180000 31.195000 ;
        RECT 10.935000 31.195000 11.235000 31.265000 ;
        RECT 11.005000 31.265000 11.305000 31.335000 ;
        RECT 11.075000 31.335000 11.375000 31.405000 ;
        RECT 11.145000 31.405000 11.445000 31.475000 ;
        RECT 11.150000 31.475000 11.515000 31.480000 ;
        RECT 11.205000 31.480000 11.520000 31.535000 ;
        RECT 11.260000 31.535000 11.520000 31.590000 ;
        RECT 11.260000 31.590000 11.520000 36.020000 ;
        RECT 11.260000 36.020000 12.150000 36.280000 ;
        RECT 14.845000  3.695000 15.145000  3.765000 ;
        RECT 14.915000  3.765000 15.215000  3.835000 ;
        RECT 14.985000  3.835000 15.285000  3.905000 ;
        RECT 15.055000  3.905000 15.355000  3.975000 ;
        RECT 15.125000  3.975000 15.425000  4.045000 ;
        RECT 15.195000  4.045000 15.495000  4.115000 ;
        RECT 15.265000  4.115000 15.565000  4.185000 ;
        RECT 15.335000  4.185000 15.635000  4.255000 ;
        RECT 15.405000  4.255000 15.705000  4.325000 ;
        RECT 15.475000  4.325000 15.775000  4.395000 ;
        RECT 15.545000  4.395000 15.845000  4.465000 ;
        RECT 15.615000  4.465000 15.915000  4.535000 ;
        RECT 15.625000  4.535000 15.985000  4.545000 ;
        RECT 15.695000  4.545000 28.765000  4.615000 ;
        RECT 15.765000  4.615000 28.835000  4.685000 ;
        RECT 15.835000  4.685000 28.905000  4.755000 ;
        RECT 15.885000  4.755000 28.975000  4.805000 ;
        RECT 22.065000  4.540000 22.940000  4.545000 ;
        RECT 22.135000  4.470000 22.870000  4.540000 ;
        RECT 22.205000  4.400000 22.800000  4.470000 ;
        RECT 22.275000  4.330000 22.730000  4.400000 ;
        RECT 22.345000  4.260000 22.660000  4.330000 ;
        RECT 22.350000  4.255000 22.660000  4.260000 ;
        RECT 22.355000  4.250000 22.660000  4.255000 ;
        RECT 22.360000  0.000000 22.660000  4.245000 ;
        RECT 22.360000  4.245000 22.660000  4.250000 ;
        RECT 28.725000  4.805000 29.025000  4.875000 ;
        RECT 28.795000  4.875000 29.095000  4.945000 ;
        RECT 28.865000  4.945000 29.165000  5.015000 ;
        RECT 28.935000  5.015000 29.235000  5.085000 ;
        RECT 29.005000  5.085000 29.305000  5.155000 ;
        RECT 29.075000  5.155000 29.375000  5.225000 ;
        RECT 29.145000  5.225000 29.445000  5.295000 ;
        RECT 29.210000  5.295000 29.515000  5.360000 ;
        RECT 29.265000  5.360000 29.580000  5.415000 ;
        RECT 29.320000  5.415000 29.580000  5.470000 ;
        RECT 29.320000  5.470000 29.580000 10.975000 ;
        RECT 29.320000 10.975000 29.580000 11.030000 ;
        RECT 29.320000 11.030000 29.635000 11.085000 ;
        RECT 29.390000 11.085000 29.690000 11.155000 ;
        RECT 29.460000 11.155000 29.760000 11.225000 ;
        RECT 29.530000 11.225000 29.830000 11.295000 ;
        RECT 29.600000 11.295000 29.900000 11.365000 ;
        RECT 29.660000 11.365000 29.970000 11.425000 ;
        RECT 29.715000 11.425000 30.030000 11.480000 ;
        RECT 29.770000 11.480000 30.030000 11.535000 ;
        RECT 29.770000 11.535000 30.030000 15.645000 ;
        RECT 29.770000 15.645000 30.030000 15.700000 ;
        RECT 29.770000 15.700000 30.085000 15.755000 ;
        RECT 29.840000 15.755000 30.140000 15.825000 ;
        RECT 29.910000 15.825000 30.210000 15.895000 ;
        RECT 29.980000 15.895000 30.280000 15.965000 ;
        RECT 30.050000 15.965000 30.350000 16.035000 ;
        RECT 30.120000 16.035000 30.420000 16.105000 ;
        RECT 30.190000 16.105000 30.490000 16.175000 ;
        RECT 30.255000 16.175000 30.560000 16.240000 ;
        RECT 30.310000 16.240000 30.625000 16.295000 ;
        RECT 30.365000 16.295000 30.625000 16.350000 ;
        RECT 30.365000 16.350000 30.625000 20.495000 ;
    END
  END EN_VDDIO_SIG_H
  PIN FILT_IN_H
    ANTENNAPARTIALCUTAREA  0.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.075000 0.000000 21.225000 3.455000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075000 0.000000 21.225000  6.670000 ;
        RECT 20.075000 6.670000 21.225000  6.820000 ;
        RECT 20.075000 6.820000 21.375000  6.970000 ;
        RECT 20.075000 6.970000 21.525000  7.120000 ;
        RECT 20.075000 7.120000 21.675000  7.150000 ;
        RECT 20.225000 7.150000 21.705000  7.300000 ;
        RECT 20.375000 7.300000 21.855000  7.450000 ;
        RECT 20.525000 7.450000 22.005000  7.600000 ;
        RECT 20.675000 7.600000 22.155000  7.750000 ;
        RECT 20.825000 7.750000 22.305000  7.900000 ;
        RECT 20.975000 7.900000 22.455000  8.050000 ;
        RECT 21.125000 8.050000 22.605000  8.200000 ;
        RECT 21.275000 8.200000 22.755000  8.350000 ;
        RECT 21.425000 8.350000 22.905000  8.500000 ;
        RECT 21.575000 8.500000 23.055000  8.650000 ;
        RECT 21.725000 8.650000 23.205000  8.800000 ;
        RECT 21.875000 8.800000 23.355000  8.950000 ;
        RECT 22.025000 8.950000 23.505000  9.100000 ;
        RECT 22.175000 9.100000 23.655000  9.250000 ;
        RECT 22.325000 9.250000 23.805000  9.400000 ;
        RECT 22.420000 9.400000 23.955000  9.495000 ;
        RECT 22.570000 9.495000 24.050000  9.645000 ;
        RECT 22.720000 9.645000 24.050000  9.795000 ;
        RECT 22.870000 9.795000 24.050000  9.945000 ;
        RECT 22.905000 9.945000 24.050000  9.980000 ;
        RECT 22.905000 9.980000 24.050000 12.265000 ;
    END
  END FILT_IN_H
  PIN INP_SEL_H
    ANTENNAGATEAREA  6.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.600000 11.420000 16.830000 12.310000 ;
        RECT 16.600000 12.310000 16.830000 12.360000 ;
        RECT 16.600000 12.360000 16.880000 12.410000 ;
        RECT 16.670000 12.410000 16.930000 12.480000 ;
        RECT 16.740000 12.480000 17.000000 12.550000 ;
        RECT 16.810000 12.550000 17.070000 12.620000 ;
        RECT 16.825000 12.620000 17.140000 12.635000 ;
        RECT 16.870000 12.635000 25.295000 12.680000 ;
        RECT 16.915000 12.680000 25.340000 12.725000 ;
        RECT 16.985000 12.725000 25.385000 12.795000 ;
        RECT 17.055000 12.795000 25.385000 12.865000 ;
        RECT 24.640000 12.615000 25.275000 12.635000 ;
        RECT 24.710000 12.545000 25.205000 12.615000 ;
        RECT 24.780000 12.475000 25.135000 12.545000 ;
        RECT 24.785000 12.470000 25.135000 12.475000 ;
        RECT 24.845000 12.410000 25.135000 12.470000 ;
        RECT 24.905000  0.000000 25.135000 12.350000 ;
        RECT 24.905000 12.350000 25.135000 12.410000 ;
        RECT 24.975000 12.865000 25.385000 12.935000 ;
        RECT 25.045000 12.935000 25.385000 13.005000 ;
        RECT 25.115000 13.005000 25.385000 13.075000 ;
        RECT 25.155000 13.075000 25.385000 13.115000 ;
        RECT 25.155000 13.115000 25.385000 15.035000 ;
        RECT 25.155000 15.035000 25.385000 15.085000 ;
        RECT 25.155000 15.085000 25.435000 15.135000 ;
        RECT 25.225000 15.135000 25.485000 15.205000 ;
        RECT 25.295000 15.205000 25.555000 15.275000 ;
        RECT 25.365000 15.275000 25.625000 15.345000 ;
        RECT 25.435000 15.345000 25.695000 15.415000 ;
        RECT 25.505000 15.415000 25.765000 15.485000 ;
        RECT 25.575000 15.485000 25.835000 15.555000 ;
        RECT 25.635000 15.555000 25.905000 15.615000 ;
        RECT 25.705000 15.615000 29.965000 15.685000 ;
        RECT 25.775000 15.685000 30.035000 15.755000 ;
        RECT 25.845000 15.755000 30.105000 15.825000 ;
        RECT 25.865000 15.825000 30.175000 15.845000 ;
        RECT 29.935000 15.845000 30.195000 15.915000 ;
        RECT 30.005000 15.915000 30.265000 15.985000 ;
        RECT 30.075000 15.985000 30.335000 16.055000 ;
        RECT 30.145000 16.055000 30.405000 16.125000 ;
        RECT 30.215000 16.125000 30.475000 16.195000 ;
        RECT 30.285000 16.195000 30.545000 16.265000 ;
        RECT 30.355000 16.265000 30.615000 16.335000 ;
        RECT 30.425000 16.335000 30.685000 16.405000 ;
        RECT 30.495000 16.405000 30.755000 16.475000 ;
        RECT 30.565000 16.475000 30.825000 16.545000 ;
        RECT 30.635000 16.545000 30.895000 16.615000 ;
        RECT 30.705000 16.615000 30.965000 16.685000 ;
        RECT 30.755000 16.685000 31.035000 16.735000 ;
        RECT 30.805000 16.735000 31.035000 16.785000 ;
        RECT 30.805000 16.785000 31.035000 19.345000 ;
    END
  END INP_SEL_H
  PIN PAD
    ANTENNAPARTIALMETALSIDEAREA  245.6270 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 29.695000 127.115000 41.990000 145.625000 ;
    END
  END PAD
  PIN PAD_A_ESD_H
    ANTENNAPARTIALCUTAREA  0.960000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.245000 0.000000 18.910000 3.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.245000 0.000000 18.910000 3.135000 ;
    END
  END PAD_A_ESD_H
  PIN PULLUP_H
    ANTENNAPARTIALCUTAREA  0.270000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  6.065000 43.285000 24.570000 43.355000 ;
        RECT  6.065000 43.355000 24.500000 43.425000 ;
        RECT  6.065000 43.425000 24.430000 43.495000 ;
        RECT  6.065000 43.495000 24.380000 43.545000 ;
        RECT 14.555000  0.000000 15.135000 12.210000 ;
        RECT 14.555000 12.210000 15.135000 12.275000 ;
        RECT 14.555000 12.275000 15.200000 12.340000 ;
        RECT 14.625000 12.340000 15.265000 12.410000 ;
        RECT 14.695000 12.410000 15.335000 12.480000 ;
        RECT 14.765000 12.480000 15.405000 12.550000 ;
        RECT 14.835000 12.550000 15.475000 12.620000 ;
        RECT 14.905000 12.620000 15.545000 12.690000 ;
        RECT 14.975000 12.690000 15.615000 12.760000 ;
        RECT 15.045000 12.760000 15.685000 12.830000 ;
        RECT 15.115000 12.830000 15.755000 12.900000 ;
        RECT 15.185000 12.900000 15.825000 12.970000 ;
        RECT 15.255000 12.970000 15.895000 13.040000 ;
        RECT 15.325000 13.040000 15.965000 13.110000 ;
        RECT 15.395000 13.110000 16.035000 13.180000 ;
        RECT 15.465000 13.180000 16.105000 13.250000 ;
        RECT 15.535000 13.250000 16.175000 13.320000 ;
        RECT 15.605000 13.320000 16.245000 13.390000 ;
        RECT 15.675000 13.390000 16.315000 13.460000 ;
        RECT 15.745000 13.460000 16.385000 13.530000 ;
        RECT 15.815000 13.530000 16.455000 13.600000 ;
        RECT 15.885000 13.600000 16.525000 13.670000 ;
        RECT 15.955000 13.670000 16.595000 13.740000 ;
        RECT 16.025000 13.740000 16.665000 13.810000 ;
        RECT 16.095000 13.810000 16.735000 13.880000 ;
        RECT 16.165000 13.880000 16.805000 13.950000 ;
        RECT 16.235000 13.950000 16.875000 14.020000 ;
        RECT 16.305000 14.020000 16.945000 14.090000 ;
        RECT 16.375000 14.090000 17.015000 14.160000 ;
        RECT 16.445000 14.160000 17.085000 14.230000 ;
        RECT 16.515000 14.230000 17.155000 14.300000 ;
        RECT 16.585000 14.300000 17.225000 14.370000 ;
        RECT 16.655000 14.370000 17.295000 14.440000 ;
        RECT 16.725000 14.440000 17.365000 14.510000 ;
        RECT 16.795000 14.510000 17.435000 14.580000 ;
        RECT 16.865000 14.580000 17.505000 14.650000 ;
        RECT 16.935000 14.650000 17.575000 14.720000 ;
        RECT 17.005000 14.720000 17.645000 14.790000 ;
        RECT 17.075000 14.790000 17.715000 14.860000 ;
        RECT 17.145000 14.860000 17.785000 14.930000 ;
        RECT 17.215000 14.930000 17.855000 15.000000 ;
        RECT 17.285000 15.000000 17.925000 15.070000 ;
        RECT 17.355000 15.070000 17.995000 15.140000 ;
        RECT 17.425000 15.140000 18.065000 15.210000 ;
        RECT 17.495000 15.210000 18.135000 15.280000 ;
        RECT 17.565000 15.280000 18.205000 15.350000 ;
        RECT 17.635000 15.350000 18.275000 15.420000 ;
        RECT 17.705000 15.420000 21.745000 15.490000 ;
        RECT 17.775000 15.490000 21.815000 15.560000 ;
        RECT 17.845000 15.560000 21.885000 15.630000 ;
        RECT 17.915000 15.630000 21.955000 15.700000 ;
        RECT 17.985000 15.700000 22.025000 15.770000 ;
        RECT 18.055000 15.770000 22.095000 15.840000 ;
        RECT 18.125000 15.840000 22.165000 15.910000 ;
        RECT 18.135000 15.910000 22.235000 15.920000 ;
        RECT 21.605000 15.920000 22.245000 15.990000 ;
        RECT 21.675000 15.990000 22.315000 16.060000 ;
        RECT 21.745000 16.060000 22.385000 16.130000 ;
        RECT 21.815000 16.130000 22.455000 16.200000 ;
        RECT 21.885000 16.200000 22.525000 16.270000 ;
        RECT 21.955000 16.270000 22.595000 16.340000 ;
        RECT 22.025000 16.340000 22.665000 16.410000 ;
        RECT 22.095000 16.410000 22.735000 16.480000 ;
        RECT 22.165000 16.480000 22.805000 16.550000 ;
        RECT 22.235000 16.550000 22.875000 16.620000 ;
        RECT 22.305000 16.620000 22.945000 16.690000 ;
        RECT 22.375000 16.690000 23.015000 16.760000 ;
        RECT 22.445000 16.760000 23.085000 16.830000 ;
        RECT 22.515000 16.830000 23.155000 16.900000 ;
        RECT 22.585000 16.900000 23.225000 16.970000 ;
        RECT 22.655000 16.970000 23.295000 17.040000 ;
        RECT 22.725000 17.040000 23.365000 17.110000 ;
        RECT 22.795000 17.110000 23.435000 17.180000 ;
        RECT 22.865000 17.180000 23.505000 17.250000 ;
        RECT 22.935000 17.250000 23.575000 17.320000 ;
        RECT 23.005000 17.320000 23.645000 17.390000 ;
        RECT 23.075000 17.390000 23.715000 17.460000 ;
        RECT 23.145000 17.460000 23.785000 17.530000 ;
        RECT 23.215000 17.530000 23.855000 17.600000 ;
        RECT 23.285000 17.600000 23.925000 17.670000 ;
        RECT 23.355000 17.670000 23.995000 17.740000 ;
        RECT 23.425000 17.740000 24.065000 17.810000 ;
        RECT 23.495000 17.810000 24.135000 17.880000 ;
        RECT 23.565000 17.880000 24.205000 17.950000 ;
        RECT 23.635000 17.950000 24.275000 18.020000 ;
        RECT 23.705000 18.020000 24.345000 18.090000 ;
        RECT 23.775000 18.090000 24.415000 18.160000 ;
        RECT 23.845000 18.160000 24.485000 18.230000 ;
        RECT 23.915000 18.230000 24.555000 18.300000 ;
        RECT 23.985000 18.300000 24.625000 18.370000 ;
        RECT 24.015000 18.370000 24.695000 18.400000 ;
        RECT 24.085000 18.400000 24.725000 18.470000 ;
        RECT 24.155000 18.470000 24.725000 18.540000 ;
        RECT 24.225000 18.540000 24.725000 18.610000 ;
        RECT 24.225000 18.610000 24.725000 25.145000 ;
        RECT 24.225000 25.145000 24.725000 25.215000 ;
        RECT 24.225000 25.215000 24.795000 25.285000 ;
        RECT 24.225000 25.285000 24.865000 25.355000 ;
        RECT 24.295000 25.355000 24.935000 25.425000 ;
        RECT 24.325000 43.230000 24.640000 43.285000 ;
        RECT 24.365000 25.425000 25.005000 25.495000 ;
        RECT 24.395000 43.160000 24.695000 43.230000 ;
        RECT 24.435000 25.495000 25.075000 25.565000 ;
        RECT 24.465000 43.090000 24.765000 43.160000 ;
        RECT 24.505000 25.565000 25.145000 25.635000 ;
        RECT 24.535000 43.020000 24.835000 43.090000 ;
        RECT 24.575000 25.635000 25.215000 25.705000 ;
        RECT 24.605000 25.705000 25.285000 25.735000 ;
        RECT 24.605000 42.950000 24.905000 43.020000 ;
        RECT 24.675000 25.735000 25.315000 25.805000 ;
        RECT 24.675000 42.880000 24.975000 42.950000 ;
        RECT 24.745000 25.805000 25.315000 25.875000 ;
        RECT 24.745000 42.810000 25.045000 42.880000 ;
        RECT 24.815000 25.875000 25.315000 25.945000 ;
        RECT 24.815000 25.945000 25.315000 42.610000 ;
        RECT 24.815000 42.610000 25.250000 42.675000 ;
        RECT 24.815000 42.675000 25.185000 42.740000 ;
        RECT 24.815000 42.740000 25.115000 42.810000 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.555000 0.000000 15.135000 0.985000 ;
    END
  END PULLUP_H
  PIN TIE_HI_ESD
    ANTENNAPARTIALCUTAREA  0.045000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 28.185000 4.895000 30.220000 4.965000 ;
        RECT 28.185000 4.965000 30.150000 5.035000 ;
        RECT 28.185000 5.035000 30.080000 5.105000 ;
        RECT 28.185000 5.105000 30.010000 5.175000 ;
        RECT 28.185000 5.175000 29.940000 5.245000 ;
        RECT 28.185000 5.245000 29.870000 5.315000 ;
        RECT 28.185000 5.315000 29.800000 5.385000 ;
        RECT 28.185000 5.385000 29.730000 5.455000 ;
        RECT 28.185000 5.455000 29.660000 5.525000 ;
        RECT 28.185000 5.525000 29.640000 5.545000 ;
        RECT 29.395000 4.870000 30.290000 4.895000 ;
        RECT 29.465000 4.800000 30.315000 4.870000 ;
        RECT 29.535000 4.730000 30.385000 4.800000 ;
        RECT 29.605000 4.660000 30.455000 4.730000 ;
        RECT 29.675000 4.590000 30.525000 4.660000 ;
        RECT 29.745000 4.520000 30.595000 4.590000 ;
        RECT 29.815000 4.450000 30.665000 4.520000 ;
        RECT 29.885000 4.380000 30.735000 4.450000 ;
        RECT 29.955000 4.310000 30.805000 4.380000 ;
        RECT 30.025000 4.240000 30.875000 4.310000 ;
        RECT 30.095000 4.170000 30.945000 4.240000 ;
        RECT 30.165000 4.100000 31.015000 4.170000 ;
        RECT 30.235000 4.030000 31.085000 4.100000 ;
        RECT 30.295000 3.970000 31.155000 4.030000 ;
        RECT 30.365000 3.900000 31.155000 3.970000 ;
        RECT 30.435000 3.830000 31.155000 3.900000 ;
        RECT 30.505000 0.000000 31.155000 3.760000 ;
        RECT 30.505000 3.760000 31.155000 3.830000 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.505000 0.000000 31.155000 0.330000 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    ANTENNAPARTIALCUTAREA  0.045000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 27.580000 0.000000 28.230000 2.855000 ;
        RECT 27.580000 2.855000 28.230000 2.925000 ;
        RECT 27.580000 2.925000 28.300000 2.995000 ;
        RECT 27.580000 2.995000 28.370000 3.065000 ;
        RECT 27.580000 3.065000 28.440000 3.125000 ;
        RECT 27.650000 3.125000 28.500000 3.195000 ;
        RECT 27.720000 3.195000 28.570000 3.265000 ;
        RECT 27.790000 3.265000 28.640000 3.335000 ;
        RECT 27.860000 3.335000 28.710000 3.405000 ;
        RECT 27.915000 3.405000 28.780000 3.460000 ;
        RECT 27.985000 3.460000 28.835000 3.530000 ;
        RECT 28.055000 3.530000 28.835000 3.600000 ;
        RECT 28.125000 3.600000 28.835000 3.670000 ;
        RECT 28.185000 3.670000 28.835000 3.730000 ;
        RECT 28.185000 3.730000 28.835000 4.105000 ;
    END
    PORT
      LAYER met2 ;
        RECT 27.580000 0.000000 28.230000 0.330000 ;
    END
  END TIE_LO_ESD
  PIN TIE_WEAK_HI_H
    ANTENNAPARTIALCUTAREA  0.520000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.215000 0.000000 73.235000 0.770000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.860000 71.930000 66.310000 72.080000 ;
        RECT 64.860000 72.080000 66.160000 72.230000 ;
        RECT 64.860000 72.230000 66.010000 72.380000 ;
        RECT 64.860000 72.380000 65.990000 72.400000 ;
        RECT 64.860000 72.400000 65.990000 94.645000 ;
        RECT 64.990000 71.800000 66.460000 71.930000 ;
        RECT 65.140000 71.650000 66.590000 71.800000 ;
        RECT 65.290000 71.500000 66.740000 71.650000 ;
        RECT 65.440000 71.350000 66.890000 71.500000 ;
        RECT 65.590000 71.200000 67.040000 71.350000 ;
        RECT 65.740000 71.050000 67.190000 71.200000 ;
        RECT 65.890000 70.900000 67.340000 71.050000 ;
        RECT 66.040000 70.750000 67.490000 70.900000 ;
        RECT 66.190000 70.600000 67.640000 70.750000 ;
        RECT 66.340000 70.450000 67.790000 70.600000 ;
        RECT 66.490000 70.300000 67.940000 70.450000 ;
        RECT 66.640000 70.150000 68.090000 70.300000 ;
        RECT 66.790000 70.000000 68.240000 70.150000 ;
        RECT 66.940000 69.850000 68.390000 70.000000 ;
        RECT 67.090000 69.700000 68.540000 69.850000 ;
        RECT 67.240000 69.550000 68.690000 69.700000 ;
        RECT 67.390000 69.400000 68.840000 69.550000 ;
        RECT 67.540000 69.250000 68.990000 69.400000 ;
        RECT 67.690000 69.100000 69.140000 69.250000 ;
        RECT 67.840000 68.950000 69.290000 69.100000 ;
        RECT 67.990000 68.800000 69.440000 68.950000 ;
        RECT 68.140000 68.650000 69.590000 68.800000 ;
        RECT 68.290000 68.500000 69.740000 68.650000 ;
        RECT 68.440000 68.350000 69.890000 68.500000 ;
        RECT 68.590000 68.200000 70.040000 68.350000 ;
        RECT 68.740000 68.050000 70.190000 68.200000 ;
        RECT 68.890000 67.900000 70.340000 68.050000 ;
        RECT 69.040000 67.750000 70.490000 67.900000 ;
        RECT 69.190000 67.600000 70.640000 67.750000 ;
        RECT 69.340000 67.450000 70.790000 67.600000 ;
        RECT 69.490000 67.300000 70.940000 67.450000 ;
        RECT 69.640000 67.150000 71.090000 67.300000 ;
        RECT 69.790000 67.000000 71.240000 67.150000 ;
        RECT 69.940000 66.850000 71.390000 67.000000 ;
        RECT 70.090000 66.700000 71.540000 66.850000 ;
        RECT 70.240000 66.550000 71.690000 66.700000 ;
        RECT 70.390000 66.400000 71.840000 66.550000 ;
        RECT 70.540000 66.250000 71.990000 66.400000 ;
        RECT 70.690000 66.100000 72.140000 66.250000 ;
        RECT 70.840000 65.950000 72.290000 66.100000 ;
        RECT 70.990000 65.800000 72.440000 65.950000 ;
        RECT 71.140000 65.650000 72.590000 65.800000 ;
        RECT 71.290000 65.500000 72.740000 65.650000 ;
        RECT 71.440000 65.350000 72.890000 65.500000 ;
        RECT 71.590000 65.200000 73.040000 65.350000 ;
        RECT 71.740000 65.050000 73.190000 65.200000 ;
        RECT 71.890000 64.900000 73.340000 65.050000 ;
        RECT 72.040000 64.750000 73.490000 64.900000 ;
        RECT 72.190000  0.000000 73.260000 49.320000 ;
        RECT 72.190000 49.320000 73.260000 49.470000 ;
        RECT 72.190000 49.470000 73.410000 49.620000 ;
        RECT 72.190000 49.620000 73.560000 49.770000 ;
        RECT 72.190000 49.770000 73.710000 49.920000 ;
        RECT 72.190000 49.920000 73.860000 49.985000 ;
        RECT 72.190000 49.985000 73.925000 64.465000 ;
        RECT 72.190000 64.465000 73.860000 64.530000 ;
        RECT 72.190000 64.530000 73.795000 64.595000 ;
        RECT 72.190000 64.595000 73.790000 64.600000 ;
        RECT 72.190000 64.600000 73.640000 64.750000 ;
    END
  END TIE_WEAK_HI_H
  PIN XRES_H_N
    ANTENNAPARTIALCUTAREA  0.240000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.915000 0.000000 29.685000 0.335000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.170000 10.610000 29.050000 10.760000 ;
        RECT 28.170000 10.760000 28.900000 10.910000 ;
        RECT 28.170000 10.910000 28.900000 14.770000 ;
        RECT 28.185000 10.595000 29.200000 10.610000 ;
        RECT 28.335000 10.445000 29.215000 10.595000 ;
        RECT 28.485000 10.295000 29.365000 10.445000 ;
        RECT 28.635000 10.145000 29.515000 10.295000 ;
        RECT 28.785000  9.995000 29.665000 10.145000 ;
        RECT 28.935000  0.000000 29.665000  9.845000 ;
        RECT 28.935000  9.845000 29.665000  9.995000 ;
    END
  END XRES_H_N
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 41.655000 ;
        RECT 0.000000 41.655000 3.720000 46.170000 ;
        RECT 0.000000 46.170000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.655000 41.630000 75.000000 46.190000 ;
        RECT 73.730000 41.585000 75.000000 41.630000 ;
        RECT 73.730000 46.190000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT -0.265000 125.265000 75.000000 129.185000 ;
      RECT -0.265000 129.185000 41.620000 130.225000 ;
      RECT -0.160000 140.815000 75.160000 144.435000 ;
      RECT  0.000000  96.860000 58.340000  96.865000 ;
      RECT  0.000000  96.865000 75.000000  97.865000 ;
      RECT  0.000000  97.865000 58.340000  99.360000 ;
      RECT  0.000000  99.360000 75.000000 101.740000 ;
      RECT  0.000000 101.740000 58.340000 101.780000 ;
      RECT  0.000000 101.780000  0.165000 102.385000 ;
      RECT  0.000000 102.385000  0.455000 102.395000 ;
      RECT  0.000000 102.395000  0.595000 125.265000 ;
      RECT  0.000000 130.995000 38.355000 131.325000 ;
      RECT  0.000000 131.325000 13.200000 134.390000 ;
      RECT  0.000000 134.390000 75.000000 134.950000 ;
      RECT  0.000000 134.950000 52.445000 136.970000 ;
      RECT  0.000000 136.970000  1.045000 138.600000 ;
      RECT  0.000000 138.600000 75.000000 140.050000 ;
      RECT  0.700000 130.425000 42.015000 130.795000 ;
      RECT  0.700000 130.795000 38.355000 130.995000 ;
      RECT  0.985000   0.185000 33.890000   0.645000 ;
      RECT  0.985000   0.645000  4.525000   3.740000 ;
      RECT  0.985000   3.740000  7.065000   4.105000 ;
      RECT  0.985000 101.780000  2.645000 102.395000 ;
      RECT  1.015000   4.105000  7.065000   8.600000 ;
      RECT  1.015000   8.600000  5.625000  12.860000 ;
      RECT  1.015000  12.860000  6.055000  13.870000 ;
      RECT  1.015000  13.870000  5.625000  17.770000 ;
      RECT  1.015000  17.770000 14.130000  18.870000 ;
      RECT  1.015000  18.870000  5.605000  37.435000 ;
      RECT  1.015000  37.435000 14.270000  38.625000 ;
      RECT  1.015000  38.625000  4.525000  71.780000 ;
      RECT  1.015000  71.780000 31.450000  84.665000 ;
      RECT  1.100000  85.320000  2.790000  96.860000 ;
      RECT  1.145000  84.665000 31.450000  85.320000 ;
      RECT 11.005000  17.765000 11.270000  17.770000 ;
      RECT 11.270000  18.870000 14.130000  25.580000 ;
      RECT 13.095000   3.770000 16.800000   6.465000 ;
      RECT 13.095000   6.465000 32.410000   6.520000 ;
      RECT 13.095000   6.520000 32.395000   8.665000 ;
      RECT 13.460000  25.580000 14.130000  27.375000 ;
      RECT 13.460000  27.375000 20.685000  27.545000 ;
      RECT 13.460000  27.545000 14.130000  34.045000 ;
      RECT 14.130000 136.970000 52.445000 137.930000 ;
      RECT 14.130000 137.930000 75.000000 138.600000 ;
      RECT 14.165000  13.360000 14.435000  13.735000 ;
      RECT 14.185000   8.665000 14.385000  12.750000 ;
      RECT 14.480000  13.050000 24.760000  15.670000 ;
      RECT 16.115000  10.105000 16.285000  10.160000 ;
      RECT 16.115000  10.160000 16.800000  10.330000 ;
      RECT 16.115000  10.330000 16.285000  10.635000 ;
      RECT 16.130000  11.590000 16.800000  11.760000 ;
      RECT 16.630000  11.480000 16.800000  11.590000 ;
      RECT 16.630000  11.760000 16.800000  12.010000 ;
      RECT 16.950000  15.670000 24.760000  15.930000 ;
      RECT 16.950000  15.930000 32.350000  16.600000 ;
      RECT 16.950000  16.600000 26.460000  18.815000 ;
      RECT 17.885000   0.645000 33.890000   3.235000 ;
      RECT 18.700000  18.815000 26.460000  20.255000 ;
      RECT 18.885000  24.405000 20.685000  27.375000 ;
      RECT 19.155000  39.220000 26.270000  41.890000 ;
      RECT 19.155000  41.890000 32.495000  42.120000 ;
      RECT 19.155000  42.120000 32.435000  43.020000 ;
      RECT 20.685000  20.255000 26.460000  20.490000 ;
      RECT 20.855000  20.490000 26.460000  21.035000 ;
      RECT 20.855000  24.480000 26.460000  25.800000 ;
      RECT 21.135000  37.530000 26.270000  39.220000 ;
      RECT 23.730000  21.035000 26.460000  24.480000 ;
      RECT 24.035000 131.325000 25.835000 134.390000 ;
      RECT 24.435000  11.465000 25.140000  11.995000 ;
      RECT 24.470000   9.975000 25.105000  10.160000 ;
      RECT 24.470000  10.160000 25.140000  10.330000 ;
      RECT 24.470000  10.330000 25.105000  10.505000 ;
      RECT 25.070000  25.800000 26.460000  26.780000 ;
      RECT 25.070000  26.780000 32.625000  27.950000 ;
      RECT 25.070000  27.950000 27.385000  33.830000 ;
      RECT 25.070000  33.830000 32.435000  33.940000 ;
      RECT 25.070000  33.940000 32.495000  34.170000 ;
      RECT 25.070000  34.170000 26.270000  37.530000 ;
      RECT 25.140000  47.770000 31.450000  71.780000 ;
      RECT 26.480000  14.880000 26.650000  15.410000 ;
      RECT 26.975000  34.730000 31.525000  34.960000 ;
      RECT 26.975000  34.960000 27.205000  40.965000 ;
      RECT 26.975000  40.965000 31.525000  41.195000 ;
      RECT 27.370000  17.445000 27.540000  25.820000 ;
      RECT 27.760000  14.880000 27.930000  15.410000 ;
      RECT 27.850000  35.215000 30.690000  35.385000 ;
      RECT 28.665000  30.760000 28.835000  31.290000 ;
      RECT 28.665000  31.845000 28.835000  32.375000 ;
      RECT 29.035000  28.960000 29.205000  29.490000 ;
      RECT 29.035000  30.070000 29.205000  30.600000 ;
      RECT 29.065000  31.460000 29.595000  31.630000 ;
      RECT 29.150000  18.365000 29.680000  18.535000 ;
      RECT 29.150000  20.125000 29.680000  20.295000 ;
      RECT 29.330000  24.890000 30.490000  25.220000 ;
      RECT 29.455000   3.235000 32.410000   6.465000 ;
      RECT 30.105000  25.405000 30.635000  25.575000 ;
      RECT 30.115000  29.700000 30.645000  29.870000 ;
      RECT 30.215000  14.720000 30.385000  15.250000 ;
      RECT 30.415000  19.390000 30.585000  19.920000 ;
      RECT 30.415000  20.510000 30.585000  21.040000 ;
      RECT 30.835000  17.635000 31.005000  18.165000 ;
      RECT 30.835000  18.755000 31.005000  19.285000 ;
      RECT 30.960000  46.750000 31.490000  46.920000 ;
      RECT 31.130000  46.485000 31.490000  46.750000 ;
      RECT 31.130000  46.920000 31.490000  47.155000 ;
      RECT 31.295000  34.960000 31.525000  40.965000 ;
      RECT 31.495000  14.720000 31.665000  15.250000 ;
      RECT 32.155000  28.780000 32.325000  32.550000 ;
      RECT 32.265000  34.170000 32.495000  41.890000 ;
      RECT 33.420000  73.960000 33.870000  81.465000 ;
      RECT 33.445000  82.260000 34.600000  83.340000 ;
      RECT 33.535000  81.905000 34.065000  82.075000 ;
      RECT 34.850000  83.100000 35.380000  83.270000 ;
      RECT 35.090000   0.900000 38.860000   1.070000 ;
      RECT 35.160000   1.070000 38.860000   1.080000 ;
      RECT 36.555000 131.325000 38.355000 134.390000 ;
      RECT 38.970000 133.145000 40.600000 133.825000 ;
      RECT 40.040000   0.195000 74.560000   5.755000 ;
      RECT 40.335000   5.755000 74.560000   5.960000 ;
      RECT 40.495000 130.795000 42.015000 130.995000 ;
      RECT 40.495000 130.995000 75.000000 132.595000 ;
      RECT 42.840000 129.770000 43.730000 130.440000 ;
      RECT 43.350000  60.495000 43.720000  78.760000 ;
      RECT 48.290000 129.770000 50.440000 130.440000 ;
      RECT 51.880000 133.145000 52.770000 133.815000 ;
      RECT 53.575000 135.430000 55.095000 137.450000 ;
      RECT 53.970000   5.960000 74.560000   6.580000 ;
      RECT 55.000000 129.770000 56.460000 130.440000 ;
      RECT 58.340000 102.310000 72.060000 102.395000 ;
      RECT 60.770000 133.145000 61.800000 133.815000 ;
      RECT 60.855000 129.760000 61.780000 130.430000 ;
      RECT 62.040000 129.185000 75.000000 130.225000 ;
      RECT 62.065000 132.595000 75.000000 134.390000 ;
      RECT 62.730000   6.580000 63.170000  59.670000 ;
      RECT 63.130000  60.940000 63.180000  85.005000 ;
      RECT 67.105000 134.950000 75.000000 137.930000 ;
      RECT 68.960000  85.895000 71.490000  86.125000 ;
      RECT 68.960000  86.125000 74.315000  94.410000 ;
      RECT 69.260000  94.410000 74.315000  96.865000 ;
      RECT 72.060000  97.865000 75.000000  99.360000 ;
      RECT 72.060000 101.740000 75.000000 101.780000 ;
      RECT 73.265000   6.580000 74.560000  84.995000 ;
      RECT 73.265000  84.995000 73.855000  85.020000 ;
      RECT 74.355000 101.780000 75.000000 125.265000 ;
    LAYER met1 ;
      RECT -0.145000  95.895000  2.680000  95.965000 ;
      RECT -0.145000  95.965000  2.750000  96.035000 ;
      RECT -0.145000  96.035000  2.820000  96.105000 ;
      RECT -0.145000  96.105000  2.890000  96.175000 ;
      RECT -0.145000  96.175000  2.960000  96.245000 ;
      RECT -0.145000  96.245000  3.030000  96.315000 ;
      RECT -0.145000  96.315000  3.100000  96.385000 ;
      RECT -0.145000  96.385000  3.170000  96.455000 ;
      RECT -0.145000  96.455000  3.240000  96.525000 ;
      RECT -0.145000  96.525000  3.310000  96.595000 ;
      RECT -0.145000  96.545000  3.325000  96.610000 ;
      RECT -0.145000  96.545000  3.325000  96.610000 ;
      RECT -0.145000  96.595000  3.380000  96.665000 ;
      RECT -0.145000  96.610000  3.395000  96.680000 ;
      RECT -0.145000  96.610000  3.395000  96.680000 ;
      RECT -0.145000  96.665000  3.450000  96.735000 ;
      RECT -0.145000  96.680000  3.465000  96.750000 ;
      RECT -0.145000  96.680000  3.465000  96.750000 ;
      RECT -0.145000  96.735000  3.520000  96.805000 ;
      RECT -0.145000  96.750000  3.535000  96.820000 ;
      RECT -0.145000  96.750000  3.535000  96.820000 ;
      RECT -0.145000  96.805000  3.590000  96.875000 ;
      RECT -0.145000  96.820000  3.605000  96.890000 ;
      RECT -0.145000  96.820000  3.605000  96.890000 ;
      RECT -0.145000  96.875000  3.660000  96.945000 ;
      RECT -0.145000  96.890000  3.675000  96.960000 ;
      RECT -0.145000  96.890000  3.675000  96.960000 ;
      RECT -0.145000  96.945000  3.730000  97.015000 ;
      RECT -0.145000  96.960000  3.745000  97.030000 ;
      RECT -0.145000  96.960000  3.745000  97.030000 ;
      RECT -0.145000  97.015000  3.800000  97.085000 ;
      RECT -0.145000  97.030000  3.815000  97.100000 ;
      RECT -0.145000  97.030000  3.815000  97.100000 ;
      RECT -0.145000  97.085000  3.870000  97.155000 ;
      RECT -0.145000  97.100000  3.885000  97.170000 ;
      RECT -0.145000  97.100000  3.885000  97.170000 ;
      RECT -0.145000  97.155000  3.940000  97.225000 ;
      RECT -0.145000  97.170000  3.955000  97.240000 ;
      RECT -0.145000  97.170000  3.955000  97.240000 ;
      RECT -0.145000  97.225000  4.010000  97.295000 ;
      RECT -0.145000  97.240000  4.025000  97.310000 ;
      RECT -0.145000  97.240000  4.025000  97.310000 ;
      RECT -0.145000  97.295000  4.080000  97.365000 ;
      RECT -0.145000  97.310000  4.095000  97.380000 ;
      RECT -0.145000  97.310000  4.095000  97.380000 ;
      RECT -0.145000  97.365000  4.150000  97.435000 ;
      RECT -0.145000  97.380000  4.165000  97.450000 ;
      RECT -0.145000  97.380000  4.165000  97.450000 ;
      RECT -0.145000  97.435000  4.220000  97.505000 ;
      RECT -0.145000  97.450000  4.235000  97.520000 ;
      RECT -0.145000  97.450000  4.235000  97.520000 ;
      RECT -0.145000  97.505000  4.290000  97.530000 ;
      RECT -0.145000  97.520000  4.305000  97.530000 ;
      RECT -0.145000  97.520000  4.305000  97.530000 ;
      RECT -0.145000  97.530000 56.545000 100.330000 ;
      RECT -0.145000 100.330000 56.545000 101.420000 ;
      RECT -0.145000 125.440000 14.680000 125.510000 ;
      RECT -0.145000 125.440000 14.680000 125.510000 ;
      RECT -0.145000 125.510000 14.610000 125.580000 ;
      RECT -0.145000 125.510000 14.610000 125.580000 ;
      RECT -0.145000 125.580000 14.540000 125.650000 ;
      RECT -0.145000 125.580000 14.540000 125.650000 ;
      RECT -0.145000 125.650000 14.470000 125.720000 ;
      RECT -0.145000 125.650000 14.470000 125.720000 ;
      RECT -0.145000 125.720000 14.400000 125.790000 ;
      RECT -0.145000 125.720000 14.400000 125.790000 ;
      RECT -0.145000 125.790000 14.330000 125.860000 ;
      RECT -0.145000 125.790000 14.330000 125.860000 ;
      RECT -0.145000 125.860000 14.260000 125.930000 ;
      RECT -0.145000 125.860000 14.260000 125.930000 ;
      RECT -0.145000 125.930000 14.190000 126.000000 ;
      RECT -0.145000 125.930000 14.190000 126.000000 ;
      RECT -0.145000 126.000000 14.120000 126.070000 ;
      RECT -0.145000 126.000000 14.120000 126.070000 ;
      RECT -0.145000 126.070000 14.050000 126.140000 ;
      RECT -0.145000 126.070000 14.050000 126.140000 ;
      RECT -0.145000 126.140000 13.980000 126.210000 ;
      RECT -0.145000 126.140000 13.980000 126.210000 ;
      RECT -0.145000 126.210000 13.910000 126.280000 ;
      RECT -0.145000 126.210000 13.910000 126.280000 ;
      RECT -0.145000 126.280000 13.840000 126.350000 ;
      RECT -0.145000 126.280000 13.840000 126.350000 ;
      RECT -0.145000 126.350000 13.770000 126.420000 ;
      RECT -0.145000 126.350000 13.770000 126.420000 ;
      RECT -0.145000 126.420000 13.700000 126.490000 ;
      RECT -0.145000 126.420000 13.700000 126.490000 ;
      RECT -0.145000 126.490000 13.630000 126.560000 ;
      RECT -0.145000 126.490000 13.630000 126.560000 ;
      RECT -0.145000 126.560000 13.560000 126.630000 ;
      RECT -0.145000 126.560000 13.560000 126.630000 ;
      RECT -0.145000 126.630000 13.490000 126.700000 ;
      RECT -0.145000 126.630000 13.490000 126.700000 ;
      RECT -0.145000 126.700000 13.420000 126.770000 ;
      RECT -0.145000 126.700000 13.420000 126.770000 ;
      RECT -0.145000 126.770000 13.350000 126.840000 ;
      RECT -0.145000 126.770000 13.350000 126.840000 ;
      RECT -0.145000 126.840000 13.280000 126.910000 ;
      RECT -0.145000 126.840000 13.280000 126.910000 ;
      RECT -0.145000 126.910000 13.210000 126.980000 ;
      RECT -0.145000 126.910000 13.210000 126.980000 ;
      RECT -0.145000 126.980000 13.140000 127.050000 ;
      RECT -0.145000 126.980000 13.140000 127.050000 ;
      RECT -0.145000 127.050000 13.070000 127.120000 ;
      RECT -0.145000 127.050000 13.070000 127.120000 ;
      RECT -0.145000 127.120000 13.000000 127.190000 ;
      RECT -0.145000 127.120000 13.000000 127.190000 ;
      RECT -0.145000 127.190000 12.930000 127.260000 ;
      RECT -0.145000 127.190000 12.930000 127.260000 ;
      RECT -0.145000 127.260000 12.860000 127.330000 ;
      RECT -0.145000 127.260000 12.860000 127.330000 ;
      RECT -0.145000 127.330000 12.790000 127.400000 ;
      RECT -0.145000 127.330000 12.790000 127.400000 ;
      RECT -0.145000 127.400000 12.720000 127.470000 ;
      RECT -0.145000 127.400000 12.720000 127.470000 ;
      RECT -0.145000 127.470000 12.650000 127.540000 ;
      RECT -0.145000 127.470000 12.650000 127.540000 ;
      RECT -0.145000 127.540000 12.580000 127.610000 ;
      RECT -0.145000 127.540000 12.580000 127.610000 ;
      RECT -0.145000 127.610000 12.510000 127.680000 ;
      RECT -0.145000 127.610000 12.510000 127.680000 ;
      RECT -0.145000 127.680000 12.440000 127.750000 ;
      RECT -0.145000 127.680000 12.440000 127.750000 ;
      RECT -0.145000 127.750000 12.370000 127.820000 ;
      RECT -0.145000 127.750000 12.370000 127.820000 ;
      RECT -0.145000 127.820000 12.300000 127.890000 ;
      RECT -0.145000 127.820000 12.300000 127.890000 ;
      RECT -0.145000 127.890000 12.230000 127.960000 ;
      RECT -0.145000 127.890000 12.230000 127.960000 ;
      RECT -0.145000 127.960000 12.160000 128.030000 ;
      RECT -0.145000 127.960000 12.160000 128.030000 ;
      RECT -0.145000 128.030000 12.090000 128.100000 ;
      RECT -0.145000 128.030000 12.090000 128.100000 ;
      RECT -0.145000 128.100000 12.020000 128.170000 ;
      RECT -0.145000 128.100000 12.020000 128.170000 ;
      RECT -0.145000 128.170000 11.950000 128.240000 ;
      RECT -0.145000 128.170000 11.950000 128.240000 ;
      RECT -0.145000 128.240000 11.930000 128.260000 ;
      RECT -0.145000 128.240000 11.930000 128.260000 ;
      RECT -0.145000 128.260000 11.860000 128.330000 ;
      RECT -0.145000 128.260000 11.860000 128.330000 ;
      RECT -0.145000 128.330000 11.790000 128.400000 ;
      RECT -0.145000 128.330000 11.790000 128.400000 ;
      RECT -0.145000 128.400000 11.720000 128.470000 ;
      RECT -0.145000 128.400000 11.720000 128.470000 ;
      RECT -0.145000 128.470000 11.650000 128.540000 ;
      RECT -0.145000 128.470000 11.650000 128.540000 ;
      RECT -0.145000 128.540000 11.580000 128.610000 ;
      RECT -0.145000 128.540000 11.580000 128.610000 ;
      RECT -0.145000 128.610000 11.510000 128.680000 ;
      RECT -0.145000 128.610000 11.510000 128.680000 ;
      RECT -0.145000 128.680000 11.440000 128.750000 ;
      RECT -0.145000 128.680000 11.440000 128.750000 ;
      RECT -0.145000 128.750000 11.370000 128.820000 ;
      RECT -0.145000 128.750000 11.370000 128.820000 ;
      RECT -0.145000 128.820000 11.300000 128.890000 ;
      RECT -0.145000 128.820000 11.300000 128.890000 ;
      RECT -0.145000 128.890000 11.230000 128.960000 ;
      RECT -0.145000 128.890000 11.230000 128.960000 ;
      RECT -0.145000 128.960000 11.160000 129.030000 ;
      RECT -0.145000 128.960000 11.160000 129.030000 ;
      RECT -0.145000 129.030000 11.090000 129.100000 ;
      RECT -0.145000 129.030000 11.090000 129.100000 ;
      RECT -0.145000 129.100000 11.020000 129.170000 ;
      RECT -0.145000 129.100000 11.020000 129.170000 ;
      RECT -0.145000 129.170000 10.950000 129.240000 ;
      RECT -0.145000 129.170000 10.950000 129.240000 ;
      RECT -0.145000 129.240000 10.880000 129.310000 ;
      RECT -0.145000 129.240000 10.880000 129.310000 ;
      RECT -0.145000 129.310000 10.810000 129.380000 ;
      RECT -0.145000 129.310000 10.810000 129.380000 ;
      RECT -0.145000 129.380000 10.740000 129.450000 ;
      RECT -0.145000 129.380000 10.740000 129.450000 ;
      RECT -0.145000 129.450000 10.670000 129.520000 ;
      RECT -0.145000 129.450000 10.670000 129.520000 ;
      RECT -0.145000 129.520000 10.600000 129.590000 ;
      RECT -0.145000 129.520000 10.600000 129.590000 ;
      RECT -0.145000 129.590000 10.530000 129.660000 ;
      RECT -0.145000 129.590000 10.530000 129.660000 ;
      RECT -0.145000 129.660000 10.460000 129.730000 ;
      RECT -0.145000 129.660000 10.460000 129.730000 ;
      RECT -0.145000 129.730000 10.390000 129.800000 ;
      RECT -0.145000 129.730000 10.390000 129.800000 ;
      RECT -0.145000 129.800000 10.320000 129.870000 ;
      RECT -0.145000 129.800000 10.320000 129.870000 ;
      RECT -0.145000 129.870000 10.250000 129.940000 ;
      RECT -0.145000 129.870000 10.250000 129.940000 ;
      RECT -0.145000 129.940000 10.180000 130.010000 ;
      RECT -0.145000 129.940000 10.180000 130.010000 ;
      RECT -0.145000 130.010000 10.110000 130.080000 ;
      RECT -0.145000 130.010000 10.110000 130.080000 ;
      RECT -0.145000 130.080000 10.040000 130.150000 ;
      RECT -0.145000 130.080000 10.040000 130.150000 ;
      RECT -0.145000 130.150000  9.970000 130.220000 ;
      RECT -0.145000 130.150000  9.970000 130.220000 ;
      RECT -0.145000 131.275000  0.940000 131.345000 ;
      RECT -0.145000 131.275000  0.940000 131.345000 ;
      RECT -0.145000 131.345000  1.010000 131.415000 ;
      RECT -0.145000 131.345000  1.010000 131.415000 ;
      RECT -0.145000 131.415000  1.080000 131.485000 ;
      RECT -0.145000 131.415000  1.080000 131.485000 ;
      RECT -0.145000 131.485000  1.150000 131.555000 ;
      RECT -0.145000 131.485000  1.150000 131.555000 ;
      RECT -0.145000 131.555000  1.220000 131.625000 ;
      RECT -0.145000 131.555000  1.220000 131.625000 ;
      RECT -0.145000 131.625000  1.290000 131.695000 ;
      RECT -0.145000 131.625000  1.290000 131.695000 ;
      RECT -0.145000 131.695000  1.360000 131.765000 ;
      RECT -0.145000 131.695000  1.360000 131.765000 ;
      RECT -0.145000 131.765000  1.430000 131.835000 ;
      RECT -0.145000 131.765000  1.430000 131.835000 ;
      RECT -0.145000 131.835000  1.500000 131.905000 ;
      RECT -0.145000 131.835000  1.500000 131.905000 ;
      RECT -0.145000 131.905000  1.570000 131.975000 ;
      RECT -0.145000 131.905000  1.570000 131.975000 ;
      RECT -0.145000 131.975000  1.640000 132.045000 ;
      RECT -0.145000 131.975000  1.640000 132.045000 ;
      RECT -0.145000 132.045000  1.710000 132.115000 ;
      RECT -0.145000 132.045000  1.710000 132.115000 ;
      RECT -0.145000 132.115000  1.780000 132.185000 ;
      RECT -0.145000 132.115000  1.780000 132.185000 ;
      RECT -0.145000 132.185000  1.850000 132.255000 ;
      RECT -0.145000 132.185000  1.850000 132.255000 ;
      RECT -0.145000 132.255000  1.920000 132.325000 ;
      RECT -0.145000 132.255000  1.920000 132.325000 ;
      RECT -0.145000 132.325000  1.990000 132.395000 ;
      RECT -0.145000 132.325000  1.990000 132.395000 ;
      RECT -0.145000 132.395000  2.060000 132.465000 ;
      RECT -0.145000 132.395000  2.060000 132.465000 ;
      RECT -0.145000 132.465000  2.130000 132.535000 ;
      RECT -0.145000 132.465000  2.130000 132.535000 ;
      RECT -0.145000 132.535000  2.200000 132.605000 ;
      RECT -0.145000 132.535000  2.200000 132.605000 ;
      RECT -0.145000 132.605000  2.270000 132.675000 ;
      RECT -0.145000 132.605000  2.270000 132.675000 ;
      RECT -0.145000 132.675000  2.340000 132.740000 ;
      RECT -0.145000 132.675000  2.340000 132.740000 ;
      RECT -0.145000 132.740000  2.405000 132.810000 ;
      RECT -0.145000 132.740000  2.405000 132.810000 ;
      RECT -0.145000 132.810000  2.475000 132.880000 ;
      RECT -0.145000 132.810000  2.475000 132.880000 ;
      RECT -0.145000 132.880000  2.545000 132.950000 ;
      RECT -0.145000 132.880000  2.545000 132.950000 ;
      RECT -0.145000 132.950000  2.615000 133.020000 ;
      RECT -0.145000 132.950000  2.615000 133.020000 ;
      RECT -0.145000 133.020000  2.685000 133.090000 ;
      RECT -0.145000 133.020000  2.685000 133.090000 ;
      RECT -0.145000 133.090000  2.755000 133.160000 ;
      RECT -0.145000 133.090000  2.755000 133.160000 ;
      RECT -0.145000 133.160000  2.825000 133.230000 ;
      RECT -0.145000 133.160000  2.825000 133.230000 ;
      RECT -0.145000 133.230000  2.895000 133.300000 ;
      RECT -0.145000 133.230000  2.895000 133.300000 ;
      RECT -0.145000 133.300000  2.965000 133.370000 ;
      RECT -0.145000 133.300000  2.965000 133.370000 ;
      RECT -0.145000 133.370000  3.035000 133.440000 ;
      RECT -0.145000 133.370000  3.035000 133.440000 ;
      RECT -0.145000 133.440000  3.105000 133.510000 ;
      RECT -0.145000 133.440000  3.105000 133.510000 ;
      RECT -0.145000 133.510000  3.175000 133.580000 ;
      RECT -0.145000 133.510000  3.175000 133.580000 ;
      RECT -0.145000 133.580000  3.245000 133.650000 ;
      RECT -0.145000 133.580000  3.245000 133.650000 ;
      RECT -0.145000 133.650000  3.315000 133.720000 ;
      RECT -0.145000 133.650000  3.315000 133.720000 ;
      RECT -0.145000 133.720000  3.385000 133.790000 ;
      RECT -0.145000 133.720000  3.385000 133.790000 ;
      RECT -0.145000 133.790000  3.455000 133.860000 ;
      RECT -0.145000 133.790000  3.455000 133.860000 ;
      RECT -0.145000 133.860000  3.525000 133.930000 ;
      RECT -0.145000 133.860000  3.525000 133.930000 ;
      RECT -0.145000 133.930000  3.595000 134.000000 ;
      RECT -0.145000 133.930000  3.595000 134.000000 ;
      RECT -0.145000 134.000000  3.665000 134.070000 ;
      RECT -0.145000 134.000000  3.665000 134.070000 ;
      RECT -0.145000 134.070000  3.735000 134.140000 ;
      RECT -0.145000 134.070000  3.735000 134.140000 ;
      RECT -0.145000 134.140000  3.805000 134.180000 ;
      RECT -0.145000 134.140000  3.805000 134.180000 ;
      RECT -0.145000 134.180000  3.775000 134.250000 ;
      RECT -0.145000 134.180000  3.775000 134.250000 ;
      RECT -0.145000 134.250000  3.700000 134.320000 ;
      RECT -0.145000 134.250000  3.700000 134.320000 ;
      RECT -0.145000 134.320000  3.635000 134.390000 ;
      RECT -0.145000 134.320000  3.635000 134.390000 ;
      RECT -0.145000 134.390000  3.560000 134.460000 ;
      RECT -0.145000 134.390000  3.560000 134.460000 ;
      RECT -0.145000 134.460000  3.490000 134.530000 ;
      RECT -0.145000 134.460000  3.490000 134.530000 ;
      RECT -0.145000 134.530000  3.420000 134.600000 ;
      RECT -0.145000 134.530000  3.420000 134.600000 ;
      RECT -0.145000 134.600000  3.350000 134.670000 ;
      RECT -0.145000 134.600000  3.350000 134.670000 ;
      RECT -0.145000 134.670000  3.280000 134.740000 ;
      RECT -0.145000 134.670000  3.280000 134.740000 ;
      RECT -0.145000 134.740000  3.210000 134.810000 ;
      RECT -0.145000 134.740000  3.210000 134.810000 ;
      RECT -0.145000 134.810000  3.140000 134.880000 ;
      RECT -0.145000 134.810000  3.140000 134.880000 ;
      RECT -0.145000 134.880000  3.070000 134.950000 ;
      RECT -0.145000 134.880000  3.070000 134.950000 ;
      RECT -0.145000 134.950000  3.000000 135.020000 ;
      RECT -0.145000 134.950000  3.000000 135.020000 ;
      RECT -0.145000 135.020000  2.930000 135.090000 ;
      RECT -0.145000 135.020000  2.930000 135.090000 ;
      RECT -0.145000 135.090000  2.860000 135.160000 ;
      RECT -0.145000 135.090000  2.860000 135.160000 ;
      RECT -0.145000 135.160000  2.790000 135.230000 ;
      RECT -0.145000 135.160000  2.790000 135.230000 ;
      RECT -0.145000 135.230000  2.720000 135.300000 ;
      RECT -0.145000 135.230000  2.720000 135.300000 ;
      RECT -0.145000 135.300000  2.650000 135.370000 ;
      RECT -0.145000 135.300000  2.650000 135.370000 ;
      RECT -0.145000 135.370000  2.580000 135.440000 ;
      RECT -0.145000 135.370000  2.580000 135.440000 ;
      RECT -0.145000 135.440000  2.550000 135.470000 ;
      RECT -0.145000 135.440000  2.550000 135.470000 ;
      RECT -0.145000 135.470000  2.480000 135.540000 ;
      RECT -0.145000 135.470000  2.480000 135.540000 ;
      RECT -0.145000 135.540000  2.410000 135.610000 ;
      RECT -0.145000 135.540000  2.410000 135.610000 ;
      RECT -0.145000 135.610000  2.340000 135.680000 ;
      RECT -0.145000 135.610000  2.340000 135.680000 ;
      RECT -0.145000 135.680000  2.270000 135.750000 ;
      RECT -0.145000 135.680000  2.270000 135.750000 ;
      RECT -0.145000 135.750000  2.200000 135.820000 ;
      RECT -0.145000 135.750000  2.200000 135.820000 ;
      RECT -0.145000 135.820000  2.130000 135.890000 ;
      RECT -0.145000 135.820000  2.130000 135.890000 ;
      RECT -0.145000 135.890000  2.060000 135.960000 ;
      RECT -0.145000 135.890000  2.060000 135.960000 ;
      RECT -0.145000 135.960000  1.990000 136.030000 ;
      RECT -0.145000 135.960000  1.990000 136.030000 ;
      RECT -0.145000 136.030000  1.920000 136.100000 ;
      RECT -0.145000 136.030000  1.920000 136.100000 ;
      RECT -0.145000 136.100000  1.850000 136.170000 ;
      RECT -0.145000 136.100000  1.850000 136.170000 ;
      RECT -0.145000 136.170000  1.780000 136.240000 ;
      RECT -0.145000 136.170000  1.780000 136.240000 ;
      RECT -0.145000 136.240000  1.710000 136.310000 ;
      RECT -0.145000 136.240000  1.710000 136.310000 ;
      RECT -0.145000 136.310000  1.640000 136.380000 ;
      RECT -0.145000 136.310000  1.640000 136.380000 ;
      RECT -0.145000 136.380000  1.570000 136.450000 ;
      RECT -0.145000 136.380000  1.570000 136.450000 ;
      RECT -0.145000 136.450000  1.495000 136.520000 ;
      RECT -0.145000 136.450000  1.495000 136.520000 ;
      RECT -0.145000 136.520000  1.425000 136.590000 ;
      RECT -0.145000 136.520000  1.425000 136.590000 ;
      RECT -0.145000 136.590000  1.355000 136.660000 ;
      RECT -0.145000 136.590000  1.355000 136.660000 ;
      RECT -0.145000 136.660000  1.285000 136.730000 ;
      RECT -0.145000 136.660000  1.285000 136.730000 ;
      RECT -0.145000 136.730000  1.215000 136.800000 ;
      RECT -0.145000 136.730000  1.215000 136.800000 ;
      RECT -0.145000 136.800000  1.145000 136.870000 ;
      RECT -0.145000 136.800000  1.145000 136.870000 ;
      RECT -0.145000 136.870000  1.075000 136.940000 ;
      RECT -0.145000 136.870000  1.075000 136.940000 ;
      RECT -0.145000 136.940000  1.005000 137.010000 ;
      RECT -0.145000 136.940000  1.005000 137.010000 ;
      RECT -0.145000 137.010000  0.935000 137.080000 ;
      RECT -0.145000 137.010000  0.935000 137.080000 ;
      RECT -0.145000 137.080000  0.865000 137.150000 ;
      RECT -0.145000 137.080000  0.865000 137.150000 ;
      RECT -0.145000 137.150000  0.795000 137.220000 ;
      RECT -0.145000 137.150000  0.795000 137.220000 ;
      RECT -0.145000 137.220000  0.725000 137.290000 ;
      RECT -0.145000 137.220000  0.725000 137.290000 ;
      RECT -0.145000 137.290000  0.655000 137.360000 ;
      RECT -0.145000 137.290000  0.655000 137.360000 ;
      RECT -0.145000 137.360000  0.585000 137.430000 ;
      RECT -0.145000 137.360000  0.585000 137.430000 ;
      RECT -0.145000 137.430000  0.515000 137.500000 ;
      RECT -0.145000 137.430000  0.515000 137.500000 ;
      RECT -0.145000 137.500000  0.445000 137.570000 ;
      RECT -0.145000 137.500000  0.445000 137.570000 ;
      RECT -0.145000 137.570000  0.375000 137.640000 ;
      RECT -0.145000 137.570000  0.375000 137.640000 ;
      RECT -0.145000 137.640000  0.305000 137.710000 ;
      RECT -0.145000 137.640000  0.305000 137.710000 ;
      RECT -0.145000 137.710000  0.235000 137.780000 ;
      RECT -0.145000 137.710000  0.235000 137.780000 ;
      RECT -0.145000 137.780000  0.165000 137.850000 ;
      RECT -0.145000 137.780000  0.165000 137.850000 ;
      RECT -0.145000 137.850000  0.095000 137.920000 ;
      RECT -0.145000 137.850000  0.095000 137.920000 ;
      RECT -0.145000 137.920000  0.025000 137.990000 ;
      RECT -0.145000 137.920000  0.025000 137.990000 ;
      RECT -0.145000 137.990000 -0.045000 138.060000 ;
      RECT -0.145000 137.990000 -0.045000 138.060000 ;
      RECT -0.145000 138.060000 -0.115000 138.130000 ;
      RECT -0.145000 138.060000 -0.115000 138.130000 ;
      RECT -0.145000 138.160000  0.940000 139.015000 ;
      RECT -0.145000 139.015000  0.940000 139.085000 ;
      RECT -0.145000 139.085000  1.010000 139.155000 ;
      RECT -0.145000 139.155000  1.080000 139.225000 ;
      RECT -0.145000 139.225000  1.150000 139.295000 ;
      RECT -0.145000 139.295000  1.220000 139.365000 ;
      RECT -0.145000 139.365000  1.290000 139.435000 ;
      RECT -0.145000 139.435000  1.360000 139.505000 ;
      RECT -0.145000 139.505000 11.105000 139.540000 ;
      RECT -0.145000 139.540000 11.140000 139.575000 ;
      RECT -0.145000 139.575000 69.715000 139.645000 ;
      RECT -0.145000 139.645000 69.785000 139.715000 ;
      RECT -0.145000 139.715000 69.855000 139.785000 ;
      RECT -0.145000 139.785000 69.925000 139.850000 ;
      RECT -0.145000 139.850000  1.385000 139.920000 ;
      RECT -0.145000 139.920000  1.315000 139.990000 ;
      RECT -0.145000 139.990000  1.245000 140.060000 ;
      RECT -0.145000 140.060000  1.175000 140.130000 ;
      RECT -0.145000 140.130000  1.105000 140.200000 ;
      RECT -0.145000 140.200000  1.035000 140.270000 ;
      RECT -0.145000 140.270000  0.965000 140.340000 ;
      RECT -0.145000 140.340000  0.940000 140.365000 ;
      RECT -0.145000 140.365000  0.940000 143.640000 ;
      RECT -0.145000 143.640000  0.940000 143.710000 ;
      RECT -0.145000 143.710000  1.010000 143.780000 ;
      RECT -0.145000 143.780000  1.080000 143.850000 ;
      RECT -0.145000 143.850000  1.150000 143.920000 ;
      RECT -0.145000 143.920000  1.220000 143.990000 ;
      RECT -0.145000 143.990000  1.290000 144.060000 ;
      RECT -0.145000 144.060000  1.360000 144.130000 ;
      RECT -0.145000 144.130000  1.430000 144.200000 ;
      RECT -0.145000 144.200000  1.500000 144.270000 ;
      RECT -0.145000 144.270000  1.570000 144.340000 ;
      RECT -0.145000 144.340000  1.640000 144.410000 ;
      RECT -0.145000 144.410000  1.710000 144.480000 ;
      RECT -0.145000 144.480000  1.780000 144.550000 ;
      RECT -0.145000 144.550000  1.850000 144.620000 ;
      RECT -0.145000 144.620000  1.920000 144.690000 ;
      RECT -0.145000 144.690000  1.990000 144.760000 ;
      RECT -0.145000 144.760000  2.060000 144.830000 ;
      RECT -0.145000 144.830000  2.130000 144.900000 ;
      RECT -0.145000 144.900000  2.200000 144.970000 ;
      RECT -0.145000 144.970000  2.270000 145.040000 ;
      RECT -0.145000 145.040000  2.340000 145.110000 ;
      RECT -0.145000 145.110000  2.410000 145.130000 ;
      RECT -0.125000  96.525000  3.310000  96.545000 ;
      RECT -0.125000  96.525000  3.310000  96.545000 ;
      RECT -0.115000 138.130000  0.940000 138.160000 ;
      RECT -0.055000  96.455000  3.240000  96.525000 ;
      RECT -0.055000  96.455000  3.240000  96.525000 ;
      RECT -0.045000 138.060000  0.940000 138.130000 ;
      RECT  0.000000   0.000000  0.705000  84.590000 ;
      RECT  0.000000   0.000000 12.145000   6.435000 ;
      RECT  0.000000   6.435000 11.775000   6.805000 ;
      RECT  0.000000   6.805000 12.230000   6.980000 ;
      RECT  0.000000   6.980000 12.555000   7.310000 ;
      RECT  0.000000   7.310000 12.555000  10.370000 ;
      RECT  0.000000  10.370000 12.660000  10.445000 ;
      RECT  0.000000  10.445000 14.415000  12.400000 ;
      RECT  0.000000  12.400000 18.075000  16.060000 ;
      RECT  0.000000  16.060000 24.085000  18.665000 ;
      RECT  0.000000  18.665000 24.085000  25.415000 ;
      RECT  0.000000  25.415000 24.675000  26.005000 ;
      RECT  0.000000  26.005000 24.675000  42.680000 ;
      RECT  0.000000  42.680000 24.210000  43.145000 ;
      RECT  0.000000  43.145000  5.925000  43.685000 ;
      RECT  0.000000  43.685000 75.000000 200.000000 ;
      RECT  0.000000  84.590000  0.705000  84.660000 ;
      RECT  0.000000  84.660000  0.775000  84.730000 ;
      RECT  0.000000  84.730000  0.845000  84.800000 ;
      RECT  0.000000  84.800000  0.915000  84.825000 ;
      RECT  0.000000  84.825000  0.940000  95.065000 ;
      RECT  0.000000  95.065000  0.870000  95.135000 ;
      RECT  0.000000  95.135000  0.800000  95.205000 ;
      RECT  0.000000  95.205000  0.730000  95.275000 ;
      RECT  0.000000  95.275000  0.660000  95.345000 ;
      RECT  0.000000  95.345000  0.590000  95.415000 ;
      RECT  0.000000  95.415000  0.520000  95.485000 ;
      RECT  0.000000  95.485000  0.450000  95.555000 ;
      RECT  0.000000  95.555000  0.390000  95.615000 ;
      RECT  0.000000 101.700000 73.490000 104.845000 ;
      RECT  0.000000 104.845000 74.035000 125.160000 ;
      RECT  0.000000 130.500000 10.015000 130.570000 ;
      RECT  0.000000 130.570000  9.945000 130.640000 ;
      RECT  0.000000 130.640000  9.875000 130.710000 ;
      RECT  0.000000 130.710000  9.805000 130.780000 ;
      RECT  0.000000 130.780000  9.735000 130.850000 ;
      RECT  0.000000 130.850000  9.665000 130.920000 ;
      RECT  0.000000 130.920000  9.595000 130.990000 ;
      RECT  0.000000 130.990000  9.590000 130.995000 ;
      RECT  0.000000 145.410000  2.595000 146.420000 ;
      RECT  0.000000 146.420000 59.500000 199.490000 ;
      RECT  0.000000 146.420000 70.525000 146.425000 ;
      RECT  0.000000 146.420000 70.525000 195.970000 ;
      RECT  0.000000 146.425000 73.405000 195.970000 ;
      RECT  0.000000 146.425000 75.000000 174.220000 ;
      RECT  0.000000 174.220000 73.405000 175.420000 ;
      RECT  0.000000 175.420000 75.000000 195.970000 ;
      RECT  0.000000 195.970000 59.500000 199.490000 ;
      RECT  0.000000 199.490000 59.500000 200.000000 ;
      RECT  0.015000  96.385000  3.170000  96.455000 ;
      RECT  0.015000  96.385000  3.170000  96.455000 ;
      RECT  0.025000 137.990000  0.940000 138.060000 ;
      RECT  0.085000  96.315000  3.100000  96.385000 ;
      RECT  0.085000  96.315000  3.100000  96.385000 ;
      RECT  0.095000 137.920000  0.940000 137.990000 ;
      RECT  0.155000  96.245000  3.030000  96.315000 ;
      RECT  0.155000  96.245000  3.030000  96.315000 ;
      RECT  0.165000 137.850000  0.940000 137.920000 ;
      RECT  0.225000  96.175000  2.960000  96.245000 ;
      RECT  0.225000  96.175000  2.960000  96.245000 ;
      RECT  0.235000 137.780000  0.940000 137.850000 ;
      RECT  0.295000  96.105000  2.890000  96.175000 ;
      RECT  0.295000  96.105000  2.890000  96.175000 ;
      RECT  0.305000 137.710000  0.940000 137.780000 ;
      RECT  0.365000  96.035000  2.820000  96.105000 ;
      RECT  0.365000  96.035000  2.820000  96.105000 ;
      RECT  0.375000 137.640000  0.940000 137.710000 ;
      RECT  0.435000  95.965000  2.750000  96.035000 ;
      RECT  0.435000  95.965000  2.750000  96.035000 ;
      RECT  0.445000 137.570000  0.940000 137.640000 ;
      RECT  0.505000  95.895000  2.680000  95.965000 ;
      RECT  0.505000  95.895000  2.680000  95.965000 ;
      RECT  0.515000 137.500000  0.940000 137.570000 ;
      RECT  0.520000  95.880000  2.665000  95.895000 ;
      RECT  0.520000  95.880000  2.665000  95.895000 ;
      RECT  0.520000  95.880000  2.665000  95.895000 ;
      RECT  0.535000  95.865000  2.650000  95.880000 ;
      RECT  0.535000  95.865000  2.650000  95.880000 ;
      RECT  0.535000  95.865000  2.650000  95.880000 ;
      RECT  0.585000 137.430000  0.940000 137.500000 ;
      RECT  0.590000  95.810000  2.595000  95.865000 ;
      RECT  0.590000  95.810000  2.595000  95.865000 ;
      RECT  0.590000  95.810000  2.650000  95.865000 ;
      RECT  0.655000 137.360000  0.940000 137.430000 ;
      RECT  0.660000  95.740000  2.525000  95.810000 ;
      RECT  0.660000  95.740000  2.525000  95.810000 ;
      RECT  0.660000  95.740000  2.650000  95.810000 ;
      RECT  0.725000 137.290000  0.940000 137.360000 ;
      RECT  0.730000  95.670000  2.455000  95.740000 ;
      RECT  0.730000  95.670000  2.455000  95.740000 ;
      RECT  0.730000  95.670000  2.650000  95.740000 ;
      RECT  0.795000 137.220000  0.940000 137.290000 ;
      RECT  0.800000  95.600000  2.385000  95.670000 ;
      RECT  0.800000  95.600000  2.385000  95.670000 ;
      RECT  0.800000  95.600000  2.650000  95.670000 ;
      RECT  0.865000 137.150000  0.940000 137.220000 ;
      RECT  0.870000  95.530000  2.315000  95.600000 ;
      RECT  0.870000  95.530000  2.315000  95.600000 ;
      RECT  0.870000  95.530000  2.650000  95.600000 ;
      RECT  0.935000 137.080000  0.940000 137.150000 ;
      RECT  0.940000  95.460000  2.650000  95.530000 ;
      RECT  0.945000  95.460000  2.245000  95.530000 ;
      RECT  0.945000  95.460000  2.245000  95.530000 ;
      RECT  0.985000   0.240000 11.975000   0.590000 ;
      RECT  0.985000   0.590000  3.300000   0.660000 ;
      RECT  0.985000   0.660000  3.230000   0.730000 ;
      RECT  0.985000   0.730000  3.160000   0.800000 ;
      RECT  0.985000   0.800000  3.090000   0.870000 ;
      RECT  0.985000   0.870000  3.020000   0.940000 ;
      RECT  0.985000   0.940000  2.950000   1.010000 ;
      RECT  0.985000   1.010000  2.880000   1.080000 ;
      RECT  0.985000   1.080000  2.810000   1.150000 ;
      RECT  0.985000   1.150000  2.740000   1.220000 ;
      RECT  0.985000   1.220000  2.670000   1.290000 ;
      RECT  0.985000   1.290000  2.600000   1.360000 ;
      RECT  0.985000   1.360000  2.530000   1.430000 ;
      RECT  0.985000   1.430000  2.460000   1.500000 ;
      RECT  0.985000   1.500000  2.415000   1.545000 ;
      RECT  0.985000   1.545000  2.415000   3.150000 ;
      RECT  0.985000   3.150000  2.415000   3.220000 ;
      RECT  0.985000   3.220000  2.485000   3.290000 ;
      RECT  0.985000   3.290000  2.555000   3.360000 ;
      RECT  0.985000   3.360000  2.625000   3.430000 ;
      RECT  0.985000   3.430000  2.695000   3.500000 ;
      RECT  0.985000   3.500000  2.765000   3.570000 ;
      RECT  0.985000   3.570000  2.835000   3.640000 ;
      RECT  0.985000   3.640000  2.905000   3.710000 ;
      RECT  0.985000   3.710000  2.975000   3.780000 ;
      RECT  0.985000   3.780000  3.045000   3.850000 ;
      RECT  0.985000   3.850000  3.115000   3.920000 ;
      RECT  0.985000   3.920000  3.185000   3.990000 ;
      RECT  0.985000   3.990000  3.255000   4.060000 ;
      RECT  0.985000   4.060000  3.325000   4.105000 ;
      RECT  0.985000   4.105000  4.515000  71.340000 ;
      RECT  0.985000  71.910000 19.260000  79.760000 ;
      RECT  0.985000  80.435000 30.155000  84.475000 ;
      RECT  1.010000  95.390000  2.175000  95.460000 ;
      RECT  1.010000  95.390000  2.175000  95.460000 ;
      RECT  1.010000  95.390000  2.650000  95.460000 ;
      RECT  1.055000  84.475000  3.865000  84.545000 ;
      RECT  1.055000  84.475000  3.865000  84.545000 ;
      RECT  1.080000  95.320000  2.650000  95.390000 ;
      RECT  1.085000  95.320000  2.105000  95.390000 ;
      RECT  1.085000  95.320000  2.105000  95.390000 ;
      RECT  1.125000  84.545000  3.795000  84.615000 ;
      RECT  1.125000  84.545000  3.795000  84.615000 ;
      RECT  1.125000 130.995000 72.380000 131.065000 ;
      RECT  1.150000  95.250000  2.650000  95.320000 ;
      RECT  1.155000  95.250000  2.035000  95.320000 ;
      RECT  1.155000  95.250000  2.035000  95.320000 ;
      RECT  1.195000  84.615000  3.725000  84.685000 ;
      RECT  1.195000  84.615000  3.725000  84.685000 ;
      RECT  1.195000 131.065000 72.380000 131.135000 ;
      RECT  1.220000  81.705000  2.650000  85.760000 ;
      RECT  1.220000  84.685000  3.700000  84.710000 ;
      RECT  1.220000  84.685000  3.700000  84.710000 ;
      RECT  1.220000  84.710000  3.630000  84.780000 ;
      RECT  1.220000  84.780000  3.560000  84.850000 ;
      RECT  1.220000  84.850000  3.490000  84.920000 ;
      RECT  1.220000  84.920000  3.420000  84.990000 ;
      RECT  1.220000  84.990000  3.350000  85.060000 ;
      RECT  1.220000  85.060000  3.280000  85.130000 ;
      RECT  1.220000  85.130000  3.210000  85.200000 ;
      RECT  1.220000  85.200000  3.140000  85.270000 ;
      RECT  1.220000  85.270000  3.070000  85.340000 ;
      RECT  1.220000  85.340000  3.000000  85.410000 ;
      RECT  1.220000  85.410000  2.930000  85.480000 ;
      RECT  1.220000  85.480000  2.860000  85.550000 ;
      RECT  1.220000  85.550000  2.790000  85.620000 ;
      RECT  1.220000  85.620000  2.720000  85.690000 ;
      RECT  1.220000  85.690000  2.650000  85.760000 ;
      RECT  1.220000  85.760000  2.580000  85.830000 ;
      RECT  1.220000  85.760000  2.580000  85.830000 ;
      RECT  1.220000  85.830000  2.510000  85.900000 ;
      RECT  1.220000  85.830000  2.510000  85.900000 ;
      RECT  1.220000  85.900000  2.440000  85.970000 ;
      RECT  1.220000  85.900000  2.440000  85.970000 ;
      RECT  1.220000  85.970000  2.370000  86.040000 ;
      RECT  1.220000  85.970000  2.370000  86.040000 ;
      RECT  1.220000  86.040000  2.300000  86.110000 ;
      RECT  1.220000  86.040000  2.300000  86.110000 ;
      RECT  1.220000  86.110000  2.230000  86.180000 ;
      RECT  1.220000  86.110000  2.230000  86.180000 ;
      RECT  1.220000  86.180000  2.160000  86.250000 ;
      RECT  1.220000  86.180000  2.160000  86.250000 ;
      RECT  1.220000  86.250000  2.090000  86.320000 ;
      RECT  1.220000  86.250000  2.090000  86.320000 ;
      RECT  1.220000  86.320000  2.020000  86.390000 ;
      RECT  1.220000  86.320000  2.020000  86.390000 ;
      RECT  1.220000  86.390000  1.950000  86.460000 ;
      RECT  1.220000  86.390000  1.950000  86.460000 ;
      RECT  1.220000  86.460000  1.880000  86.530000 ;
      RECT  1.220000  86.460000  1.880000  86.530000 ;
      RECT  1.220000  86.530000  1.810000  86.600000 ;
      RECT  1.220000  86.530000  1.810000  86.600000 ;
      RECT  1.220000  86.600000  1.740000  86.670000 ;
      RECT  1.220000  86.600000  1.740000  86.670000 ;
      RECT  1.220000  86.670000  1.670000  86.740000 ;
      RECT  1.220000  86.670000  1.670000  86.740000 ;
      RECT  1.220000  86.740000  1.600000  86.810000 ;
      RECT  1.220000  86.740000  1.600000  86.810000 ;
      RECT  1.220000  86.810000  1.530000  86.880000 ;
      RECT  1.220000  86.810000  1.530000  86.880000 ;
      RECT  1.220000  86.880000  1.460000  86.950000 ;
      RECT  1.220000  86.880000  1.460000  86.950000 ;
      RECT  1.220000  86.950000  1.390000  87.020000 ;
      RECT  1.220000  86.950000  1.390000  87.020000 ;
      RECT  1.220000  87.020000  1.320000  87.090000 ;
      RECT  1.220000  87.020000  1.320000  87.090000 ;
      RECT  1.220000  87.090000  1.250000  87.160000 ;
      RECT  1.220000  87.090000  1.250000  87.160000 ;
      RECT  1.220000  87.190000  2.650000  94.810000 ;
      RECT  1.220000  94.810000  1.525000  94.880000 ;
      RECT  1.220000  94.880000  1.455000  94.950000 ;
      RECT  1.220000  94.950000  1.385000  95.020000 ;
      RECT  1.220000  95.020000  1.315000  95.090000 ;
      RECT  1.220000  95.090000  1.245000  95.160000 ;
      RECT  1.220000  95.160000  1.225000  95.180000 ;
      RECT  1.220000  95.180000  2.650000  95.250000 ;
      RECT  1.220000 135.750000 14.920000 139.225000 ;
      RECT  1.220000 137.195000 70.400000 137.265000 ;
      RECT  1.220000 137.195000 70.400000 137.265000 ;
      RECT  1.220000 137.265000 70.330000 137.335000 ;
      RECT  1.220000 137.265000 70.330000 137.335000 ;
      RECT  1.220000 137.335000 70.260000 137.405000 ;
      RECT  1.220000 137.335000 70.260000 137.405000 ;
      RECT  1.220000 137.405000 70.190000 137.475000 ;
      RECT  1.220000 137.405000 70.190000 137.475000 ;
      RECT  1.220000 137.475000 70.120000 137.545000 ;
      RECT  1.220000 137.475000 70.120000 137.545000 ;
      RECT  1.220000 137.545000 70.050000 137.615000 ;
      RECT  1.220000 137.545000 70.050000 137.615000 ;
      RECT  1.220000 137.615000 69.980000 137.685000 ;
      RECT  1.220000 137.615000 69.980000 137.685000 ;
      RECT  1.220000 137.685000 69.910000 137.755000 ;
      RECT  1.220000 137.685000 69.910000 137.755000 ;
      RECT  1.220000 137.755000 69.840000 137.825000 ;
      RECT  1.220000 137.755000 69.840000 137.825000 ;
      RECT  1.220000 137.825000 69.770000 137.895000 ;
      RECT  1.220000 137.825000 69.770000 137.895000 ;
      RECT  1.220000 137.895000 69.700000 137.965000 ;
      RECT  1.220000 137.895000 69.700000 137.965000 ;
      RECT  1.220000 137.965000 69.630000 138.035000 ;
      RECT  1.220000 137.965000 69.630000 138.035000 ;
      RECT  1.220000 138.035000 69.560000 138.105000 ;
      RECT  1.220000 138.035000 69.560000 138.105000 ;
      RECT  1.220000 138.105000 69.490000 138.175000 ;
      RECT  1.220000 138.105000 69.490000 138.175000 ;
      RECT  1.220000 138.175000 69.420000 138.245000 ;
      RECT  1.220000 138.175000 69.420000 138.245000 ;
      RECT  1.220000 138.245000 69.350000 138.315000 ;
      RECT  1.220000 138.245000 69.350000 138.315000 ;
      RECT  1.220000 138.315000 69.280000 138.385000 ;
      RECT  1.220000 138.315000 69.280000 138.385000 ;
      RECT  1.220000 138.385000 69.210000 138.455000 ;
      RECT  1.220000 138.385000 69.210000 138.455000 ;
      RECT  1.220000 138.455000 69.140000 138.525000 ;
      RECT  1.220000 138.455000 69.140000 138.525000 ;
      RECT  1.220000 138.525000 69.070000 138.595000 ;
      RECT  1.220000 138.525000 69.070000 138.595000 ;
      RECT  1.220000 138.595000 69.000000 138.665000 ;
      RECT  1.220000 138.595000 69.000000 138.665000 ;
      RECT  1.220000 138.665000 16.790000 138.685000 ;
      RECT  1.220000 138.665000 16.790000 138.685000 ;
      RECT  1.220000 138.685000 16.770000 138.705000 ;
      RECT  1.220000 138.685000 16.770000 138.705000 ;
      RECT  1.220000 138.705000 16.765000 138.710000 ;
      RECT  1.220000 138.705000 16.765000 138.710000 ;
      RECT  1.220000 138.710000 14.920000 138.900000 ;
      RECT  1.220000 140.480000 70.225000 140.550000 ;
      RECT  1.220000 140.550000 70.295000 140.620000 ;
      RECT  1.220000 140.620000 70.365000 140.690000 ;
      RECT  1.220000 140.690000 70.435000 140.760000 ;
      RECT  1.220000 140.760000 70.505000 140.780000 ;
      RECT  1.220000 140.780000 70.525000 141.095000 ;
      RECT  1.225000  95.180000  1.965000  95.250000 ;
      RECT  1.225000  95.180000  1.965000  95.250000 ;
      RECT  1.245000  95.160000  1.945000  95.180000 ;
      RECT  1.245000  95.160000  1.945000  95.180000 ;
      RECT  1.265000 131.135000 72.380000 131.205000 ;
      RECT  1.265000 137.150000 70.470000 137.195000 ;
      RECT  1.265000 137.150000 70.470000 137.195000 ;
      RECT  1.290000 138.900000 14.920000 138.970000 ;
      RECT  1.290000 138.900000 14.920000 138.970000 ;
      RECT  1.290000 140.410000 70.155000 140.480000 ;
      RECT  1.315000  95.090000  1.875000  95.160000 ;
      RECT  1.315000  95.090000  1.875000  95.160000 ;
      RECT  1.335000 131.205000 72.380000 131.275000 ;
      RECT  1.335000 137.080000 70.515000 137.150000 ;
      RECT  1.335000 137.080000 70.515000 137.150000 ;
      RECT  1.340000 141.375000 69.645000 143.595000 ;
      RECT  1.360000 138.970000 14.920000 139.040000 ;
      RECT  1.360000 138.970000 14.920000 139.040000 ;
      RECT  1.360000 140.340000 70.085000 140.410000 ;
      RECT  1.385000  95.020000  1.805000  95.090000 ;
      RECT  1.385000  95.020000  1.805000  95.090000 ;
      RECT  1.405000 131.275000 72.380000 131.345000 ;
      RECT  1.405000 137.010000 70.585000 137.080000 ;
      RECT  1.405000 137.010000 70.585000 137.080000 ;
      RECT  1.430000 139.040000 14.920000 139.110000 ;
      RECT  1.430000 139.040000 14.920000 139.110000 ;
      RECT  1.430000 140.270000 70.015000 140.340000 ;
      RECT  1.455000  94.950000  1.735000  95.020000 ;
      RECT  1.455000  94.950000  1.735000  95.020000 ;
      RECT  1.475000 131.345000 72.380000 131.415000 ;
      RECT  1.475000 136.940000 70.655000 137.010000 ;
      RECT  1.475000 136.940000 70.655000 137.010000 ;
      RECT  1.500000 139.110000 14.920000 139.180000 ;
      RECT  1.500000 139.110000 14.920000 139.180000 ;
      RECT  1.500000 140.200000 69.945000 140.270000 ;
      RECT  1.525000  94.880000  1.665000  94.950000 ;
      RECT  1.525000  94.880000  1.665000  94.950000 ;
      RECT  1.545000 131.415000 72.380000 131.485000 ;
      RECT  1.545000 136.870000 70.725000 136.940000 ;
      RECT  1.545000 136.870000 70.725000 136.940000 ;
      RECT  1.545000 139.180000 14.920000 139.225000 ;
      RECT  1.545000 139.180000 14.920000 139.225000 ;
      RECT  1.570000 140.130000 69.875000 140.200000 ;
      RECT  1.615000 131.485000 72.380000 131.555000 ;
      RECT  1.615000 136.800000 70.795000 136.870000 ;
      RECT  1.615000 136.800000 70.795000 136.870000 ;
      RECT  1.640000 143.875000 70.525000 143.945000 ;
      RECT  1.665000  94.810000  2.650000  94.880000 ;
      RECT  1.685000 131.555000 72.380000 131.625000 ;
      RECT  1.685000 136.730000 70.865000 136.800000 ;
      RECT  1.685000 136.730000 70.865000 136.800000 ;
      RECT  1.710000 143.945000 70.525000 144.015000 ;
      RECT  1.735000  94.880000  2.650000  94.950000 ;
      RECT  1.755000 131.625000 72.380000 131.695000 ;
      RECT  1.755000 136.660000 70.935000 136.730000 ;
      RECT  1.755000 136.660000 70.935000 136.730000 ;
      RECT  1.780000 144.015000 70.525000 144.085000 ;
      RECT  1.805000  94.950000  2.650000  95.020000 ;
      RECT  1.825000 131.695000 72.380000 131.765000 ;
      RECT  1.825000 136.590000 71.005000 136.660000 ;
      RECT  1.825000 136.590000 71.005000 136.660000 ;
      RECT  1.850000 144.085000 70.525000 144.155000 ;
      RECT  1.875000  95.020000  2.650000  95.090000 ;
      RECT  1.895000 131.765000 72.380000 131.835000 ;
      RECT  1.895000 136.520000 71.075000 136.590000 ;
      RECT  1.895000 136.520000 71.075000 136.590000 ;
      RECT  1.920000 144.155000 70.525000 144.225000 ;
      RECT  1.945000  95.090000  2.650000  95.160000 ;
      RECT  1.965000  95.160000  2.650000  95.180000 ;
      RECT  1.965000 131.835000 72.380000 131.905000 ;
      RECT  1.965000 136.450000 71.145000 136.520000 ;
      RECT  1.965000 136.450000 71.145000 136.520000 ;
      RECT  1.980000 144.225000 70.525000 144.285000 ;
      RECT  2.035000 131.905000 72.380000 131.975000 ;
      RECT  2.035000 136.380000 71.215000 136.450000 ;
      RECT  2.035000 136.380000 71.215000 136.450000 ;
      RECT  2.050000 144.285000 70.455000 144.355000 ;
      RECT  2.105000 131.975000 72.380000 132.045000 ;
      RECT  2.105000 136.310000 71.285000 136.380000 ;
      RECT  2.105000 136.310000 71.285000 136.380000 ;
      RECT  2.120000 144.355000 70.385000 144.425000 ;
      RECT  2.175000 132.045000 72.380000 132.115000 ;
      RECT  2.175000 136.240000 71.355000 136.310000 ;
      RECT  2.175000 136.240000 71.355000 136.310000 ;
      RECT  2.190000 144.425000 70.315000 144.495000 ;
      RECT  2.245000 132.115000 72.380000 132.185000 ;
      RECT  2.245000 136.170000 71.425000 136.240000 ;
      RECT  2.245000 136.170000 71.425000 136.240000 ;
      RECT  2.260000 144.495000 70.245000 144.565000 ;
      RECT  2.315000 132.185000 72.380000 132.255000 ;
      RECT  2.315000 136.100000 71.495000 136.170000 ;
      RECT  2.315000 136.100000 71.495000 136.170000 ;
      RECT  2.330000 144.565000 70.175000 144.635000 ;
      RECT  2.385000 132.255000 72.380000 132.325000 ;
      RECT  2.385000 136.030000 71.565000 136.100000 ;
      RECT  2.385000 136.030000 71.565000 136.100000 ;
      RECT  2.400000 144.635000 70.105000 144.705000 ;
      RECT  2.455000 132.325000 72.380000 132.395000 ;
      RECT  2.455000 135.960000 71.635000 136.030000 ;
      RECT  2.455000 135.960000 71.635000 136.030000 ;
      RECT  2.470000 144.705000 70.035000 144.775000 ;
      RECT  2.475000 132.740000 13.110000 132.810000 ;
      RECT  2.520000 132.395000 72.380000 132.460000 ;
      RECT  2.525000 135.890000 71.705000 135.960000 ;
      RECT  2.525000 135.890000 71.705000 135.960000 ;
      RECT  2.540000 144.775000 69.965000 144.845000 ;
      RECT  2.545000 132.810000 13.110000 132.880000 ;
      RECT  2.545000 144.845000 69.960000 144.850000 ;
      RECT  2.580000 135.440000 13.110000 135.470000 ;
      RECT  2.595000 135.820000 71.775000 135.890000 ;
      RECT  2.595000 135.820000 71.775000 135.890000 ;
      RECT  2.615000 132.880000 13.110000 132.950000 ;
      RECT  2.650000 135.370000 13.110000 135.440000 ;
      RECT  2.665000 135.750000 71.845000 135.820000 ;
      RECT  2.665000 135.750000 71.845000 135.820000 ;
      RECT  2.685000 132.950000 13.110000 133.020000 ;
      RECT  2.695000   1.660000  3.625000   3.035000 ;
      RECT  2.715000   1.640000  3.625000   1.660000 ;
      RECT  2.720000 135.300000 13.110000 135.370000 ;
      RECT  2.755000 133.020000 13.110000 133.090000 ;
      RECT  2.765000   3.035000  3.625000   3.105000 ;
      RECT  2.785000   1.570000  3.625000   1.640000 ;
      RECT  2.790000 135.230000 13.110000 135.300000 ;
      RECT  2.825000 133.090000 13.110000 133.160000 ;
      RECT  2.835000   3.105000  3.625000   3.175000 ;
      RECT  2.855000   1.500000  3.625000   1.570000 ;
      RECT  2.860000 135.160000 13.110000 135.230000 ;
      RECT  2.875000 145.130000  5.945000 146.140000 ;
      RECT  2.895000 133.160000 13.110000 133.230000 ;
      RECT  2.905000   3.175000  3.625000   3.245000 ;
      RECT  2.925000   1.430000  3.625000   1.500000 ;
      RECT  2.930000  85.875000 71.475000  94.750000 ;
      RECT  2.930000  94.750000 75.000000  95.615000 ;
      RECT  2.930000  95.615000 73.545000  95.680000 ;
      RECT  2.930000  95.680000 73.480000  95.745000 ;
      RECT  2.930000  95.745000 73.475000  95.750000 ;
      RECT  2.930000 135.090000 13.110000 135.160000 ;
      RECT  2.965000 133.230000 13.110000 133.300000 ;
      RECT  2.970000  85.835000 71.475000  85.875000 ;
      RECT  2.970000  85.835000 71.475000  85.875000 ;
      RECT  2.975000   3.245000  3.625000   3.315000 ;
      RECT  2.995000   1.360000  3.625000   1.430000 ;
      RECT  3.000000  95.750000 71.475000  95.820000 ;
      RECT  3.000000  95.750000 71.475000  95.820000 ;
      RECT  3.000000  95.750000 73.405000  95.820000 ;
      RECT  3.000000 135.020000 13.110000 135.090000 ;
      RECT  3.035000 133.300000 13.110000 133.370000 ;
      RECT  3.040000  85.765000 71.475000  85.835000 ;
      RECT  3.040000  85.765000 71.475000  85.835000 ;
      RECT  3.045000   3.315000  3.625000   3.385000 ;
      RECT  3.065000   1.290000  3.625000   1.360000 ;
      RECT  3.070000  95.820000 71.475000  95.890000 ;
      RECT  3.070000  95.820000 71.475000  95.890000 ;
      RECT  3.070000  95.820000 73.335000  95.890000 ;
      RECT  3.070000 134.950000 13.110000 135.020000 ;
      RECT  3.090000   3.385000  3.625000   3.430000 ;
      RECT  3.105000 133.370000 13.110000 133.440000 ;
      RECT  3.110000  85.695000 71.475000  85.765000 ;
      RECT  3.110000  85.695000 71.475000  85.765000 ;
      RECT  3.135000   1.220000  3.625000   1.290000 ;
      RECT  3.140000  95.890000 71.475000  95.960000 ;
      RECT  3.140000  95.890000 71.475000  95.960000 ;
      RECT  3.140000  95.890000 73.265000  95.960000 ;
      RECT  3.140000 134.880000 13.110000 134.950000 ;
      RECT  3.160000   3.430000 12.005000   3.500000 ;
      RECT  3.175000 133.440000 13.110000 133.510000 ;
      RECT  3.180000  85.625000 71.475000  85.695000 ;
      RECT  3.180000  85.625000 71.475000  85.695000 ;
      RECT  3.205000   1.150000  3.625000   1.220000 ;
      RECT  3.210000  95.960000 71.475000  96.030000 ;
      RECT  3.210000  95.960000 71.475000  96.030000 ;
      RECT  3.210000  95.960000 73.195000  96.030000 ;
      RECT  3.210000 134.810000 13.110000 134.880000 ;
      RECT  3.230000   3.500000 12.005000   3.570000 ;
      RECT  3.245000 133.510000 13.110000 133.580000 ;
      RECT  3.250000  85.555000 71.475000  85.625000 ;
      RECT  3.250000  85.555000 71.475000  85.625000 ;
      RECT  3.260000  85.545000 71.475000  85.555000 ;
      RECT  3.260000  85.545000 71.475000  85.555000 ;
      RECT  3.260000  85.545000 75.000000  85.555000 ;
      RECT  3.275000   1.080000  3.625000   1.150000 ;
      RECT  3.280000  96.030000 71.475000  96.100000 ;
      RECT  3.280000  96.030000 71.475000  96.100000 ;
      RECT  3.280000  96.030000 73.125000  96.100000 ;
      RECT  3.280000 134.740000 13.110000 134.810000 ;
      RECT  3.300000   3.570000 12.005000   3.640000 ;
      RECT  3.315000 133.580000 13.110000 133.650000 ;
      RECT  3.330000  85.475000 71.475000  85.545000 ;
      RECT  3.330000  85.475000 71.475000  85.545000 ;
      RECT  3.330000  85.475000 75.000000  85.545000 ;
      RECT  3.345000   1.010000  3.625000   1.080000 ;
      RECT  3.350000  96.100000 71.475000  96.170000 ;
      RECT  3.350000  96.100000 71.475000  96.170000 ;
      RECT  3.350000  96.100000 73.055000  96.170000 ;
      RECT  3.350000 134.670000 13.110000 134.740000 ;
      RECT  3.370000   3.640000 12.005000   3.710000 ;
      RECT  3.385000 133.650000 13.110000 133.720000 ;
      RECT  3.400000  85.405000 71.475000  85.475000 ;
      RECT  3.400000  85.405000 71.475000  85.475000 ;
      RECT  3.400000  85.405000 75.000000  85.475000 ;
      RECT  3.415000   0.940000  3.625000   1.010000 ;
      RECT  3.420000  96.170000 71.475000  96.240000 ;
      RECT  3.420000  96.170000 71.475000  96.240000 ;
      RECT  3.420000  96.170000 72.985000  96.240000 ;
      RECT  3.420000 134.600000 13.110000 134.670000 ;
      RECT  3.440000   3.710000 12.005000   3.780000 ;
      RECT  3.455000 133.720000 13.110000 133.790000 ;
      RECT  3.470000  85.335000 71.475000  85.405000 ;
      RECT  3.470000  85.335000 71.475000  85.405000 ;
      RECT  3.470000  85.335000 75.000000  85.405000 ;
      RECT  3.485000   0.870000  3.625000   0.940000 ;
      RECT  3.485000   3.780000 12.005000   3.825000 ;
      RECT  3.490000  85.315000 33.105000  85.335000 ;
      RECT  3.490000  85.315000 33.105000  85.335000 ;
      RECT  3.490000  96.240000 71.475000  96.310000 ;
      RECT  3.490000  96.240000 71.475000  96.310000 ;
      RECT  3.490000  96.240000 72.915000  96.310000 ;
      RECT  3.490000 134.530000 13.110000 134.600000 ;
      RECT  3.525000 133.790000 13.110000 133.860000 ;
      RECT  3.560000  85.245000 33.105000  85.315000 ;
      RECT  3.560000  85.245000 33.105000  85.315000 ;
      RECT  3.560000  96.310000 71.475000  96.380000 ;
      RECT  3.560000  96.310000 71.475000  96.380000 ;
      RECT  3.560000  96.310000 72.845000  96.380000 ;
      RECT  3.560000 134.460000 13.110000 134.530000 ;
      RECT  3.595000 133.860000 13.110000 133.930000 ;
      RECT  3.630000  85.175000 33.105000  85.245000 ;
      RECT  3.630000  85.175000 33.105000  85.245000 ;
      RECT  3.630000  96.380000 71.475000  96.450000 ;
      RECT  3.630000  96.380000 71.475000  96.450000 ;
      RECT  3.630000  96.380000 72.775000  96.450000 ;
      RECT  3.635000 134.390000 13.110000 134.460000 ;
      RECT  3.665000 133.930000 13.110000 134.000000 ;
      RECT  3.700000  85.105000 33.105000  85.175000 ;
      RECT  3.700000  85.105000 33.105000  85.175000 ;
      RECT  3.700000  96.450000 71.475000  96.520000 ;
      RECT  3.700000  96.450000 71.475000  96.520000 ;
      RECT  3.700000  96.450000 72.705000  96.520000 ;
      RECT  3.700000 134.320000 13.110000 134.390000 ;
      RECT  3.735000 134.000000 13.110000 134.070000 ;
      RECT  3.770000  85.035000 33.105000  85.105000 ;
      RECT  3.770000  85.035000 33.105000  85.105000 ;
      RECT  3.770000  96.520000 71.475000  96.590000 ;
      RECT  3.770000  96.520000 71.475000  96.590000 ;
      RECT  3.770000  96.520000 72.635000  96.590000 ;
      RECT  3.775000 134.250000 13.110000 134.320000 ;
      RECT  3.805000 134.070000 13.110000 134.140000 ;
      RECT  3.840000  84.965000 33.105000  85.035000 ;
      RECT  3.840000  84.965000 33.105000  85.035000 ;
      RECT  3.840000  96.590000 71.475000  96.660000 ;
      RECT  3.840000  96.590000 71.475000  96.660000 ;
      RECT  3.840000  96.590000 72.565000  96.660000 ;
      RECT  3.845000 134.140000 13.110000 134.180000 ;
      RECT  3.845000 134.180000 13.110000 134.250000 ;
      RECT  3.905000   1.140000  5.710000   3.150000 ;
      RECT  3.910000  84.895000 33.105000  84.965000 ;
      RECT  3.910000  84.895000 33.105000  84.965000 ;
      RECT  3.910000  96.660000 71.475000  96.730000 ;
      RECT  3.910000  96.660000 71.475000  96.730000 ;
      RECT  3.910000  96.660000 72.495000  96.730000 ;
      RECT  3.980000  84.825000 33.105000  84.895000 ;
      RECT  3.980000  84.825000 33.105000  84.895000 ;
      RECT  3.980000  96.730000 71.475000  96.800000 ;
      RECT  3.980000  96.730000 71.475000  96.800000 ;
      RECT  3.980000  96.730000 72.425000  96.800000 ;
      RECT  4.050000  84.755000 33.105000  84.825000 ;
      RECT  4.050000  84.755000 33.105000  84.825000 ;
      RECT  4.050000  96.800000 71.475000  96.870000 ;
      RECT  4.050000  96.800000 71.475000  96.870000 ;
      RECT  4.050000  96.800000 72.355000  96.870000 ;
      RECT  4.120000  96.870000 71.475000  96.940000 ;
      RECT  4.120000  96.870000 71.475000  96.940000 ;
      RECT  4.120000  96.870000 72.285000  96.940000 ;
      RECT  4.190000  96.940000 71.475000  97.010000 ;
      RECT  4.190000  96.940000 71.475000  97.010000 ;
      RECT  4.190000  96.940000 72.215000  97.010000 ;
      RECT  4.260000  97.010000 71.475000  97.080000 ;
      RECT  4.260000  97.010000 71.475000  97.080000 ;
      RECT  4.260000  97.010000 72.145000  97.080000 ;
      RECT  4.330000  97.080000 71.475000  97.150000 ;
      RECT  4.330000  97.080000 71.475000  97.150000 ;
      RECT  4.330000  97.080000 72.075000  97.150000 ;
      RECT  4.400000  97.150000 71.475000  97.220000 ;
      RECT  4.400000  97.150000 71.475000  97.220000 ;
      RECT  4.400000  97.150000 72.005000  97.220000 ;
      RECT  4.430000  97.220000 71.475000  97.250000 ;
      RECT  4.430000  97.220000 71.475000  97.250000 ;
      RECT  4.430000  97.220000 71.975000  97.250000 ;
      RECT  4.795000   3.430000 12.005000   3.825000 ;
      RECT  4.795000   3.825000 12.005000   6.380000 ;
      RECT  4.795000   6.380000 11.935000   6.450000 ;
      RECT  4.795000   6.380000 11.935000   6.450000 ;
      RECT  4.795000   6.450000 11.865000   6.520000 ;
      RECT  4.795000   6.450000 11.865000   6.520000 ;
      RECT  4.795000   6.520000 11.795000   6.590000 ;
      RECT  4.795000   6.520000 11.795000   6.590000 ;
      RECT  4.795000   6.590000 11.725000   6.660000 ;
      RECT  4.795000   6.590000 11.725000   6.660000 ;
      RECT  4.795000   6.660000 11.655000   6.730000 ;
      RECT  4.795000   6.660000 11.655000   6.730000 ;
      RECT  4.795000   6.730000 11.585000   6.800000 ;
      RECT  4.795000   6.730000 11.585000   6.800000 ;
      RECT  4.795000   6.800000 11.515000   6.870000 ;
      RECT  4.795000   6.800000 11.515000   6.870000 ;
      RECT  4.795000   6.870000 11.445000   6.940000 ;
      RECT  4.795000   6.870000 11.445000   6.940000 ;
      RECT  4.795000   6.940000 11.440000   6.945000 ;
      RECT  4.795000   6.940000 11.440000   6.945000 ;
      RECT  4.795000   6.945000 12.090000   7.040000 ;
      RECT  4.795000   7.040000 12.090000   7.110000 ;
      RECT  4.795000   7.040000 12.090000   7.110000 ;
      RECT  4.795000   7.110000 12.160000   7.180000 ;
      RECT  4.795000   7.110000 12.160000   7.180000 ;
      RECT  4.795000   7.180000 12.230000   7.250000 ;
      RECT  4.795000   7.180000 12.230000   7.250000 ;
      RECT  4.795000   7.250000 12.300000   7.320000 ;
      RECT  4.795000   7.250000 12.300000   7.320000 ;
      RECT  4.795000   7.320000 12.370000   7.365000 ;
      RECT  4.795000   7.320000 12.370000   7.365000 ;
      RECT  4.795000   7.365000 12.415000  10.510000 ;
      RECT  4.795000   7.365000 12.415000  12.455000 ;
      RECT  4.795000   7.365000 12.415000  12.455000 ;
      RECT  4.795000  10.510000 12.520000  10.585000 ;
      RECT  4.795000  10.585000 14.275000  12.455000 ;
      RECT  4.795000  10.585000 14.275000  16.200000 ;
      RECT  4.795000  12.455000 14.275000  12.525000 ;
      RECT  4.795000  12.455000 14.275000  12.525000 ;
      RECT  4.795000  12.525000 14.345000  12.595000 ;
      RECT  4.795000  12.525000 14.345000  12.595000 ;
      RECT  4.795000  12.595000 14.415000  12.665000 ;
      RECT  4.795000  12.595000 14.415000  12.665000 ;
      RECT  4.795000  12.665000 14.485000  12.735000 ;
      RECT  4.795000  12.665000 14.485000  12.735000 ;
      RECT  4.795000  12.735000 14.555000  12.805000 ;
      RECT  4.795000  12.735000 14.555000  12.805000 ;
      RECT  4.795000  12.805000 14.625000  12.875000 ;
      RECT  4.795000  12.805000 14.625000  12.875000 ;
      RECT  4.795000  12.875000 14.695000  12.945000 ;
      RECT  4.795000  12.875000 14.695000  12.945000 ;
      RECT  4.795000  12.945000 14.765000  13.015000 ;
      RECT  4.795000  12.945000 14.765000  13.015000 ;
      RECT  4.795000  13.015000 14.835000  13.085000 ;
      RECT  4.795000  13.015000 14.835000  13.085000 ;
      RECT  4.795000  13.085000 14.905000  13.155000 ;
      RECT  4.795000  13.085000 14.905000  13.155000 ;
      RECT  4.795000  13.155000 14.975000  13.225000 ;
      RECT  4.795000  13.155000 14.975000  13.225000 ;
      RECT  4.795000  13.225000 15.045000  13.295000 ;
      RECT  4.795000  13.225000 15.045000  13.295000 ;
      RECT  4.795000  13.295000 15.115000  13.365000 ;
      RECT  4.795000  13.295000 15.115000  13.365000 ;
      RECT  4.795000  13.365000 15.185000  13.435000 ;
      RECT  4.795000  13.365000 15.185000  13.435000 ;
      RECT  4.795000  13.435000 15.255000  13.505000 ;
      RECT  4.795000  13.435000 15.255000  13.505000 ;
      RECT  4.795000  13.505000 15.325000  13.575000 ;
      RECT  4.795000  13.505000 15.325000  13.575000 ;
      RECT  4.795000  13.575000 15.395000  13.645000 ;
      RECT  4.795000  13.575000 15.395000  13.645000 ;
      RECT  4.795000  13.645000 15.465000  13.715000 ;
      RECT  4.795000  13.645000 15.465000  13.715000 ;
      RECT  4.795000  13.715000 15.535000  13.785000 ;
      RECT  4.795000  13.715000 15.535000  13.785000 ;
      RECT  4.795000  13.785000 15.605000  13.855000 ;
      RECT  4.795000  13.785000 15.605000  13.855000 ;
      RECT  4.795000  13.855000 15.675000  13.925000 ;
      RECT  4.795000  13.855000 15.675000  13.925000 ;
      RECT  4.795000  13.925000 15.745000  13.995000 ;
      RECT  4.795000  13.925000 15.745000  13.995000 ;
      RECT  4.795000  13.995000 15.815000  14.065000 ;
      RECT  4.795000  13.995000 15.815000  14.065000 ;
      RECT  4.795000  14.065000 15.885000  14.135000 ;
      RECT  4.795000  14.065000 15.885000  14.135000 ;
      RECT  4.795000  14.135000 15.955000  14.205000 ;
      RECT  4.795000  14.135000 15.955000  14.205000 ;
      RECT  4.795000  14.205000 16.025000  14.275000 ;
      RECT  4.795000  14.205000 16.025000  14.275000 ;
      RECT  4.795000  14.275000 16.095000  14.345000 ;
      RECT  4.795000  14.275000 16.095000  14.345000 ;
      RECT  4.795000  14.345000 16.165000  14.415000 ;
      RECT  4.795000  14.345000 16.165000  14.415000 ;
      RECT  4.795000  14.415000 16.235000  14.485000 ;
      RECT  4.795000  14.415000 16.235000  14.485000 ;
      RECT  4.795000  14.485000 16.305000  14.555000 ;
      RECT  4.795000  14.485000 16.305000  14.555000 ;
      RECT  4.795000  14.555000 16.375000  14.625000 ;
      RECT  4.795000  14.555000 16.375000  14.625000 ;
      RECT  4.795000  14.625000 16.445000  14.695000 ;
      RECT  4.795000  14.625000 16.445000  14.695000 ;
      RECT  4.795000  14.695000 16.515000  14.765000 ;
      RECT  4.795000  14.695000 16.515000  14.765000 ;
      RECT  4.795000  14.765000 16.585000  14.835000 ;
      RECT  4.795000  14.765000 16.585000  14.835000 ;
      RECT  4.795000  14.835000 16.655000  14.905000 ;
      RECT  4.795000  14.835000 16.655000  14.905000 ;
      RECT  4.795000  14.905000 16.725000  14.975000 ;
      RECT  4.795000  14.905000 16.725000  14.975000 ;
      RECT  4.795000  14.975000 16.795000  15.045000 ;
      RECT  4.795000  14.975000 16.795000  15.045000 ;
      RECT  4.795000  15.045000 16.865000  15.115000 ;
      RECT  4.795000  15.045000 16.865000  15.115000 ;
      RECT  4.795000  15.115000 16.935000  15.185000 ;
      RECT  4.795000  15.115000 16.935000  15.185000 ;
      RECT  4.795000  15.185000 17.005000  15.255000 ;
      RECT  4.795000  15.185000 17.005000  15.255000 ;
      RECT  4.795000  15.255000 17.075000  15.325000 ;
      RECT  4.795000  15.255000 17.075000  15.325000 ;
      RECT  4.795000  15.325000 17.145000  15.395000 ;
      RECT  4.795000  15.325000 17.145000  15.395000 ;
      RECT  4.795000  15.395000 17.215000  15.465000 ;
      RECT  4.795000  15.395000 17.215000  15.465000 ;
      RECT  4.795000  15.465000 17.285000  15.535000 ;
      RECT  4.795000  15.465000 17.285000  15.535000 ;
      RECT  4.795000  15.535000 17.355000  15.605000 ;
      RECT  4.795000  15.535000 17.355000  15.605000 ;
      RECT  4.795000  15.605000 17.425000  15.675000 ;
      RECT  4.795000  15.605000 17.425000  15.675000 ;
      RECT  4.795000  15.675000 17.495000  15.745000 ;
      RECT  4.795000  15.675000 17.495000  15.745000 ;
      RECT  4.795000  15.745000 17.565000  15.815000 ;
      RECT  4.795000  15.745000 17.565000  15.815000 ;
      RECT  4.795000  15.815000 17.635000  15.885000 ;
      RECT  4.795000  15.815000 17.635000  15.885000 ;
      RECT  4.795000  15.885000 17.705000  15.955000 ;
      RECT  4.795000  15.885000 17.705000  15.955000 ;
      RECT  4.795000  15.955000 17.775000  16.025000 ;
      RECT  4.795000  15.955000 17.775000  16.025000 ;
      RECT  4.795000  16.025000 17.845000  16.095000 ;
      RECT  4.795000  16.025000 17.845000  16.095000 ;
      RECT  4.795000  16.095000 17.915000  16.165000 ;
      RECT  4.795000  16.095000 17.915000  16.165000 ;
      RECT  4.795000  16.165000 17.985000  16.200000 ;
      RECT  4.795000  16.165000 17.985000  16.200000 ;
      RECT  4.795000  16.200000 21.420000  16.270000 ;
      RECT  4.795000  16.200000 21.420000  16.270000 ;
      RECT  4.795000  16.270000 21.490000  16.340000 ;
      RECT  4.795000  16.270000 21.490000  16.340000 ;
      RECT  4.795000  16.340000 21.560000  16.410000 ;
      RECT  4.795000  16.340000 21.560000  16.410000 ;
      RECT  4.795000  16.410000 21.630000  16.480000 ;
      RECT  4.795000  16.410000 21.630000  16.480000 ;
      RECT  4.795000  16.480000 21.700000  16.550000 ;
      RECT  4.795000  16.480000 21.700000  16.550000 ;
      RECT  4.795000  16.550000 21.770000  16.620000 ;
      RECT  4.795000  16.550000 21.770000  16.620000 ;
      RECT  4.795000  16.620000 21.840000  16.690000 ;
      RECT  4.795000  16.620000 21.840000  16.690000 ;
      RECT  4.795000  16.690000 21.910000  16.760000 ;
      RECT  4.795000  16.690000 21.910000  16.760000 ;
      RECT  4.795000  16.760000 21.980000  16.830000 ;
      RECT  4.795000  16.760000 21.980000  16.830000 ;
      RECT  4.795000  16.830000 22.050000  16.900000 ;
      RECT  4.795000  16.830000 22.050000  16.900000 ;
      RECT  4.795000  16.900000 22.120000  16.970000 ;
      RECT  4.795000  16.900000 22.120000  16.970000 ;
      RECT  4.795000  16.970000 22.190000  17.040000 ;
      RECT  4.795000  16.970000 22.190000  17.040000 ;
      RECT  4.795000  17.040000 22.260000  17.110000 ;
      RECT  4.795000  17.040000 22.260000  17.110000 ;
      RECT  4.795000  17.110000 22.330000  17.180000 ;
      RECT  4.795000  17.110000 22.330000  17.180000 ;
      RECT  4.795000  17.180000 22.400000  17.250000 ;
      RECT  4.795000  17.180000 22.400000  17.250000 ;
      RECT  4.795000  17.250000 22.470000  17.320000 ;
      RECT  4.795000  17.250000 22.470000  17.320000 ;
      RECT  4.795000  17.320000 22.540000  17.390000 ;
      RECT  4.795000  17.320000 22.540000  17.390000 ;
      RECT  4.795000  17.390000 22.610000  17.460000 ;
      RECT  4.795000  17.390000 22.610000  17.460000 ;
      RECT  4.795000  17.460000 22.680000  17.530000 ;
      RECT  4.795000  17.460000 22.680000  17.530000 ;
      RECT  4.795000  17.530000 22.750000  17.600000 ;
      RECT  4.795000  17.530000 22.750000  17.600000 ;
      RECT  4.795000  17.600000 22.820000  17.670000 ;
      RECT  4.795000  17.600000 22.820000  17.670000 ;
      RECT  4.795000  17.670000 22.890000  17.740000 ;
      RECT  4.795000  17.670000 22.890000  17.740000 ;
      RECT  4.795000  17.740000 22.960000  17.810000 ;
      RECT  4.795000  17.740000 22.960000  17.810000 ;
      RECT  4.795000  17.810000 23.030000  17.880000 ;
      RECT  4.795000  17.810000 23.030000  17.880000 ;
      RECT  4.795000  17.880000 23.100000  17.950000 ;
      RECT  4.795000  17.880000 23.100000  17.950000 ;
      RECT  4.795000  17.950000 23.170000  18.020000 ;
      RECT  4.795000  17.950000 23.170000  18.020000 ;
      RECT  4.795000  18.020000 23.240000  18.090000 ;
      RECT  4.795000  18.020000 23.240000  18.090000 ;
      RECT  4.795000  18.090000 23.310000  18.160000 ;
      RECT  4.795000  18.090000 23.310000  18.160000 ;
      RECT  4.795000  18.160000 23.380000  18.230000 ;
      RECT  4.795000  18.160000 23.380000  18.230000 ;
      RECT  4.795000  18.230000 23.450000  18.300000 ;
      RECT  4.795000  18.230000 23.450000  18.300000 ;
      RECT  4.795000  18.300000 23.520000  18.370000 ;
      RECT  4.795000  18.300000 23.520000  18.370000 ;
      RECT  4.795000  18.370000 23.590000  18.440000 ;
      RECT  4.795000  18.370000 23.590000  18.440000 ;
      RECT  4.795000  18.440000 23.660000  18.510000 ;
      RECT  4.795000  18.440000 23.660000  18.510000 ;
      RECT  4.795000  18.510000 23.730000  18.580000 ;
      RECT  4.795000  18.510000 23.730000  18.580000 ;
      RECT  4.795000  18.580000 23.800000  18.650000 ;
      RECT  4.795000  18.580000 23.800000  18.650000 ;
      RECT  4.795000  18.650000 23.870000  18.720000 ;
      RECT  4.795000  18.650000 23.870000  18.720000 ;
      RECT  4.795000  18.720000 23.940000  18.725000 ;
      RECT  4.795000  18.720000 23.940000  18.725000 ;
      RECT  4.795000  18.725000 23.945000  25.470000 ;
      RECT  4.795000  18.725000 23.945000  26.060000 ;
      RECT  4.795000  25.470000 23.945000  25.540000 ;
      RECT  4.795000  25.470000 23.945000  25.540000 ;
      RECT  4.795000  25.540000 24.015000  25.610000 ;
      RECT  4.795000  25.540000 24.015000  25.610000 ;
      RECT  4.795000  25.610000 24.085000  25.680000 ;
      RECT  4.795000  25.610000 24.085000  25.680000 ;
      RECT  4.795000  25.680000 24.155000  25.750000 ;
      RECT  4.795000  25.680000 24.155000  25.750000 ;
      RECT  4.795000  25.750000 24.225000  25.820000 ;
      RECT  4.795000  25.750000 24.225000  25.820000 ;
      RECT  4.795000  25.820000 24.295000  25.890000 ;
      RECT  4.795000  25.820000 24.295000  25.890000 ;
      RECT  4.795000  25.890000 24.365000  25.960000 ;
      RECT  4.795000  25.890000 24.365000  25.960000 ;
      RECT  4.795000  25.960000 24.435000  26.030000 ;
      RECT  4.795000  25.960000 24.435000  26.030000 ;
      RECT  4.795000  26.030000 24.505000  26.060000 ;
      RECT  4.795000  26.030000 24.505000  26.060000 ;
      RECT  4.795000  26.060000 24.535000  42.625000 ;
      RECT  4.795000  42.625000 24.465000  42.695000 ;
      RECT  4.795000  42.625000 24.465000  42.695000 ;
      RECT  4.795000  42.695000 24.395000  42.765000 ;
      RECT  4.795000  42.695000 24.395000  42.765000 ;
      RECT  4.795000  42.765000 24.325000  42.835000 ;
      RECT  4.795000  42.765000 24.325000  42.835000 ;
      RECT  4.795000  42.835000 24.255000  42.905000 ;
      RECT  4.795000  42.835000 24.255000  42.905000 ;
      RECT  4.795000  42.905000 24.185000  42.975000 ;
      RECT  4.795000  42.905000 24.185000  42.975000 ;
      RECT  4.795000  42.975000 24.155000  43.005000 ;
      RECT  4.795000  42.975000 24.155000  43.005000 ;
      RECT  4.795000  43.005000  5.785000  43.825000 ;
      RECT  4.795000  43.825000 73.380000  71.630000 ;
      RECT  5.990000   0.870000 12.005000   3.430000 ;
      RECT  6.225000 143.875000 70.525000 144.285000 ;
      RECT  6.225000 144.285000 70.455000 144.355000 ;
      RECT  6.225000 144.285000 70.455000 144.355000 ;
      RECT  6.225000 144.355000 70.385000 144.425000 ;
      RECT  6.225000 144.355000 70.385000 144.425000 ;
      RECT  6.225000 144.425000 70.315000 144.495000 ;
      RECT  6.225000 144.425000 70.315000 144.495000 ;
      RECT  6.225000 144.495000 70.245000 144.565000 ;
      RECT  6.225000 144.495000 70.245000 144.565000 ;
      RECT  6.225000 144.565000 70.175000 144.635000 ;
      RECT  6.225000 144.565000 70.175000 144.635000 ;
      RECT  6.225000 144.635000 70.105000 144.705000 ;
      RECT  6.225000 144.635000 70.105000 144.705000 ;
      RECT  6.225000 144.705000 70.035000 144.775000 ;
      RECT  6.225000 144.705000 70.035000 144.775000 ;
      RECT  6.225000 144.775000 69.965000 144.845000 ;
      RECT  6.225000 144.775000 69.965000 144.845000 ;
      RECT  6.225000 144.845000 69.960000 144.850000 ;
      RECT  6.225000 144.845000 69.960000 144.850000 ;
      RECT  6.225000 144.850000 69.890000 144.920000 ;
      RECT  6.225000 144.850000 69.890000 144.920000 ;
      RECT  6.225000 144.920000 69.820000 144.990000 ;
      RECT  6.225000 144.920000 69.820000 144.990000 ;
      RECT  6.225000 144.990000 69.750000 145.060000 ;
      RECT  6.225000 144.990000 69.750000 145.060000 ;
      RECT  6.225000 145.060000 69.680000 145.130000 ;
      RECT  6.225000 145.060000 69.680000 145.130000 ;
      RECT  6.225000 145.130000 69.610000 145.200000 ;
      RECT  6.225000 145.130000 69.610000 145.200000 ;
      RECT  6.225000 145.200000 69.540000 145.270000 ;
      RECT  6.225000 145.200000 69.540000 145.270000 ;
      RECT  6.225000 145.270000 69.470000 145.340000 ;
      RECT  6.225000 145.270000 69.470000 145.340000 ;
      RECT  6.225000 145.340000 69.400000 145.410000 ;
      RECT  6.225000 145.340000 69.400000 145.410000 ;
      RECT  6.225000 145.410000 70.525000 146.420000 ;
      RECT  6.225000 145.410000 70.525000 195.970000 ;
      RECT  8.190000 132.395000 72.380000 132.460000 ;
      RECT  8.190000 132.395000 72.380000 132.460000 ;
      RECT  8.260000 132.325000 72.380000 132.395000 ;
      RECT  8.260000 132.325000 72.380000 132.395000 ;
      RECT  8.330000 132.255000 72.380000 132.325000 ;
      RECT  8.330000 132.255000 72.380000 132.325000 ;
      RECT  8.400000 132.185000 72.380000 132.255000 ;
      RECT  8.400000 132.185000 72.380000 132.255000 ;
      RECT  8.470000 132.115000 72.380000 132.185000 ;
      RECT  8.470000 132.115000 72.380000 132.185000 ;
      RECT  8.540000 132.045000 72.380000 132.115000 ;
      RECT  8.540000 132.045000 72.380000 132.115000 ;
      RECT  8.610000 131.975000 72.380000 132.045000 ;
      RECT  8.610000 131.975000 72.380000 132.045000 ;
      RECT  8.680000 131.905000 72.380000 131.975000 ;
      RECT  8.680000 131.905000 72.380000 131.975000 ;
      RECT  8.750000 131.835000 72.380000 131.905000 ;
      RECT  8.750000 131.835000 72.380000 131.905000 ;
      RECT  8.820000 131.765000 72.380000 131.835000 ;
      RECT  8.820000 131.765000 72.380000 131.835000 ;
      RECT  8.890000 131.695000 72.380000 131.765000 ;
      RECT  8.890000 131.695000 72.380000 131.765000 ;
      RECT  8.960000 131.625000 72.380000 131.695000 ;
      RECT  8.960000 131.625000 72.380000 131.695000 ;
      RECT  9.030000 131.555000 72.380000 131.625000 ;
      RECT  9.030000 131.555000 72.380000 131.625000 ;
      RECT  9.100000 131.485000 72.380000 131.555000 ;
      RECT  9.100000 131.485000 72.380000 131.555000 ;
      RECT  9.170000 131.415000 72.380000 131.485000 ;
      RECT  9.170000 131.415000 72.380000 131.485000 ;
      RECT  9.240000 131.345000 72.380000 131.415000 ;
      RECT  9.240000 131.345000 72.380000 131.415000 ;
      RECT  9.310000 131.275000 72.380000 131.345000 ;
      RECT  9.310000 131.275000 72.380000 131.345000 ;
      RECT  9.380000 131.205000 72.380000 131.275000 ;
      RECT  9.380000 131.205000 72.380000 131.275000 ;
      RECT  9.450000 131.135000 72.380000 131.205000 ;
      RECT  9.450000 131.135000 72.380000 131.205000 ;
      RECT  9.520000 131.065000 72.380000 131.135000 ;
      RECT  9.520000 131.065000 72.380000 131.135000 ;
      RECT  9.590000 130.995000 72.380000 131.065000 ;
      RECT  9.590000 130.995000 72.380000 131.065000 ;
      RECT  9.595000 130.990000 72.380000 130.995000 ;
      RECT  9.595000 130.990000 72.380000 130.995000 ;
      RECT  9.665000 130.920000 72.380000 130.990000 ;
      RECT  9.665000 130.920000 72.380000 130.990000 ;
      RECT  9.735000 130.850000 72.380000 130.920000 ;
      RECT  9.735000 130.850000 72.380000 130.920000 ;
      RECT  9.805000 130.780000 72.380000 130.850000 ;
      RECT  9.805000 130.780000 72.380000 130.850000 ;
      RECT  9.875000 130.710000 72.380000 130.780000 ;
      RECT  9.875000 130.710000 72.380000 130.780000 ;
      RECT  9.945000 130.640000 72.380000 130.710000 ;
      RECT  9.945000 130.640000 72.380000 130.710000 ;
      RECT 10.015000 130.570000 72.380000 130.640000 ;
      RECT 10.015000 130.570000 72.380000 130.640000 ;
      RECT 10.085000 130.500000 72.380000 130.570000 ;
      RECT 10.085000 130.500000 72.380000 130.570000 ;
      RECT 10.155000 130.430000 64.845000 130.500000 ;
      RECT 10.155000 130.430000 64.845000 130.500000 ;
      RECT 10.225000 130.360000 64.775000 130.430000 ;
      RECT 10.225000 130.360000 64.775000 130.430000 ;
      RECT 10.295000 130.290000 64.705000 130.360000 ;
      RECT 10.295000 130.290000 64.705000 130.360000 ;
      RECT 10.365000 130.220000 64.635000 130.290000 ;
      RECT 10.365000 130.220000 64.635000 130.290000 ;
      RECT 10.435000 130.150000 64.565000 130.220000 ;
      RECT 10.435000 130.150000 64.565000 130.220000 ;
      RECT 10.505000 130.080000 64.495000 130.150000 ;
      RECT 10.505000 130.080000 64.495000 130.150000 ;
      RECT 10.575000 130.010000 64.425000 130.080000 ;
      RECT 10.575000 130.010000 64.425000 130.080000 ;
      RECT 10.645000 129.940000 64.355000 130.010000 ;
      RECT 10.645000 129.940000 64.355000 130.010000 ;
      RECT 10.715000 129.870000 64.285000 129.940000 ;
      RECT 10.715000 129.870000 64.285000 129.940000 ;
      RECT 10.785000 129.800000 64.215000 129.870000 ;
      RECT 10.785000 129.800000 64.215000 129.870000 ;
      RECT 10.855000 129.730000 64.145000 129.800000 ;
      RECT 10.855000 129.730000 64.145000 129.800000 ;
      RECT 10.925000 129.660000 64.075000 129.730000 ;
      RECT 10.925000 129.660000 64.075000 129.730000 ;
      RECT 10.995000 129.590000 64.005000 129.660000 ;
      RECT 10.995000 129.590000 64.005000 129.660000 ;
      RECT 11.065000 129.520000 63.935000 129.590000 ;
      RECT 11.065000 129.520000 63.935000 129.590000 ;
      RECT 11.135000 129.450000 63.865000 129.520000 ;
      RECT 11.135000 129.450000 63.865000 129.520000 ;
      RECT 11.205000 129.380000 63.795000 129.450000 ;
      RECT 11.205000 129.380000 63.795000 129.450000 ;
      RECT 11.255000 139.225000 14.920000 139.260000 ;
      RECT 11.255000 139.225000 14.920000 139.260000 ;
      RECT 11.275000 129.310000 63.725000 129.380000 ;
      RECT 11.275000 129.310000 63.725000 129.380000 ;
      RECT 11.290000 139.260000 14.920000 139.295000 ;
      RECT 11.290000 139.260000 14.920000 139.295000 ;
      RECT 11.345000 129.240000 63.655000 129.310000 ;
      RECT 11.345000 129.240000 63.655000 129.310000 ;
      RECT 11.415000 129.170000 63.585000 129.240000 ;
      RECT 11.415000 129.170000 63.585000 129.240000 ;
      RECT 11.485000 129.100000 63.515000 129.170000 ;
      RECT 11.485000 129.100000 63.515000 129.170000 ;
      RECT 11.555000 129.030000 63.445000 129.100000 ;
      RECT 11.555000 129.030000 63.445000 129.100000 ;
      RECT 11.625000 128.960000 63.375000 129.030000 ;
      RECT 11.625000 128.960000 63.375000 129.030000 ;
      RECT 11.695000 128.890000 63.305000 128.960000 ;
      RECT 11.695000 128.890000 63.305000 128.960000 ;
      RECT 11.765000 128.820000 63.235000 128.890000 ;
      RECT 11.765000 128.820000 63.235000 128.890000 ;
      RECT 11.835000 128.750000 63.165000 128.820000 ;
      RECT 11.835000 128.750000 63.165000 128.820000 ;
      RECT 11.905000 128.680000 63.095000 128.750000 ;
      RECT 11.905000 128.680000 63.095000 128.750000 ;
      RECT 11.950000 128.240000 63.050000 128.260000 ;
      RECT 11.975000 128.610000 63.025000 128.680000 ;
      RECT 11.975000 128.610000 63.025000 128.680000 ;
      RECT 12.020000 128.170000 62.980000 128.240000 ;
      RECT 12.045000 128.540000 62.955000 128.610000 ;
      RECT 12.045000 128.540000 62.955000 128.610000 ;
      RECT 12.090000 128.100000 62.910000 128.170000 ;
      RECT 12.160000 128.030000 62.840000 128.100000 ;
      RECT 12.230000 127.960000 62.770000 128.030000 ;
      RECT 12.300000 127.890000 62.700000 127.960000 ;
      RECT 12.370000 127.820000 62.630000 127.890000 ;
      RECT 12.440000 127.750000 62.560000 127.820000 ;
      RECT 12.510000 127.680000 62.490000 127.750000 ;
      RECT 12.580000 127.610000 62.420000 127.680000 ;
      RECT 12.650000 127.540000 62.350000 127.610000 ;
      RECT 12.685000   0.000000 14.415000   6.715000 ;
      RECT 12.685000   6.715000 14.415000   7.070000 ;
      RECT 12.720000 127.470000 62.280000 127.540000 ;
      RECT 12.790000 127.400000 62.210000 127.470000 ;
      RECT 12.825000   3.550000 14.275000   6.660000 ;
      RECT 12.860000 127.330000 62.140000 127.400000 ;
      RECT 12.895000   6.660000 14.275000   6.730000 ;
      RECT 12.920000   0.240000 13.915000   3.270000 ;
      RECT 12.930000 127.260000 62.070000 127.330000 ;
      RECT 12.965000   6.730000 14.275000   6.800000 ;
      RECT 12.970000  10.555000 14.275000  10.585000 ;
      RECT 13.000000 127.190000 62.000000 127.260000 ;
      RECT 13.035000   6.800000 14.275000   6.870000 ;
      RECT 13.040000   7.070000 14.415000  10.290000 ;
      RECT 13.040000  10.290000 14.415000  10.445000 ;
      RECT 13.040000  10.485000 14.275000  10.555000 ;
      RECT 13.070000 127.120000 61.930000 127.190000 ;
      RECT 13.105000   6.870000 14.275000   6.940000 ;
      RECT 13.110000  10.415000 14.275000  10.485000 ;
      RECT 13.140000 127.050000 61.860000 127.120000 ;
      RECT 13.175000   6.940000 14.275000   7.010000 ;
      RECT 13.180000   7.010000 14.275000   7.015000 ;
      RECT 13.180000   7.015000 14.275000  10.345000 ;
      RECT 13.180000  10.345000 14.275000  10.415000 ;
      RECT 13.210000 126.980000 61.790000 127.050000 ;
      RECT 13.280000 126.910000 61.720000 126.980000 ;
      RECT 13.350000 126.840000 61.650000 126.910000 ;
      RECT 13.390000 130.500000 72.380000 135.750000 ;
      RECT 13.390000 132.460000 72.380000 135.285000 ;
      RECT 13.390000 135.285000 72.310000 135.355000 ;
      RECT 13.390000 135.285000 72.310000 135.355000 ;
      RECT 13.390000 135.355000 72.240000 135.425000 ;
      RECT 13.390000 135.355000 72.240000 135.425000 ;
      RECT 13.390000 135.425000 72.170000 135.495000 ;
      RECT 13.390000 135.425000 72.170000 135.495000 ;
      RECT 13.390000 135.495000 72.100000 135.565000 ;
      RECT 13.390000 135.495000 72.100000 135.565000 ;
      RECT 13.390000 135.565000 72.030000 135.635000 ;
      RECT 13.390000 135.565000 72.030000 135.635000 ;
      RECT 13.390000 135.635000 71.960000 135.705000 ;
      RECT 13.390000 135.635000 71.960000 135.705000 ;
      RECT 13.390000 135.705000 71.915000 135.750000 ;
      RECT 13.390000 135.705000 71.915000 135.750000 ;
      RECT 13.420000 126.770000 61.580000 126.840000 ;
      RECT 13.490000 126.700000 61.510000 126.770000 ;
      RECT 13.560000 126.630000 61.440000 126.700000 ;
      RECT 13.630000 126.560000 61.370000 126.630000 ;
      RECT 13.700000 126.490000 61.300000 126.560000 ;
      RECT 13.770000 126.420000 61.230000 126.490000 ;
      RECT 13.840000 126.350000 61.160000 126.420000 ;
      RECT 13.910000 126.280000 61.090000 126.350000 ;
      RECT 13.980000 126.210000 61.020000 126.280000 ;
      RECT 14.050000 126.140000 60.950000 126.210000 ;
      RECT 14.120000 126.070000 60.880000 126.140000 ;
      RECT 14.190000 126.000000 60.810000 126.070000 ;
      RECT 14.260000 125.930000 60.740000 126.000000 ;
      RECT 14.330000 125.860000 60.670000 125.930000 ;
      RECT 14.400000 125.790000 60.600000 125.860000 ;
      RECT 14.470000 125.720000 60.530000 125.790000 ;
      RECT 14.540000 125.650000 60.460000 125.720000 ;
      RECT 14.610000 125.580000 60.390000 125.650000 ;
      RECT 14.680000 125.510000 60.320000 125.580000 ;
      RECT 14.750000 125.440000 60.250000 125.510000 ;
      RECT 15.200000 138.990000 69.130000 139.060000 ;
      RECT 15.200000 139.060000 69.200000 139.130000 ;
      RECT 15.200000 139.130000 69.270000 139.200000 ;
      RECT 15.200000 139.200000 69.340000 139.270000 ;
      RECT 15.200000 139.270000 69.410000 139.340000 ;
      RECT 15.200000 139.340000 69.480000 139.410000 ;
      RECT 15.200000 139.410000 69.550000 139.480000 ;
      RECT 15.200000 139.480000 69.620000 139.550000 ;
      RECT 15.200000 139.550000 69.690000 139.575000 ;
      RECT 15.275000   0.000000 22.220000   1.345000 ;
      RECT 15.275000   1.345000 24.765000  11.280000 ;
      RECT 15.275000  11.280000 16.460000  12.150000 ;
      RECT 15.275000  12.150000 16.460000  12.470000 ;
      RECT 15.415000   0.830000 16.780000   3.430000 ;
      RECT 15.415000   3.430000 24.625000  11.140000 ;
      RECT 15.415000  11.140000 16.320000  12.095000 ;
      RECT 15.485000  12.095000 16.320000  12.165000 ;
      RECT 15.525000   0.200000 21.315000   0.550000 ;
      RECT 15.555000  12.165000 16.320000  12.235000 ;
      RECT 15.590000  12.470000 16.995000  13.005000 ;
      RECT 15.625000  12.235000 16.320000  12.305000 ;
      RECT 15.695000  12.305000 16.320000  12.375000 ;
      RECT 15.765000  12.375000 16.320000  12.445000 ;
      RECT 15.835000  12.445000 16.320000  12.515000 ;
      RECT 15.845000  12.515000 16.320000  12.525000 ;
      RECT 15.915000  12.525000 16.320000  12.595000 ;
      RECT 15.985000  12.595000 16.390000  12.665000 ;
      RECT 16.055000  12.665000 16.460000  12.735000 ;
      RECT 16.125000  12.735000 16.530000  12.805000 ;
      RECT 16.125000  13.005000 25.015000  13.175000 ;
      RECT 16.195000  12.805000 16.600000  12.875000 ;
      RECT 16.265000  12.875000 16.670000  12.945000 ;
      RECT 16.295000  13.175000 25.015000  15.195000 ;
      RECT 16.335000  12.945000 16.740000  13.015000 ;
      RECT 16.405000  13.015000 16.810000  13.085000 ;
      RECT 16.465000  13.085000 16.880000  13.145000 ;
      RECT 16.510000  13.145000 24.790000  13.190000 ;
      RECT 16.550000  13.190000 24.835000  13.230000 ;
      RECT 16.620000  13.230000 24.875000  13.300000 ;
      RECT 16.690000  13.300000 24.875000  13.370000 ;
      RECT 16.760000  13.370000 24.875000  13.440000 ;
      RECT 16.830000  13.440000 24.875000  13.510000 ;
      RECT 16.885000 138.985000 75.145000 138.990000 ;
      RECT 16.900000  13.510000 24.875000  13.580000 ;
      RECT 16.905000 138.965000 75.145000 138.985000 ;
      RECT 16.925000 138.945000 75.145000 138.965000 ;
      RECT 16.970000  11.280000 24.765000  12.250000 ;
      RECT 16.970000  12.250000 24.765000  12.290000 ;
      RECT 16.970000  13.580000 24.875000  13.650000 ;
      RECT 17.010000  12.290000 24.560000  12.495000 ;
      RECT 17.040000  13.650000 24.875000  13.720000 ;
      RECT 17.060000   1.140000 18.910000   3.150000 ;
      RECT 17.110000   3.430000 24.625000  12.195000 ;
      RECT 17.110000  11.140000 24.625000  12.195000 ;
      RECT 17.110000  13.720000 24.875000  13.790000 ;
      RECT 17.130000  12.195000 24.625000  12.215000 ;
      RECT 17.130000  12.195000 24.625000  12.215000 ;
      RECT 17.150000  12.215000 24.625000  12.235000 ;
      RECT 17.150000  12.215000 24.625000  12.235000 ;
      RECT 17.180000  13.790000 24.875000  13.860000 ;
      RECT 17.210000  12.235000 24.565000  12.295000 ;
      RECT 17.210000  12.235000 24.565000  12.295000 ;
      RECT 17.250000  13.860000 24.875000  13.930000 ;
      RECT 17.270000  12.295000 24.505000  12.355000 ;
      RECT 17.270000  12.295000 24.505000  12.355000 ;
      RECT 17.320000  13.930000 24.875000  14.000000 ;
      RECT 17.390000  14.000000 24.875000  14.070000 ;
      RECT 17.460000  14.070000 24.875000  14.140000 ;
      RECT 17.530000  14.140000 24.875000  14.210000 ;
      RECT 17.600000  14.210000 24.875000  14.280000 ;
      RECT 17.670000  14.280000 24.875000  14.350000 ;
      RECT 17.740000  14.350000 24.875000  14.420000 ;
      RECT 17.810000  14.420000 24.875000  14.490000 ;
      RECT 17.880000  14.490000 24.875000  14.560000 ;
      RECT 17.950000  14.560000 24.875000  14.630000 ;
      RECT 18.020000  14.630000 24.875000  14.700000 ;
      RECT 18.090000  14.700000 24.875000  14.770000 ;
      RECT 18.160000  14.770000 24.875000  14.840000 ;
      RECT 18.230000  14.840000 24.875000  14.910000 ;
      RECT 18.300000  14.910000 24.875000  14.980000 ;
      RECT 18.315000  15.195000 25.100000  15.280000 ;
      RECT 18.370000  14.980000 24.875000  15.050000 ;
      RECT 18.440000  15.050000 24.875000  15.120000 ;
      RECT 18.460000  15.120000 24.875000  15.140000 ;
      RECT 18.985000   0.550000 21.315000   0.620000 ;
      RECT 19.055000   0.620000 21.315000   0.690000 ;
      RECT 19.125000   0.690000 21.315000   0.760000 ;
      RECT 19.190000   2.785000 22.900000   2.855000 ;
      RECT 19.190000   2.785000 22.900000   2.855000 ;
      RECT 19.190000   2.855000 22.970000   2.925000 ;
      RECT 19.190000   2.855000 22.970000   2.925000 ;
      RECT 19.190000   2.925000 23.040000   2.995000 ;
      RECT 19.190000   2.925000 23.040000   2.995000 ;
      RECT 19.190000   2.995000 23.110000   3.065000 ;
      RECT 19.190000   2.995000 23.110000   3.065000 ;
      RECT 19.190000   3.065000 23.180000   3.135000 ;
      RECT 19.190000   3.065000 23.180000   3.135000 ;
      RECT 19.190000   3.135000 23.250000   3.205000 ;
      RECT 19.190000   3.135000 23.250000   3.205000 ;
      RECT 19.190000   3.205000 23.320000   3.275000 ;
      RECT 19.190000   3.205000 23.320000   3.275000 ;
      RECT 19.190000   3.275000 23.390000   3.280000 ;
      RECT 19.190000   3.275000 23.390000   3.280000 ;
      RECT 19.190000   3.280000 24.625000   3.430000 ;
      RECT 19.190000   3.280000 24.625000  11.140000 ;
      RECT 19.190000   3.280000 24.625000  11.140000 ;
      RECT 19.195000   0.760000 21.315000   0.830000 ;
      RECT 19.265000   0.830000 21.385000   0.900000 ;
      RECT 19.335000   0.900000 21.455000   0.970000 ;
      RECT 19.405000   0.970000 21.525000   1.040000 ;
      RECT 19.475000   1.040000 21.595000   1.110000 ;
      RECT 19.540000  71.630000 73.380000  80.155000 ;
      RECT 19.545000   1.110000 21.665000   1.180000 ;
      RECT 19.580000   1.180000 21.735000   1.215000 ;
      RECT 19.580000   1.215000 21.770000   1.285000 ;
      RECT 19.580000   1.285000 21.840000   1.355000 ;
      RECT 19.580000   1.355000 21.910000   1.425000 ;
      RECT 19.580000   1.425000 21.980000   1.495000 ;
      RECT 19.580000   1.495000 22.050000   1.565000 ;
      RECT 19.580000   1.565000 22.120000   1.585000 ;
      RECT 19.580000   1.585000 24.585000   2.505000 ;
      RECT 21.595000   0.000000 22.080000   0.645000 ;
      RECT 21.665000   0.645000 22.080000   0.715000 ;
      RECT 21.735000   0.715000 22.080000   0.785000 ;
      RECT 21.805000   0.785000 22.080000   0.855000 ;
      RECT 21.805000  15.280000 25.805000  15.985000 ;
      RECT 21.875000   0.855000 22.080000   0.925000 ;
      RECT 21.915000  15.140000 24.875000  15.195000 ;
      RECT 21.945000   0.925000 22.080000   0.995000 ;
      RECT 21.970000  15.195000 24.875000  15.250000 ;
      RECT 22.015000   0.995000 22.080000   1.065000 ;
      RECT 22.040000  15.250000 24.875000  15.320000 ;
      RECT 22.110000  15.320000 24.945000  15.390000 ;
      RECT 22.180000  15.390000 25.015000  15.460000 ;
      RECT 22.250000  15.460000 25.085000  15.530000 ;
      RECT 22.320000  15.530000 25.155000  15.600000 ;
      RECT 22.390000  15.600000 25.225000  15.670000 ;
      RECT 22.460000  15.670000 25.295000  15.740000 ;
      RECT 22.505000  15.985000 30.665000  16.845000 ;
      RECT 22.530000  15.740000 25.365000  15.810000 ;
      RECT 22.600000  15.810000 25.435000  15.880000 ;
      RECT 22.670000  15.880000 25.505000  15.950000 ;
      RECT 22.740000  15.950000 25.575000  16.020000 ;
      RECT 22.790000   1.560000 24.585000   1.585000 ;
      RECT 22.800000   0.000000 24.765000   1.345000 ;
      RECT 22.810000  16.020000 25.645000  16.090000 ;
      RECT 22.845000  16.090000 25.715000  16.125000 ;
      RECT 22.860000   1.490000 24.585000   1.560000 ;
      RECT 22.915000  16.125000 29.750000  16.195000 ;
      RECT 22.915000  16.125000 29.750000  16.195000 ;
      RECT 22.930000   1.420000 24.585000   1.490000 ;
      RECT 22.940000   0.000000 24.625000   0.390000 ;
      RECT 22.940000   0.390000 23.210000   0.745000 ;
      RECT 22.940000   0.745000 23.140000   0.815000 ;
      RECT 22.940000   0.815000 23.070000   0.885000 ;
      RECT 22.940000   0.885000 23.000000   0.955000 ;
      RECT 22.985000  16.195000 29.820000  16.265000 ;
      RECT 22.985000  16.195000 29.820000  16.265000 ;
      RECT 23.000000   1.350000 24.585000   1.420000 ;
      RECT 23.055000  16.265000 29.890000  16.335000 ;
      RECT 23.055000  16.265000 29.890000  16.335000 ;
      RECT 23.070000   1.280000 24.585000   1.350000 ;
      RECT 23.085000   2.505000 24.585000   2.575000 ;
      RECT 23.125000  16.335000 29.960000  16.405000 ;
      RECT 23.125000  16.335000 29.960000  16.405000 ;
      RECT 23.140000   1.210000 24.585000   1.280000 ;
      RECT 23.155000   2.575000 24.585000   2.645000 ;
      RECT 23.195000  16.405000 30.030000  16.475000 ;
      RECT 23.195000  16.405000 30.030000  16.475000 ;
      RECT 23.210000   1.140000 24.585000   1.210000 ;
      RECT 23.225000   2.645000 24.585000   2.715000 ;
      RECT 23.265000  16.475000 30.100000  16.545000 ;
      RECT 23.265000  16.475000 30.100000  16.545000 ;
      RECT 23.280000   1.070000 24.585000   1.140000 ;
      RECT 23.295000   2.715000 24.585000   2.785000 ;
      RECT 23.335000  16.545000 30.170000  16.615000 ;
      RECT 23.335000  16.545000 30.170000  16.615000 ;
      RECT 23.350000   1.000000 24.585000   1.070000 ;
      RECT 23.365000   2.785000 24.585000   2.855000 ;
      RECT 23.365000  16.845000 30.665000  18.340000 ;
      RECT 23.405000  16.615000 30.240000  16.685000 ;
      RECT 23.405000  16.615000 30.240000  16.685000 ;
      RECT 23.420000   0.930000 24.585000   1.000000 ;
      RECT 23.435000   2.855000 24.585000   2.925000 ;
      RECT 23.475000  16.685000 30.310000  16.755000 ;
      RECT 23.475000  16.685000 30.310000  16.755000 ;
      RECT 23.490000   0.670000 24.585000   0.860000 ;
      RECT 23.490000   0.860000 24.585000   0.930000 ;
      RECT 23.505000   2.925000 24.585000   2.995000 ;
      RECT 23.510000   2.995000 24.585000   3.000000 ;
      RECT 23.545000  16.755000 30.380000  16.825000 ;
      RECT 23.545000  16.755000 30.380000  16.825000 ;
      RECT 23.615000  16.825000 30.450000  16.895000 ;
      RECT 23.615000  16.825000 30.450000  16.895000 ;
      RECT 23.620000  16.895000 30.520000  16.900000 ;
      RECT 23.620000  16.895000 30.520000  16.900000 ;
      RECT 23.690000  16.900000 30.525000  16.970000 ;
      RECT 23.690000  16.900000 30.525000  16.970000 ;
      RECT 23.760000  16.970000 30.525000  17.040000 ;
      RECT 23.760000  16.970000 30.525000  17.040000 ;
      RECT 23.830000  17.040000 30.525000  17.110000 ;
      RECT 23.830000  17.040000 30.525000  17.110000 ;
      RECT 23.900000  17.110000 30.525000  17.180000 ;
      RECT 23.900000  17.110000 30.525000  17.180000 ;
      RECT 23.970000  17.180000 30.525000  17.250000 ;
      RECT 23.970000  17.180000 30.525000  17.250000 ;
      RECT 24.040000  17.250000 30.525000  17.320000 ;
      RECT 24.040000  17.250000 30.525000  17.320000 ;
      RECT 24.110000  17.320000 30.525000  17.390000 ;
      RECT 24.110000  17.320000 30.525000  17.390000 ;
      RECT 24.180000  17.390000 30.525000  17.460000 ;
      RECT 24.180000  17.390000 30.525000  17.460000 ;
      RECT 24.250000  17.460000 30.525000  17.530000 ;
      RECT 24.250000  17.460000 30.525000  17.530000 ;
      RECT 24.320000  17.530000 30.525000  17.600000 ;
      RECT 24.320000  17.530000 30.525000  17.600000 ;
      RECT 24.390000  17.600000 30.525000  17.670000 ;
      RECT 24.390000  17.600000 30.525000  17.670000 ;
      RECT 24.460000  17.670000 30.525000  17.740000 ;
      RECT 24.460000  17.670000 30.525000  17.740000 ;
      RECT 24.530000  17.740000 30.525000  17.810000 ;
      RECT 24.530000  17.740000 30.525000  17.810000 ;
      RECT 24.545000  43.775000 73.380000  43.825000 ;
      RECT 24.545000  43.775000 73.380000  43.825000 ;
      RECT 24.600000  17.810000 30.525000  17.880000 ;
      RECT 24.600000  17.810000 30.525000  17.880000 ;
      RECT 24.615000  43.705000 73.380000  43.775000 ;
      RECT 24.615000  43.705000 73.380000  43.775000 ;
      RECT 24.670000  17.880000 30.525000  17.950000 ;
      RECT 24.670000  17.880000 30.525000  17.950000 ;
      RECT 24.685000  43.635000 73.380000  43.705000 ;
      RECT 24.685000  43.635000 73.380000  43.705000 ;
      RECT 24.740000  17.950000 30.525000  18.020000 ;
      RECT 24.740000  17.950000 30.525000  18.020000 ;
      RECT 24.755000  43.565000 73.380000  43.635000 ;
      RECT 24.755000  43.565000 73.380000  43.635000 ;
      RECT 24.810000  18.020000 30.525000  18.090000 ;
      RECT 24.810000  18.020000 30.525000  18.090000 ;
      RECT 24.825000  43.495000 73.380000  43.565000 ;
      RECT 24.825000  43.495000 73.380000  43.565000 ;
      RECT 24.865000  18.340000 30.665000  19.485000 ;
      RECT 24.865000  19.485000 32.625000  25.085000 ;
      RECT 24.865000  25.085000 32.625000  25.675000 ;
      RECT 24.880000  18.090000 30.525000  18.160000 ;
      RECT 24.880000  18.090000 30.525000  18.160000 ;
      RECT 24.895000  43.425000 73.380000  43.495000 ;
      RECT 24.895000  43.425000 73.380000  43.495000 ;
      RECT 24.950000  18.160000 30.525000  18.230000 ;
      RECT 24.950000  18.160000 30.525000  18.230000 ;
      RECT 24.965000  43.355000 73.380000  43.425000 ;
      RECT 24.965000  43.355000 73.380000  43.425000 ;
      RECT 25.005000  16.900000 30.525000  25.030000 ;
      RECT 25.005000  18.230000 30.525000  18.285000 ;
      RECT 25.005000  18.230000 30.525000  18.285000 ;
      RECT 25.005000  18.285000 30.525000  19.625000 ;
      RECT 25.005000  19.625000 32.485000  25.030000 ;
      RECT 25.035000  43.285000 73.380000  43.355000 ;
      RECT 25.035000  43.285000 73.380000  43.355000 ;
      RECT 25.075000  25.030000 32.485000  25.100000 ;
      RECT 25.075000  25.030000 32.485000  25.100000 ;
      RECT 25.105000  43.215000 73.380000  43.285000 ;
      RECT 25.105000  43.215000 73.380000  43.285000 ;
      RECT 25.145000  25.100000 32.485000  25.170000 ;
      RECT 25.145000  25.100000 32.485000  25.170000 ;
      RECT 25.175000  43.145000 73.380000  43.215000 ;
      RECT 25.175000  43.145000 73.380000  43.215000 ;
      RECT 25.215000  25.170000 32.485000  25.240000 ;
      RECT 25.215000  25.170000 32.485000  25.240000 ;
      RECT 25.245000  43.075000 73.380000  43.145000 ;
      RECT 25.245000  43.075000 73.380000  43.145000 ;
      RECT 25.275000   0.000000 27.440000   3.180000 ;
      RECT 25.275000   3.180000 28.045000   3.785000 ;
      RECT 25.275000   3.785000 28.045000   4.245000 ;
      RECT 25.275000   4.245000 29.310000   4.755000 ;
      RECT 25.275000   4.755000 28.045000   5.685000 ;
      RECT 25.275000   5.685000 32.620000   8.890000 ;
      RECT 25.275000   8.890000 32.625000   8.895000 ;
      RECT 25.275000   8.895000 32.625000  12.415000 ;
      RECT 25.275000  12.415000 32.625000  12.665000 ;
      RECT 25.285000  25.240000 32.485000  25.310000 ;
      RECT 25.285000  25.240000 32.485000  25.310000 ;
      RECT 25.315000  43.005000 73.380000  43.075000 ;
      RECT 25.315000  43.005000 73.380000  43.075000 ;
      RECT 25.355000  25.310000 32.485000  25.380000 ;
      RECT 25.355000  25.310000 32.485000  25.380000 ;
      RECT 25.385000  42.935000 73.380000  43.005000 ;
      RECT 25.385000  42.935000 73.380000  43.005000 ;
      RECT 25.415000   3.515000 27.575000   3.585000 ;
      RECT 25.415000   3.585000 27.645000   3.655000 ;
      RECT 25.415000   3.655000 27.715000   3.725000 ;
      RECT 25.415000   3.725000 27.785000   3.795000 ;
      RECT 25.415000   3.795000 27.855000   3.845000 ;
      RECT 25.415000   3.845000 27.905000   4.385000 ;
      RECT 25.415000   4.385000 29.415000   4.455000 ;
      RECT 25.415000   4.455000 29.345000   4.525000 ;
      RECT 25.415000   4.525000 29.275000   4.595000 ;
      RECT 25.415000   4.595000 29.255000   4.615000 ;
      RECT 25.415000   4.615000 27.905000   5.825000 ;
      RECT 25.415000   5.825000 31.165000   6.800000 ;
      RECT 25.415000   5.825000 31.165000   8.950000 ;
      RECT 25.415000   5.825000 31.165000   8.950000 ;
      RECT 25.415000   5.825000 31.165000   8.950000 ;
      RECT 25.415000   6.800000 32.480000   8.945000 ;
      RECT 25.415000   8.945000 32.480000   8.950000 ;
      RECT 25.415000   8.945000 32.480000   8.950000 ;
      RECT 25.415000   8.950000 32.485000  12.360000 ;
      RECT 25.425000  25.380000 32.485000  25.450000 ;
      RECT 25.425000  25.380000 32.485000  25.450000 ;
      RECT 25.455000  25.675000 32.625000  28.070000 ;
      RECT 25.455000  28.070000 32.485000  28.210000 ;
      RECT 25.455000  28.210000 28.495000  28.480000 ;
      RECT 25.455000  28.480000 28.495000  32.575000 ;
      RECT 25.455000  32.575000 75.000000  42.670000 ;
      RECT 25.455000  42.670000 75.000000  43.685000 ;
      RECT 25.455000  42.865000 73.380000  42.935000 ;
      RECT 25.455000  42.865000 73.380000  42.935000 ;
      RECT 25.485000  12.360000 32.485000  12.430000 ;
      RECT 25.485000  12.360000 32.485000  12.430000 ;
      RECT 25.495000  25.450000 32.485000  25.520000 ;
      RECT 25.495000  25.450000 32.485000  25.520000 ;
      RECT 25.525000  12.665000 32.625000  14.975000 ;
      RECT 25.525000  14.975000 32.625000  15.475000 ;
      RECT 25.525000  42.795000 73.380000  42.865000 ;
      RECT 25.525000  42.795000 73.380000  42.865000 ;
      RECT 25.555000  12.430000 32.485000  12.500000 ;
      RECT 25.555000  12.430000 32.485000  12.500000 ;
      RECT 25.560000   0.185000 27.265000   3.235000 ;
      RECT 25.565000  25.520000 32.485000  25.590000 ;
      RECT 25.565000  25.520000 32.485000  25.590000 ;
      RECT 25.595000  25.590000 32.485000  25.620000 ;
      RECT 25.595000  25.590000 32.485000  25.620000 ;
      RECT 25.595000  25.620000 32.485000  28.015000 ;
      RECT 25.595000  28.015000 32.460000  28.040000 ;
      RECT 25.595000  28.015000 32.460000  28.040000 ;
      RECT 25.595000  28.040000 32.430000  28.070000 ;
      RECT 25.595000  28.040000 32.430000  28.070000 ;
      RECT 25.595000  28.070000 28.640000  28.140000 ;
      RECT 25.595000  28.070000 28.640000  28.140000 ;
      RECT 25.595000  28.140000 28.570000  28.210000 ;
      RECT 25.595000  28.140000 28.570000  28.210000 ;
      RECT 25.595000  28.210000 28.500000  28.280000 ;
      RECT 25.595000  28.210000 28.500000  28.280000 ;
      RECT 25.595000  28.280000 28.430000  28.350000 ;
      RECT 25.595000  28.280000 28.430000  28.350000 ;
      RECT 25.595000  28.350000 28.360000  28.420000 ;
      RECT 25.595000  28.350000 28.360000  28.420000 ;
      RECT 25.595000  28.420000 28.355000  28.425000 ;
      RECT 25.595000  28.420000 28.355000  28.425000 ;
      RECT 25.595000  28.425000 28.355000  32.715000 ;
      RECT 25.595000  32.715000 73.380000  42.725000 ;
      RECT 25.595000  42.725000 73.380000  42.795000 ;
      RECT 25.595000  42.725000 73.380000  42.795000 ;
      RECT 25.625000  12.500000 32.485000  12.570000 ;
      RECT 25.625000  12.500000 32.485000  12.570000 ;
      RECT 25.665000  12.570000 32.485000  12.610000 ;
      RECT 25.665000  12.570000 32.485000  12.610000 ;
      RECT 25.665000  12.610000 32.485000  14.920000 ;
      RECT 25.735000  14.920000 32.485000  14.990000 ;
      RECT 25.735000  14.920000 32.485000  14.990000 ;
      RECT 25.805000  14.990000 32.485000  15.060000 ;
      RECT 25.805000  14.990000 32.485000  15.060000 ;
      RECT 25.875000  15.060000 32.485000  15.130000 ;
      RECT 25.875000  15.060000 32.485000  15.130000 ;
      RECT 25.945000  15.130000 32.485000  15.200000 ;
      RECT 25.945000  15.130000 32.485000  15.200000 ;
      RECT 26.015000  15.200000 32.485000  15.270000 ;
      RECT 26.015000  15.200000 32.485000  15.270000 ;
      RECT 26.080000  15.270000 32.485000  15.335000 ;
      RECT 26.080000  15.270000 32.485000  15.335000 ;
      RECT 28.370000   0.000000 30.365000   2.795000 ;
      RECT 28.370000   2.795000 30.365000   3.400000 ;
      RECT 28.500000   0.185000 30.205000   2.395000 ;
      RECT 28.515000   2.675000 30.225000   2.745000 ;
      RECT 28.585000   2.745000 30.225000   2.815000 ;
      RECT 28.655000   2.815000 30.225000   2.885000 ;
      RECT 28.725000   2.885000 30.225000   2.955000 ;
      RECT 28.795000   2.955000 30.225000   3.025000 ;
      RECT 28.865000   3.025000 30.225000   3.095000 ;
      RECT 28.935000   3.095000 30.225000   3.165000 ;
      RECT 28.975000   3.400000 30.365000   3.700000 ;
      RECT 28.975000   3.700000 29.820000   4.245000 ;
      RECT 29.005000   3.165000 30.225000   3.235000 ;
      RECT 29.005000  28.790000 75.000000  32.575000 ;
      RECT 29.075000   3.235000 30.225000   3.305000 ;
      RECT 29.080000  28.720000 75.000000  28.790000 ;
      RECT 29.115000   3.305000 30.225000   3.345000 ;
      RECT 29.115000   3.345000 30.225000   3.645000 ;
      RECT 29.115000   3.645000 30.155000   3.715000 ;
      RECT 29.115000   3.715000 30.085000   3.785000 ;
      RECT 29.115000   3.785000 30.015000   3.855000 ;
      RECT 29.115000   3.855000 29.945000   3.925000 ;
      RECT 29.115000   3.925000 29.875000   3.995000 ;
      RECT 29.115000   3.995000 29.805000   4.065000 ;
      RECT 29.115000   4.065000 29.735000   4.135000 ;
      RECT 29.115000   4.135000 29.665000   4.205000 ;
      RECT 29.115000   4.205000 29.595000   4.275000 ;
      RECT 29.115000   4.275000 29.525000   4.345000 ;
      RECT 29.115000   4.345000 29.485000   4.385000 ;
      RECT 29.145000  28.860000 73.380000  32.715000 ;
      RECT 29.765000   5.815000 31.165000   5.825000 ;
      RECT 29.835000   5.745000 31.165000   5.815000 ;
      RECT 29.905000   5.675000 31.165000   5.745000 ;
      RECT 29.975000   5.605000 31.165000   5.675000 ;
      RECT 30.025000  15.475000 32.625000  16.625000 ;
      RECT 30.045000   5.535000 31.165000   5.605000 ;
      RECT 30.115000   5.465000 31.165000   5.535000 ;
      RECT 30.150000  15.335000 32.485000  15.405000 ;
      RECT 30.150000  15.335000 32.485000  15.405000 ;
      RECT 30.185000   5.395000 31.165000   5.465000 ;
      RECT 30.220000  15.405000 32.485000  15.475000 ;
      RECT 30.220000  15.405000 32.485000  15.475000 ;
      RECT 30.255000   5.325000 31.165000   5.395000 ;
      RECT 30.290000  15.475000 32.485000  15.545000 ;
      RECT 30.290000  15.475000 32.485000  15.545000 ;
      RECT 30.325000   5.255000 31.165000   5.325000 ;
      RECT 30.360000  15.545000 32.485000  15.615000 ;
      RECT 30.360000  15.545000 32.485000  15.615000 ;
      RECT 30.395000   5.185000 31.165000   5.255000 ;
      RECT 30.430000  15.615000 32.485000  15.685000 ;
      RECT 30.430000  15.615000 32.485000  15.685000 ;
      RECT 30.435000  80.155000 73.380000  84.520000 ;
      RECT 30.435000  84.520000 33.105000  84.755000 ;
      RECT 30.465000   5.115000 31.165000   5.185000 ;
      RECT 30.500000  15.685000 32.485000  15.755000 ;
      RECT 30.500000  15.685000 32.485000  15.755000 ;
      RECT 30.535000   5.045000 31.165000   5.115000 ;
      RECT 30.570000  15.755000 32.485000  15.825000 ;
      RECT 30.570000  15.755000 32.485000  15.825000 ;
      RECT 30.605000   4.975000 31.165000   5.045000 ;
      RECT 30.640000  15.825000 32.485000  15.895000 ;
      RECT 30.640000  15.825000 32.485000  15.895000 ;
      RECT 30.675000   4.905000 31.165000   4.975000 ;
      RECT 30.710000  15.895000 32.485000  15.965000 ;
      RECT 30.710000  15.895000 32.485000  15.965000 ;
      RECT 30.745000   4.835000 31.165000   4.905000 ;
      RECT 30.780000  15.965000 32.485000  16.035000 ;
      RECT 30.780000  15.965000 32.485000  16.035000 ;
      RECT 30.815000   4.765000 31.165000   4.835000 ;
      RECT 30.850000  16.035000 32.485000  16.105000 ;
      RECT 30.850000  16.035000 32.485000  16.105000 ;
      RECT 30.885000   4.695000 31.165000   4.765000 ;
      RECT 30.920000  16.105000 32.485000  16.175000 ;
      RECT 30.920000  16.105000 32.485000  16.175000 ;
      RECT 30.955000   4.625000 31.165000   4.695000 ;
      RECT 30.990000  16.175000 32.485000  16.245000 ;
      RECT 30.990000  16.175000 32.485000  16.245000 ;
      RECT 31.025000   4.555000 31.165000   4.625000 ;
      RECT 31.060000  16.245000 32.485000  16.315000 ;
      RECT 31.060000  16.245000 32.485000  16.315000 ;
      RECT 31.095000   4.485000 31.165000   4.555000 ;
      RECT 31.130000  16.315000 32.485000  16.385000 ;
      RECT 31.130000  16.315000 32.485000  16.385000 ;
      RECT 31.175000  16.625000 32.625000  19.485000 ;
      RECT 31.200000  16.385000 32.485000  16.455000 ;
      RECT 31.200000  16.385000 32.485000  16.455000 ;
      RECT 31.270000  16.455000 32.485000  16.525000 ;
      RECT 31.270000  16.455000 32.485000  16.525000 ;
      RECT 31.295000   0.000000 32.620000   4.090000 ;
      RECT 31.295000   4.090000 32.620000   5.685000 ;
      RECT 31.315000  16.525000 32.485000  16.570000 ;
      RECT 31.315000  16.525000 32.485000  16.570000 ;
      RECT 31.315000  16.570000 32.485000  19.625000 ;
      RECT 31.435000   0.000000 32.480000   0.390000 ;
      RECT 31.445000   0.670000 32.410000   6.520000 ;
      RECT 33.160000   0.000000 75.000000   8.660000 ;
      RECT 33.160000   8.660000 75.000000   8.665000 ;
      RECT 33.165000   8.665000 75.000000  28.720000 ;
      RECT 33.300000   0.000000 75.000000   0.600000 ;
      RECT 33.300000   0.600000 34.820000   0.620000 ;
      RECT 33.300000   0.620000 34.615000   2.160000 ;
      RECT 33.300000   2.160000 39.940000   6.270000 ;
      RECT 33.300000   6.270000 73.110000   6.340000 ;
      RECT 33.300000   6.270000 73.110000   6.340000 ;
      RECT 33.300000   6.340000 73.180000   6.410000 ;
      RECT 33.300000   6.340000 73.180000   6.410000 ;
      RECT 33.300000   6.410000 73.250000   6.480000 ;
      RECT 33.300000   6.410000 73.250000   6.480000 ;
      RECT 33.300000   6.480000 73.320000   6.540000 ;
      RECT 33.300000   6.480000 73.320000   6.540000 ;
      RECT 33.300000   6.540000 73.380000   8.605000 ;
      RECT 33.305000   8.605000 73.380000   8.610000 ;
      RECT 33.305000   8.605000 73.380000   8.610000 ;
      RECT 33.305000   8.610000 73.380000  28.860000 ;
      RECT 33.305000   8.610000 73.380000  32.715000 ;
      RECT 33.385000  84.800000 74.700000  85.055000 ;
      RECT 34.895000   0.900000 38.965000   1.880000 ;
      RECT 35.100000   0.880000 38.920000   0.900000 ;
      RECT 39.200000   0.600000 75.000000   0.620000 ;
      RECT 39.245000   0.620000 75.000000   0.740000 ;
      RECT 39.245000   0.740000 39.940000   2.160000 ;
      RECT 40.220000   1.020000 74.590000   5.990000 ;
      RECT 56.545000 100.330000 72.090000 101.420000 ;
      RECT 56.725000  97.530000 72.090000  97.760000 ;
      RECT 56.825000  98.040000 71.245000  98.110000 ;
      RECT 56.825000  98.110000 71.315000  98.180000 ;
      RECT 56.825000  98.180000 71.385000  98.250000 ;
      RECT 56.825000  98.250000 71.455000  98.320000 ;
      RECT 56.825000  98.320000 71.525000  98.390000 ;
      RECT 56.825000  98.390000 71.595000  98.460000 ;
      RECT 56.825000  98.460000 71.665000  98.530000 ;
      RECT 56.825000  98.530000 71.735000  98.600000 ;
      RECT 56.825000  98.600000 71.805000  98.605000 ;
      RECT 56.825000  98.605000 71.810000  99.405000 ;
      RECT 56.825000  99.405000 71.740000  99.475000 ;
      RECT 56.825000  99.475000 71.670000  99.545000 ;
      RECT 56.825000  99.545000 71.600000  99.615000 ;
      RECT 56.825000  99.615000 71.530000  99.685000 ;
      RECT 56.825000  99.685000 71.460000  99.755000 ;
      RECT 56.825000  99.755000 71.390000  99.825000 ;
      RECT 56.825000  99.825000 71.320000  99.895000 ;
      RECT 56.825000  99.895000 71.250000  99.965000 ;
      RECT 56.825000  99.965000 71.180000 100.035000 ;
      RECT 56.825000 100.035000 71.165000 100.050000 ;
      RECT 59.500000 199.490000 64.600000 200.000000 ;
      RECT 59.780000 196.250000 64.320000 199.210000 ;
      RECT 60.320000 125.440000 75.145000 125.510000 ;
      RECT 60.320000 125.440000 75.145000 125.510000 ;
      RECT 60.390000 125.510000 75.145000 125.580000 ;
      RECT 60.390000 125.510000 75.145000 125.580000 ;
      RECT 60.460000 125.580000 75.145000 125.650000 ;
      RECT 60.460000 125.580000 75.145000 125.650000 ;
      RECT 60.530000 125.650000 75.145000 125.720000 ;
      RECT 60.530000 125.650000 75.145000 125.720000 ;
      RECT 60.600000 125.720000 75.145000 125.790000 ;
      RECT 60.600000 125.720000 75.145000 125.790000 ;
      RECT 60.670000 125.790000 75.145000 125.860000 ;
      RECT 60.670000 125.790000 75.145000 125.860000 ;
      RECT 60.740000 125.860000 75.145000 125.930000 ;
      RECT 60.740000 125.860000 75.145000 125.930000 ;
      RECT 60.810000 125.930000 75.145000 126.000000 ;
      RECT 60.810000 125.930000 75.145000 126.000000 ;
      RECT 60.880000 126.000000 75.145000 126.070000 ;
      RECT 60.880000 126.000000 75.145000 126.070000 ;
      RECT 60.950000 126.070000 75.145000 126.140000 ;
      RECT 60.950000 126.070000 75.145000 126.140000 ;
      RECT 61.020000 126.140000 75.145000 126.210000 ;
      RECT 61.020000 126.140000 75.145000 126.210000 ;
      RECT 61.090000 126.210000 75.145000 126.280000 ;
      RECT 61.090000 126.210000 75.145000 126.280000 ;
      RECT 61.160000 126.280000 75.145000 126.350000 ;
      RECT 61.160000 126.280000 75.145000 126.350000 ;
      RECT 61.230000 126.350000 75.145000 126.420000 ;
      RECT 61.230000 126.350000 75.145000 126.420000 ;
      RECT 61.300000 126.420000 75.145000 126.490000 ;
      RECT 61.300000 126.420000 75.145000 126.490000 ;
      RECT 61.370000 126.490000 75.145000 126.560000 ;
      RECT 61.370000 126.490000 75.145000 126.560000 ;
      RECT 61.440000 126.560000 75.145000 126.630000 ;
      RECT 61.440000 126.560000 75.145000 126.630000 ;
      RECT 61.510000 126.630000 75.145000 126.700000 ;
      RECT 61.510000 126.630000 75.145000 126.700000 ;
      RECT 61.580000 126.700000 75.145000 126.770000 ;
      RECT 61.580000 126.700000 75.145000 126.770000 ;
      RECT 61.650000 126.770000 75.145000 126.840000 ;
      RECT 61.650000 126.770000 75.145000 126.840000 ;
      RECT 61.720000 126.840000 75.145000 126.910000 ;
      RECT 61.720000 126.840000 75.145000 126.910000 ;
      RECT 61.790000 126.910000 75.145000 126.980000 ;
      RECT 61.790000 126.910000 75.145000 126.980000 ;
      RECT 61.860000 126.980000 75.145000 127.050000 ;
      RECT 61.860000 126.980000 75.145000 127.050000 ;
      RECT 61.930000 127.050000 75.145000 127.120000 ;
      RECT 61.930000 127.050000 75.145000 127.120000 ;
      RECT 62.000000 127.120000 75.145000 127.190000 ;
      RECT 62.000000 127.120000 75.145000 127.190000 ;
      RECT 62.070000 127.190000 75.145000 127.260000 ;
      RECT 62.070000 127.190000 75.145000 127.260000 ;
      RECT 62.140000 127.260000 75.145000 127.330000 ;
      RECT 62.140000 127.260000 75.145000 127.330000 ;
      RECT 62.210000 127.330000 75.145000 127.400000 ;
      RECT 62.210000 127.330000 75.145000 127.400000 ;
      RECT 62.280000 127.400000 75.145000 127.470000 ;
      RECT 62.280000 127.400000 75.145000 127.470000 ;
      RECT 62.350000 127.470000 75.145000 127.540000 ;
      RECT 62.350000 127.470000 75.145000 127.540000 ;
      RECT 62.420000 127.540000 75.145000 127.610000 ;
      RECT 62.420000 127.540000 75.145000 127.610000 ;
      RECT 62.490000 127.610000 75.145000 127.680000 ;
      RECT 62.490000 127.610000 75.145000 127.680000 ;
      RECT 62.560000 127.680000 75.145000 127.750000 ;
      RECT 62.560000 127.680000 75.145000 127.750000 ;
      RECT 62.630000 127.750000 75.145000 127.820000 ;
      RECT 62.630000 127.750000 75.145000 127.820000 ;
      RECT 62.700000 127.820000 75.145000 127.890000 ;
      RECT 62.700000 127.820000 75.145000 127.890000 ;
      RECT 62.770000 127.890000 75.145000 127.960000 ;
      RECT 62.770000 127.890000 75.145000 127.960000 ;
      RECT 62.840000 127.960000 75.145000 128.030000 ;
      RECT 62.840000 127.960000 75.145000 128.030000 ;
      RECT 62.910000 128.030000 75.145000 128.100000 ;
      RECT 62.910000 128.030000 75.145000 128.100000 ;
      RECT 62.980000 128.100000 75.145000 128.170000 ;
      RECT 62.980000 128.100000 75.145000 128.170000 ;
      RECT 63.050000 128.170000 75.145000 128.240000 ;
      RECT 63.050000 128.170000 75.145000 128.240000 ;
      RECT 63.070000 128.240000 75.145000 128.260000 ;
      RECT 63.070000 128.240000 75.145000 128.260000 ;
      RECT 63.140000 128.260000 75.145000 128.330000 ;
      RECT 63.140000 128.260000 75.145000 128.330000 ;
      RECT 63.210000 128.330000 75.145000 128.400000 ;
      RECT 63.210000 128.330000 75.145000 128.400000 ;
      RECT 63.280000 128.400000 75.145000 128.470000 ;
      RECT 63.280000 128.400000 75.145000 128.470000 ;
      RECT 63.350000 128.470000 75.145000 128.540000 ;
      RECT 63.350000 128.470000 75.145000 128.540000 ;
      RECT 63.420000 128.540000 75.145000 128.610000 ;
      RECT 63.420000 128.540000 75.145000 128.610000 ;
      RECT 63.490000 128.610000 75.145000 128.680000 ;
      RECT 63.490000 128.610000 75.145000 128.680000 ;
      RECT 63.560000 128.680000 75.145000 128.750000 ;
      RECT 63.560000 128.680000 75.145000 128.750000 ;
      RECT 63.630000 128.750000 75.145000 128.820000 ;
      RECT 63.630000 128.750000 75.145000 128.820000 ;
      RECT 63.700000 128.820000 75.145000 128.890000 ;
      RECT 63.700000 128.820000 75.145000 128.890000 ;
      RECT 63.770000 128.890000 75.145000 128.960000 ;
      RECT 63.770000 128.890000 75.145000 128.960000 ;
      RECT 63.840000 128.960000 75.145000 129.030000 ;
      RECT 63.840000 128.960000 75.145000 129.030000 ;
      RECT 63.910000 129.030000 75.145000 129.100000 ;
      RECT 63.910000 129.030000 75.145000 129.100000 ;
      RECT 63.980000 129.100000 75.145000 129.170000 ;
      RECT 63.980000 129.100000 75.145000 129.170000 ;
      RECT 64.050000 129.170000 75.145000 129.240000 ;
      RECT 64.050000 129.170000 75.145000 129.240000 ;
      RECT 64.120000 129.240000 75.145000 129.310000 ;
      RECT 64.120000 129.240000 75.145000 129.310000 ;
      RECT 64.190000 129.310000 75.145000 129.380000 ;
      RECT 64.190000 129.310000 75.145000 129.380000 ;
      RECT 64.260000 129.380000 75.145000 129.450000 ;
      RECT 64.260000 129.380000 75.145000 129.450000 ;
      RECT 64.330000 129.450000 75.145000 129.520000 ;
      RECT 64.330000 129.450000 75.145000 129.520000 ;
      RECT 64.400000 129.520000 75.145000 129.590000 ;
      RECT 64.400000 129.520000 75.145000 129.590000 ;
      RECT 64.470000 129.590000 75.145000 129.660000 ;
      RECT 64.470000 129.590000 75.145000 129.660000 ;
      RECT 64.540000 129.660000 75.145000 129.730000 ;
      RECT 64.540000 129.660000 75.145000 129.730000 ;
      RECT 64.600000 175.420000 75.000000 200.000000 ;
      RECT 64.600000 195.970000 75.000000 199.490000 ;
      RECT 64.600000 199.490000 75.000000 200.000000 ;
      RECT 64.610000 129.730000 75.145000 129.800000 ;
      RECT 64.610000 129.730000 75.145000 129.800000 ;
      RECT 64.680000 129.800000 75.145000 129.870000 ;
      RECT 64.680000 129.800000 75.145000 129.870000 ;
      RECT 64.750000 129.870000 75.145000 129.940000 ;
      RECT 64.750000 129.870000 75.145000 129.940000 ;
      RECT 64.820000 129.940000 75.145000 130.010000 ;
      RECT 64.820000 129.940000 75.145000 130.010000 ;
      RECT 64.890000 130.010000 75.145000 130.080000 ;
      RECT 64.890000 130.010000 75.145000 130.080000 ;
      RECT 64.960000 130.080000 75.145000 130.150000 ;
      RECT 64.960000 130.080000 75.145000 130.150000 ;
      RECT 65.030000 130.150000 75.145000 130.220000 ;
      RECT 65.030000 130.150000 75.145000 130.220000 ;
      RECT 69.105000 138.955000 75.145000 138.960000 ;
      RECT 69.105000 138.955000 75.145000 138.960000 ;
      RECT 69.110000 138.950000 75.145000 138.955000 ;
      RECT 69.110000 138.950000 75.145000 138.955000 ;
      RECT 69.115000 138.945000 75.145000 138.950000 ;
      RECT 69.115000 138.945000 75.145000 138.950000 ;
      RECT 69.115000 138.960000 75.145000 138.975000 ;
      RECT 69.115000 138.960000 75.145000 138.975000 ;
      RECT 69.130000 138.975000 75.145000 138.990000 ;
      RECT 69.130000 138.975000 75.145000 138.990000 ;
      RECT 69.160000 138.900000 75.145000 138.945000 ;
      RECT 69.160000 138.900000 75.145000 138.945000 ;
      RECT 69.200000 138.990000 75.145000 139.060000 ;
      RECT 69.200000 138.990000 75.145000 139.060000 ;
      RECT 69.230000 138.830000 75.145000 138.900000 ;
      RECT 69.230000 138.830000 75.145000 138.900000 ;
      RECT 69.270000 139.060000 75.145000 139.130000 ;
      RECT 69.270000 139.060000 75.145000 139.130000 ;
      RECT 69.300000 138.760000 75.145000 138.830000 ;
      RECT 69.300000 138.760000 75.145000 138.830000 ;
      RECT 69.340000 139.130000 75.145000 139.200000 ;
      RECT 69.340000 139.130000 75.145000 139.200000 ;
      RECT 69.370000 138.690000 75.145000 138.760000 ;
      RECT 69.370000 138.690000 75.145000 138.760000 ;
      RECT 69.410000 139.200000 75.145000 139.270000 ;
      RECT 69.410000 139.200000 75.145000 139.270000 ;
      RECT 69.440000 138.620000 75.145000 138.690000 ;
      RECT 69.440000 138.620000 75.145000 138.690000 ;
      RECT 69.480000 139.270000 75.145000 139.340000 ;
      RECT 69.480000 139.270000 75.145000 139.340000 ;
      RECT 69.510000 138.550000 75.145000 138.620000 ;
      RECT 69.510000 138.550000 75.145000 138.620000 ;
      RECT 69.550000 139.340000 75.145000 139.410000 ;
      RECT 69.550000 139.340000 75.145000 139.410000 ;
      RECT 69.580000 138.480000 75.145000 138.550000 ;
      RECT 69.580000 138.480000 75.145000 138.550000 ;
      RECT 69.620000 139.410000 75.145000 139.480000 ;
      RECT 69.620000 139.410000 75.145000 139.480000 ;
      RECT 69.650000 138.410000 75.145000 138.480000 ;
      RECT 69.650000 138.410000 75.145000 138.480000 ;
      RECT 69.690000 139.480000 75.145000 139.550000 ;
      RECT 69.690000 139.480000 75.145000 139.550000 ;
      RECT 69.715000 139.550000 75.145000 139.575000 ;
      RECT 69.715000 139.550000 75.145000 139.575000 ;
      RECT 69.720000 138.340000 75.145000 138.410000 ;
      RECT 69.720000 138.340000 75.145000 138.410000 ;
      RECT 69.785000 139.575000 75.145000 139.645000 ;
      RECT 69.785000 139.575000 75.145000 139.645000 ;
      RECT 69.790000 138.270000 75.145000 138.340000 ;
      RECT 69.790000 138.270000 75.145000 138.340000 ;
      RECT 69.855000 139.645000 75.145000 139.715000 ;
      RECT 69.855000 139.645000 75.145000 139.715000 ;
      RECT 69.860000 138.200000 75.145000 138.270000 ;
      RECT 69.860000 138.200000 75.145000 138.270000 ;
      RECT 69.925000 139.715000 75.145000 139.785000 ;
      RECT 69.925000 139.715000 75.145000 139.785000 ;
      RECT 69.925000 141.095000 70.525000 143.875000 ;
      RECT 69.930000 138.130000 75.145000 138.200000 ;
      RECT 69.930000 138.130000 75.145000 138.200000 ;
      RECT 69.990000 139.785000 75.145000 139.850000 ;
      RECT 69.990000 139.785000 75.145000 139.850000 ;
      RECT 70.000000 138.060000 75.145000 138.130000 ;
      RECT 70.000000 138.060000 75.145000 138.130000 ;
      RECT 70.060000 139.850000 75.145000 139.920000 ;
      RECT 70.060000 139.850000 75.145000 139.920000 ;
      RECT 70.070000 137.990000 75.145000 138.060000 ;
      RECT 70.070000 137.990000 75.145000 138.060000 ;
      RECT 70.105000 145.100000 75.145000 145.130000 ;
      RECT 70.130000 139.920000 75.145000 139.990000 ;
      RECT 70.130000 139.920000 75.145000 139.990000 ;
      RECT 70.140000 137.920000 75.145000 137.990000 ;
      RECT 70.140000 137.920000 75.145000 137.990000 ;
      RECT 70.175000 145.030000 75.145000 145.100000 ;
      RECT 70.200000 139.990000 75.145000 140.060000 ;
      RECT 70.200000 139.990000 75.145000 140.060000 ;
      RECT 70.210000 137.850000 75.145000 137.920000 ;
      RECT 70.210000 137.850000 75.145000 137.920000 ;
      RECT 70.245000 144.960000 75.145000 145.030000 ;
      RECT 70.270000 140.060000 75.145000 140.130000 ;
      RECT 70.270000 140.060000 75.145000 140.130000 ;
      RECT 70.280000 137.780000 75.145000 137.850000 ;
      RECT 70.280000 137.780000 75.145000 137.850000 ;
      RECT 70.315000 144.890000 75.145000 144.960000 ;
      RECT 70.340000 140.130000 75.145000 140.200000 ;
      RECT 70.340000 140.130000 75.145000 140.200000 ;
      RECT 70.350000 137.710000 75.145000 137.780000 ;
      RECT 70.350000 137.710000 75.145000 137.780000 ;
      RECT 70.385000 144.820000 75.145000 144.890000 ;
      RECT 70.410000 140.200000 75.145000 140.270000 ;
      RECT 70.410000 140.200000 75.145000 140.270000 ;
      RECT 70.420000 137.640000 75.145000 137.710000 ;
      RECT 70.420000 137.640000 75.145000 137.710000 ;
      RECT 70.455000 144.750000 75.145000 144.820000 ;
      RECT 70.480000 140.270000 75.145000 140.340000 ;
      RECT 70.480000 140.270000 75.145000 140.340000 ;
      RECT 70.490000 137.570000 75.145000 137.640000 ;
      RECT 70.490000 137.570000 75.145000 137.640000 ;
      RECT 70.525000 144.680000 75.145000 144.750000 ;
      RECT 70.550000 140.340000 75.145000 140.410000 ;
      RECT 70.550000 140.340000 75.145000 140.410000 ;
      RECT 70.560000 137.500000 75.145000 137.570000 ;
      RECT 70.560000 137.500000 75.145000 137.570000 ;
      RECT 70.595000 144.610000 75.145000 144.680000 ;
      RECT 70.620000 140.410000 75.145000 140.480000 ;
      RECT 70.620000 140.410000 75.145000 140.480000 ;
      RECT 70.630000 137.430000 75.145000 137.500000 ;
      RECT 70.630000 137.430000 75.145000 137.500000 ;
      RECT 70.665000 144.540000 75.145000 144.610000 ;
      RECT 70.690000 140.480000 75.145000 140.550000 ;
      RECT 70.690000 140.480000 75.145000 140.550000 ;
      RECT 70.700000 137.360000 75.145000 137.430000 ;
      RECT 70.700000 137.360000 75.145000 137.430000 ;
      RECT 70.735000 144.470000 75.145000 144.540000 ;
      RECT 70.760000 140.550000 75.145000 140.620000 ;
      RECT 70.760000 140.550000 75.145000 140.620000 ;
      RECT 70.770000 137.290000 75.145000 137.360000 ;
      RECT 70.770000 137.290000 75.145000 137.360000 ;
      RECT 70.805000 139.850000 75.145000 145.130000 ;
      RECT 70.805000 140.620000 75.145000 140.665000 ;
      RECT 70.805000 140.620000 75.145000 140.665000 ;
      RECT 70.805000 140.665000 75.145000 144.400000 ;
      RECT 70.805000 144.400000 75.145000 144.470000 ;
      RECT 70.805000 144.400000 75.145000 145.130000 ;
      RECT 70.805000 145.130000 73.195000 146.145000 ;
      RECT 70.840000 137.220000 75.145000 137.290000 ;
      RECT 70.840000 137.220000 75.145000 137.290000 ;
      RECT 70.910000 137.150000 75.145000 137.220000 ;
      RECT 70.910000 137.150000 75.145000 137.220000 ;
      RECT 70.980000 137.080000 75.145000 137.150000 ;
      RECT 70.980000 137.080000 75.145000 137.150000 ;
      RECT 71.050000 137.010000 75.145000 137.080000 ;
      RECT 71.050000 137.010000 75.145000 137.080000 ;
      RECT 71.120000 136.940000 75.145000 137.010000 ;
      RECT 71.120000 136.940000 75.145000 137.010000 ;
      RECT 71.190000 136.870000 75.145000 136.940000 ;
      RECT 71.190000 136.870000 75.145000 136.940000 ;
      RECT 71.260000 136.800000 75.145000 136.870000 ;
      RECT 71.260000 136.800000 75.145000 136.870000 ;
      RECT 71.320000 100.290000 75.145000 100.330000 ;
      RECT 71.330000 136.730000 75.145000 136.800000 ;
      RECT 71.330000 136.730000 75.145000 136.800000 ;
      RECT 71.390000 100.220000 75.145000 100.290000 ;
      RECT 71.400000 136.660000 75.145000 136.730000 ;
      RECT 71.400000 136.660000 75.145000 136.730000 ;
      RECT 71.430000  97.760000 75.145000  97.830000 ;
      RECT 71.460000 100.150000 75.145000 100.220000 ;
      RECT 71.470000 136.590000 75.145000 136.660000 ;
      RECT 71.470000 136.590000 75.145000 136.660000 ;
      RECT 71.500000  97.830000 75.145000  97.900000 ;
      RECT 71.530000 100.080000 75.145000 100.150000 ;
      RECT 71.540000 136.520000 75.145000 136.590000 ;
      RECT 71.540000 136.520000 75.145000 136.590000 ;
      RECT 71.570000  97.900000 75.145000  97.970000 ;
      RECT 71.600000 100.010000 75.145000 100.080000 ;
      RECT 71.610000 136.450000 75.145000 136.520000 ;
      RECT 71.610000 136.450000 75.145000 136.520000 ;
      RECT 71.640000  97.970000 75.145000  98.040000 ;
      RECT 71.670000  99.940000 75.145000 100.010000 ;
      RECT 71.680000 136.380000 75.145000 136.450000 ;
      RECT 71.680000 136.380000 75.145000 136.450000 ;
      RECT 71.710000  98.040000 75.145000  98.110000 ;
      RECT 71.740000  99.870000 75.145000  99.940000 ;
      RECT 71.750000 136.310000 75.145000 136.380000 ;
      RECT 71.750000 136.310000 75.145000 136.380000 ;
      RECT 71.755000  85.835000 74.700000  94.470000 ;
      RECT 71.780000  98.110000 75.145000  98.180000 ;
      RECT 71.810000  99.800000 75.145000  99.870000 ;
      RECT 71.820000 136.240000 75.145000 136.310000 ;
      RECT 71.820000 136.240000 75.145000 136.310000 ;
      RECT 71.850000  98.180000 75.145000  98.250000 ;
      RECT 71.880000  99.730000 75.145000  99.800000 ;
      RECT 71.890000 136.170000 75.145000 136.240000 ;
      RECT 71.890000 136.170000 75.145000 136.240000 ;
      RECT 71.920000  98.250000 75.145000  98.320000 ;
      RECT 71.950000  99.660000 75.145000  99.730000 ;
      RECT 71.960000 136.100000 75.145000 136.170000 ;
      RECT 71.960000 136.100000 75.145000 136.170000 ;
      RECT 71.990000  98.320000 75.145000  98.390000 ;
      RECT 72.020000  99.590000 75.145000  99.660000 ;
      RECT 72.030000 136.030000 75.145000 136.100000 ;
      RECT 72.030000 136.030000 75.145000 136.100000 ;
      RECT 72.060000  98.390000 75.145000  98.460000 ;
      RECT 72.090000  97.530000 75.145000 100.765000 ;
      RECT 72.090000  97.760000 75.145000  98.490000 ;
      RECT 72.090000  98.460000 75.145000  98.490000 ;
      RECT 72.090000  98.490000 75.145000  99.520000 ;
      RECT 72.090000  99.520000 75.145000  99.590000 ;
      RECT 72.090000  99.520000 75.145000 100.330000 ;
      RECT 72.090000 100.330000 75.145000 101.420000 ;
      RECT 72.100000 135.960000 75.145000 136.030000 ;
      RECT 72.100000 135.960000 75.145000 136.030000 ;
      RECT 72.115000  97.505000 75.145000  97.530000 ;
      RECT 72.170000 135.890000 75.145000 135.960000 ;
      RECT 72.170000 135.890000 75.145000 135.960000 ;
      RECT 72.185000  97.435000 75.145000  97.505000 ;
      RECT 72.240000 135.820000 75.145000 135.890000 ;
      RECT 72.240000 135.820000 75.145000 135.890000 ;
      RECT 72.255000  97.365000 75.145000  97.435000 ;
      RECT 72.310000 135.750000 75.145000 135.820000 ;
      RECT 72.310000 135.750000 75.145000 135.820000 ;
      RECT 72.325000  97.295000 75.145000  97.365000 ;
      RECT 72.380000 130.500000 75.000000 130.995000 ;
      RECT 72.380000 135.680000 75.145000 135.750000 ;
      RECT 72.380000 135.680000 75.145000 135.750000 ;
      RECT 72.395000  97.225000 75.145000  97.295000 ;
      RECT 72.450000 135.610000 75.145000 135.680000 ;
      RECT 72.450000 135.610000 75.145000 135.680000 ;
      RECT 72.465000  97.155000 75.145000  97.225000 ;
      RECT 72.520000 135.540000 75.145000 135.610000 ;
      RECT 72.520000 135.540000 75.145000 135.610000 ;
      RECT 72.535000  97.085000 75.145000  97.155000 ;
      RECT 72.590000 135.470000 75.145000 135.540000 ;
      RECT 72.590000 135.470000 75.145000 135.540000 ;
      RECT 72.605000  97.015000 75.145000  97.085000 ;
      RECT 72.660000 131.275000 75.145000 132.915000 ;
      RECT 72.660000 135.400000 75.145000 135.470000 ;
      RECT 72.660000 135.400000 75.145000 135.470000 ;
      RECT 72.675000  96.945000 75.145000  97.015000 ;
      RECT 72.695000 135.365000 75.145000 135.400000 ;
      RECT 72.695000 135.365000 75.145000 135.400000 ;
      RECT 72.745000  96.875000 75.145000  96.945000 ;
      RECT 72.765000 135.295000 75.145000 135.365000 ;
      RECT 72.765000 135.295000 75.145000 135.365000 ;
      RECT 72.815000  96.805000 75.145000  96.875000 ;
      RECT 72.835000 135.225000 75.145000 135.295000 ;
      RECT 72.835000 135.225000 75.145000 135.295000 ;
      RECT 72.885000  96.735000 75.145000  96.805000 ;
      RECT 72.905000 135.155000 75.145000 135.225000 ;
      RECT 72.905000 135.155000 75.145000 135.225000 ;
      RECT 72.955000  96.665000 75.145000  96.735000 ;
      RECT 72.975000 135.085000 75.145000 135.155000 ;
      RECT 72.975000 135.085000 75.145000 135.155000 ;
      RECT 73.025000  96.595000 75.145000  96.665000 ;
      RECT 73.045000 135.015000 75.145000 135.085000 ;
      RECT 73.045000 135.015000 75.145000 135.085000 ;
      RECT 73.095000  96.525000 75.145000  96.595000 ;
      RECT 73.115000 134.945000 75.145000 135.015000 ;
      RECT 73.115000 134.945000 75.145000 135.015000 ;
      RECT 73.165000  96.455000 75.145000  96.525000 ;
      RECT 73.185000 134.875000 75.145000 134.945000 ;
      RECT 73.185000 134.875000 75.145000 134.945000 ;
      RECT 73.235000  96.385000 75.145000  96.455000 ;
      RECT 73.255000 134.805000 75.145000 134.875000 ;
      RECT 73.255000 134.805000 75.145000 134.875000 ;
      RECT 73.295000   5.990000 74.590000   6.060000 ;
      RECT 73.305000  96.315000 75.145000  96.385000 ;
      RECT 73.325000 134.735000 75.145000 134.805000 ;
      RECT 73.325000 134.735000 75.145000 134.805000 ;
      RECT 73.365000   6.060000 74.590000   6.130000 ;
      RECT 73.375000  96.245000 75.145000  96.315000 ;
      RECT 73.395000 134.665000 75.145000 134.735000 ;
      RECT 73.395000 134.665000 75.145000 134.735000 ;
      RECT 73.435000   6.130000 74.590000   6.200000 ;
      RECT 73.445000  96.175000 75.145000  96.245000 ;
      RECT 73.465000 134.595000 75.145000 134.665000 ;
      RECT 73.465000 134.595000 75.145000 134.665000 ;
      RECT 73.475000 145.410000 75.000000 146.425000 ;
      RECT 73.505000   6.200000 74.590000   6.270000 ;
      RECT 73.515000  96.105000 75.145000  96.175000 ;
      RECT 73.535000 134.525000 75.145000 134.595000 ;
      RECT 73.535000 134.525000 75.145000 134.595000 ;
      RECT 73.575000   6.270000 74.590000   6.340000 ;
      RECT 73.585000  96.035000 75.145000  96.105000 ;
      RECT 73.605000 134.455000 75.145000 134.525000 ;
      RECT 73.605000 134.455000 75.145000 134.525000 ;
      RECT 73.645000   6.340000 74.590000   6.410000 ;
      RECT 73.655000  95.965000 75.145000  96.035000 ;
      RECT 73.660000   6.410000 74.590000   6.425000 ;
      RECT 73.660000   6.425000 74.590000  79.620000 ;
      RECT 73.660000  79.620000 74.590000  79.675000 ;
      RECT 73.660000  79.675000 74.645000  79.730000 ;
      RECT 73.660000  79.730000 74.700000  84.800000 ;
      RECT 73.675000 134.385000 75.145000 134.455000 ;
      RECT 73.675000 134.385000 75.145000 134.455000 ;
      RECT 73.685000 174.500000 74.745000 175.140000 ;
      RECT 73.725000  95.895000 75.145000  95.965000 ;
      RECT 73.725000  95.895000 75.145000 100.535000 ;
      RECT 73.745000 134.315000 75.145000 134.385000 ;
      RECT 73.745000 134.315000 75.145000 134.385000 ;
      RECT 73.770000 101.420000 74.700000 104.565000 ;
      RECT 73.815000 134.245000 75.145000 134.315000 ;
      RECT 73.815000 134.245000 75.145000 134.315000 ;
      RECT 73.885000 134.175000 75.145000 134.245000 ;
      RECT 73.885000 134.175000 75.145000 134.245000 ;
      RECT 73.955000 134.105000 75.145000 134.175000 ;
      RECT 73.955000 134.105000 75.145000 134.175000 ;
      RECT 74.025000 134.035000 75.145000 134.105000 ;
      RECT 74.025000 134.035000 75.145000 134.105000 ;
      RECT 74.035000 104.845000 75.000000 105.150000 ;
      RECT 74.095000 133.965000 75.145000 134.035000 ;
      RECT 74.095000 133.965000 75.145000 134.035000 ;
      RECT 74.165000 133.895000 75.145000 133.965000 ;
      RECT 74.165000 133.895000 75.145000 133.965000 ;
      RECT 74.235000 133.825000 75.145000 133.895000 ;
      RECT 74.235000 133.825000 75.145000 133.895000 ;
      RECT 74.305000 133.755000 75.145000 133.825000 ;
      RECT 74.305000 133.755000 75.145000 133.825000 ;
      RECT 74.315000 105.430000 74.915000 125.440000 ;
      RECT 74.375000 133.685000 75.145000 133.755000 ;
      RECT 74.375000 133.685000 75.145000 133.755000 ;
      RECT 74.445000 133.615000 75.145000 133.685000 ;
      RECT 74.445000 133.615000 75.145000 133.685000 ;
      RECT 74.515000 133.545000 75.145000 133.615000 ;
      RECT 74.515000 133.545000 75.145000 133.615000 ;
      RECT 74.585000 133.475000 75.145000 133.545000 ;
      RECT 74.585000 133.475000 75.145000 133.545000 ;
      RECT 74.655000 133.405000 75.145000 133.475000 ;
      RECT 74.655000 133.405000 75.145000 133.475000 ;
      RECT 74.725000 133.335000 75.145000 133.405000 ;
      RECT 74.725000 133.335000 75.145000 133.405000 ;
      RECT 74.795000 133.265000 75.145000 133.335000 ;
      RECT 74.795000 133.265000 75.145000 133.335000 ;
      RECT 74.855000 102.200000 74.925000 102.270000 ;
      RECT 74.855000 102.270000 74.995000 102.340000 ;
      RECT 74.855000 102.340000 75.065000 102.410000 ;
      RECT 74.855000 102.410000 75.135000 102.420000 ;
      RECT 74.865000 133.195000 75.145000 133.265000 ;
      RECT 74.865000 133.195000 75.145000 133.265000 ;
      RECT 74.935000 133.125000 75.145000 133.195000 ;
      RECT 74.935000 133.125000 75.145000 133.195000 ;
      RECT 75.005000 133.055000 75.145000 133.125000 ;
      RECT 75.005000 133.055000 75.145000 133.125000 ;
      RECT 75.075000 132.985000 75.145000 133.055000 ;
      RECT 75.075000 132.985000 75.145000 133.055000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  8.145000   4.405000 ;
      RECT  0.000000   0.000000  8.285000   1.320000 ;
      RECT  0.000000   1.320000 12.145000   1.610000 ;
      RECT  0.000000   1.610000 17.105000   3.275000 ;
      RECT  0.000000   3.155000 10.635000   3.225000 ;
      RECT  0.000000   3.225000 10.565000   3.295000 ;
      RECT  0.000000   3.275000 19.935000   3.295000 ;
      RECT  0.000000   3.295000  9.595000   4.460000 ;
      RECT  0.000000   3.295000 10.495000   3.365000 ;
      RECT  0.000000   3.365000 10.425000   3.435000 ;
      RECT  0.000000   3.435000 10.355000   3.505000 ;
      RECT  0.000000   3.505000 10.285000   3.575000 ;
      RECT  0.000000   3.575000 10.215000   3.645000 ;
      RECT  0.000000   3.645000 10.145000   3.715000 ;
      RECT  0.000000   3.715000 10.075000   3.785000 ;
      RECT  0.000000   3.785000 10.005000   3.855000 ;
      RECT  0.000000   3.855000  9.935000   3.925000 ;
      RECT  0.000000   3.925000  9.865000   3.995000 ;
      RECT  0.000000   3.995000  9.795000   4.065000 ;
      RECT  0.000000   4.065000  9.725000   4.135000 ;
      RECT  0.000000   4.135000  9.655000   4.205000 ;
      RECT  0.000000   4.205000  9.585000   4.275000 ;
      RECT  0.000000   4.275000  9.515000   4.345000 ;
      RECT  0.000000   4.345000  9.455000   4.405000 ;
      RECT  0.000000   4.405000  3.005000  26.495000 ;
      RECT  0.000000   4.460000  9.595000   9.030000 ;
      RECT  0.000000   9.030000 10.725000  10.160000 ;
      RECT  0.000000   9.085000  9.455000   9.155000 ;
      RECT  0.000000   9.155000  9.525000   9.225000 ;
      RECT  0.000000   9.225000  9.595000   9.295000 ;
      RECT  0.000000   9.295000  9.665000   9.365000 ;
      RECT  0.000000   9.365000  9.735000   9.435000 ;
      RECT  0.000000   9.435000  9.805000   9.505000 ;
      RECT  0.000000   9.505000  9.875000   9.575000 ;
      RECT  0.000000   9.575000  9.945000   9.645000 ;
      RECT  0.000000   9.645000 10.015000   9.715000 ;
      RECT  0.000000   9.715000 10.085000   9.785000 ;
      RECT  0.000000   9.785000 10.155000   9.855000 ;
      RECT  0.000000   9.855000 10.225000   9.925000 ;
      RECT  0.000000   9.925000 10.295000   9.995000 ;
      RECT  0.000000   9.995000 10.365000  10.065000 ;
      RECT  0.000000  10.065000 10.435000  10.135000 ;
      RECT  0.000000  10.135000 10.505000  10.205000 ;
      RECT  0.000000  10.160000 10.725000  26.550000 ;
      RECT  0.000000  10.205000 10.575000  10.215000 ;
      RECT  0.000000  26.495000 10.515000  26.565000 ;
      RECT  0.000000  26.550000 10.510000  26.765000 ;
      RECT  0.000000  26.565000 10.445000  26.635000 ;
      RECT  0.000000  26.635000 10.375000  26.705000 ;
      RECT  0.000000  26.705000 10.370000  26.710000 ;
      RECT  0.000000  26.710000  3.005000 196.995000 ;
      RECT  0.000000  26.765000 10.510000  28.470000 ;
      RECT  0.000000  28.470000 10.725000  28.685000 ;
      RECT  0.000000  28.525000 10.370000  28.595000 ;
      RECT  0.000000  28.595000 10.440000  28.665000 ;
      RECT  0.000000  28.665000 10.510000  28.735000 ;
      RECT  0.000000  28.685000 10.725000  31.255000 ;
      RECT  0.000000  28.735000 10.580000  28.740000 ;
      RECT  0.000000  31.255000 11.120000  31.650000 ;
      RECT  0.000000  31.310000 10.585000  31.380000 ;
      RECT  0.000000  31.380000 10.655000  31.450000 ;
      RECT  0.000000  31.450000 10.725000  31.520000 ;
      RECT  0.000000  31.520000 10.795000  31.590000 ;
      RECT  0.000000  31.590000 10.865000  31.660000 ;
      RECT  0.000000  31.650000 11.120000  36.420000 ;
      RECT  0.000000  31.660000 10.935000  31.705000 ;
      RECT  0.000000  36.420000 75.000000 200.000000 ;
      RECT  0.000000 196.995000 75.000000 200.000000 ;
      RECT  3.000000   3.002000  5.145000   4.460000 ;
      RECT  3.000000   4.460000  6.455000  10.330000 ;
      RECT  3.000000  10.330000  6.455000  10.400000 ;
      RECT  3.000000  10.330000  6.455000  10.400000 ;
      RECT  3.000000  10.400000  6.520000  10.470000 ;
      RECT  3.000000  10.400000  6.520000  10.470000 ;
      RECT  3.000000  10.470000  6.595000  10.540000 ;
      RECT  3.000000  10.470000  6.595000  10.540000 ;
      RECT  3.000000  10.540000  6.665000  10.610000 ;
      RECT  3.000000  10.540000  6.665000  10.610000 ;
      RECT  3.000000  10.610000  6.730000  10.680000 ;
      RECT  3.000000  10.610000  6.730000  10.680000 ;
      RECT  3.000000  10.680000  6.805000  10.750000 ;
      RECT  3.000000  10.680000  6.805000  10.750000 ;
      RECT  3.000000  10.750000  6.875000  10.820000 ;
      RECT  3.000000  10.750000  6.875000  10.820000 ;
      RECT  3.000000  10.820000  6.940000  10.890000 ;
      RECT  3.000000  10.820000  6.940000  10.890000 ;
      RECT  3.000000  10.890000  7.015000  10.960000 ;
      RECT  3.000000  10.890000  7.015000  10.960000 ;
      RECT  3.000000  10.960000  7.085000  11.030000 ;
      RECT  3.000000  10.960000  7.085000  11.030000 ;
      RECT  3.000000  11.030000  7.150000  11.100000 ;
      RECT  3.000000  11.030000  7.150000  11.100000 ;
      RECT  3.000000  11.100000  7.225000  11.170000 ;
      RECT  3.000000  11.100000  7.225000  11.170000 ;
      RECT  3.000000  11.170000  7.295000  11.240000 ;
      RECT  3.000000  11.170000  7.295000  11.240000 ;
      RECT  3.000000  11.240000  7.365000  11.310000 ;
      RECT  3.000000  11.240000  7.365000  11.310000 ;
      RECT  3.000000  11.310000  7.435000  11.380000 ;
      RECT  3.000000  11.310000  7.435000  11.380000 ;
      RECT  3.000000  11.380000  7.505000  11.450000 ;
      RECT  3.000000  11.380000  7.505000  11.450000 ;
      RECT  3.000000  11.450000  7.575000  11.460000 ;
      RECT  3.000000  11.450000  7.575000  11.460000 ;
      RECT  3.000000  11.460000  7.585000  25.250000 ;
      RECT  3.000000  25.250000  7.515000  25.320000 ;
      RECT  3.000000  25.250000  7.515000  25.320000 ;
      RECT  3.000000  25.320000  7.440000  25.390000 ;
      RECT  3.000000  25.320000  7.440000  25.390000 ;
      RECT  3.000000  25.390000  7.375000  25.460000 ;
      RECT  3.000000  25.390000  7.375000  25.460000 ;
      RECT  3.000000  25.460000  7.370000  25.465000 ;
      RECT  3.000000  25.460000  7.370000  25.465000 ;
      RECT  3.000000  25.465000  7.370000  29.770000 ;
      RECT  3.000000  29.770000  7.370000  29.840000 ;
      RECT  3.000000  29.770000  7.370000  29.840000 ;
      RECT  3.000000  29.840000  7.435000  29.910000 ;
      RECT  3.000000  29.840000  7.435000  29.910000 ;
      RECT  3.000000  29.910000  7.510000  29.980000 ;
      RECT  3.000000  29.910000  7.510000  29.980000 ;
      RECT  3.000000  29.980000  7.580000  29.985000 ;
      RECT  3.000000  29.980000  7.580000  29.985000 ;
      RECT  3.000000  29.985000  7.585000  32.555000 ;
      RECT  3.000000  32.555000  7.585000  32.625000 ;
      RECT  3.000000  32.555000  7.585000  32.625000 ;
      RECT  3.000000  32.625000  7.650000  32.695000 ;
      RECT  3.000000  32.625000  7.650000  32.695000 ;
      RECT  3.000000  32.695000  7.725000  32.765000 ;
      RECT  3.000000  32.695000  7.725000  32.765000 ;
      RECT  3.000000  32.765000  7.795000  32.835000 ;
      RECT  3.000000  32.765000  7.795000  32.835000 ;
      RECT  3.000000  32.835000  7.865000  32.905000 ;
      RECT  3.000000  32.835000  7.865000  32.905000 ;
      RECT  3.000000  32.905000  7.935000  32.950000 ;
      RECT  3.000000  32.905000  7.935000  32.950000 ;
      RECT  3.000000  32.950000  7.975000  39.560000 ;
      RECT  3.000000  39.560000 72.000000 197.000000 ;
      RECT  5.145000   4.405000  9.455000   7.410000 ;
      RECT  6.450000   1.750000 16.965000   3.155000 ;
      RECT  6.450000   3.155000  9.455000   4.405000 ;
      RECT  6.450000   7.410000  9.455000  10.215000 ;
      RECT  6.455000  10.215000 10.585000  13.220000 ;
      RECT  7.365000  26.710000 10.370000  28.740000 ;
      RECT  7.365000  28.740000 10.585000  31.310000 ;
      RECT  7.370000  23.490000 10.585000  26.495000 ;
      RECT  7.370000  31.310000 10.585000  31.705000 ;
      RECT  7.370000  31.705000 10.980000  31.745000 ;
      RECT  7.580000  13.220000 10.585000  23.490000 ;
      RECT  7.580000  31.745000 10.980000  36.560000 ;
      RECT  7.975000  36.560000 15.435000  39.560000 ;
      RECT  7.975000  39.560000 15.430000  39.565000 ;
      RECT  8.145000   1.460000 12.005000   1.750000 ;
      RECT  9.035000   0.000000 12.145000   1.320000 ;
      RECT  9.175000   0.000000 12.005000   1.460000 ;
      RECT 10.135000   4.685000 15.825000   4.945000 ;
      RECT 10.135000   4.945000 29.180000   5.525000 ;
      RECT 10.135000   5.525000 29.180000   8.800000 ;
      RECT 10.135000   8.800000 29.180000   9.930000 ;
      RECT 10.275000   4.745000 15.430000   4.815000 ;
      RECT 10.275000   4.815000 15.500000   4.885000 ;
      RECT 10.275000   4.885000 15.570000   4.955000 ;
      RECT 10.275000   4.955000 15.640000   5.025000 ;
      RECT 10.275000   5.025000 15.710000   5.085000 ;
      RECT 10.275000   5.085000 28.540000   5.155000 ;
      RECT 10.275000   5.155000 28.610000   5.225000 ;
      RECT 10.275000   5.225000 28.680000   5.295000 ;
      RECT 10.275000   5.295000 28.750000   5.365000 ;
      RECT 10.275000   5.365000 28.820000   5.435000 ;
      RECT 10.275000   5.435000 28.890000   5.505000 ;
      RECT 10.275000   5.505000 28.960000   5.575000 ;
      RECT 10.275000   5.575000 29.030000   5.585000 ;
      RECT 10.275000   5.585000 29.040000   8.590000 ;
      RECT 10.275000   8.590000 14.405000   8.745000 ;
      RECT 10.345000   4.675000 15.360000   4.745000 ;
      RECT 10.345000   8.745000 29.040000   8.815000 ;
      RECT 10.415000   4.605000 15.290000   4.675000 ;
      RECT 10.415000   8.815000 29.040000   8.885000 ;
      RECT 10.485000   4.535000 15.220000   4.605000 ;
      RECT 10.485000   8.885000 29.040000   8.955000 ;
      RECT 10.555000   4.465000 15.150000   4.535000 ;
      RECT 10.555000   8.955000 29.040000   9.025000 ;
      RECT 10.625000   4.395000 15.080000   4.465000 ;
      RECT 10.625000   9.025000 29.040000   9.095000 ;
      RECT 10.695000   4.325000 15.010000   4.395000 ;
      RECT 10.695000   9.095000 29.040000   9.165000 ;
      RECT 10.765000   4.255000 14.940000   4.325000 ;
      RECT 10.765000   9.165000 29.040000   9.235000 ;
      RECT 10.835000   4.185000 14.870000   4.255000 ;
      RECT 10.835000   9.235000 29.040000   9.305000 ;
      RECT 10.905000   4.115000 14.800000   4.185000 ;
      RECT 10.905000   9.305000 29.040000   9.375000 ;
      RECT 10.975000   4.045000 14.730000   4.115000 ;
      RECT 10.975000   9.375000 29.040000   9.445000 ;
      RECT 10.990000   3.835000 15.570000   4.685000 ;
      RECT 11.045000   3.975000 14.660000   4.045000 ;
      RECT 11.045000   9.445000 29.040000   9.515000 ;
      RECT 11.050000  27.360000 75.000000  27.875000 ;
      RECT 11.050000  27.875000 75.000000  28.090000 ;
      RECT 11.115000   9.515000 29.040000   9.585000 ;
      RECT 11.185000   9.585000 29.040000   9.655000 ;
      RECT 11.190000  27.415000 14.805000  27.820000 ;
      RECT 11.195000  27.410000 75.000000  27.415000 ;
      RECT 11.255000   9.655000 29.040000   9.725000 ;
      RECT 11.260000  27.820000 75.000000  27.890000 ;
      RECT 11.265000   9.930000 29.180000  11.145000 ;
      RECT 11.265000  11.145000 29.630000  11.595000 ;
      RECT 11.265000  11.595000 29.630000  15.815000 ;
      RECT 11.265000  15.815000 30.225000  16.410000 ;
      RECT 11.265000  16.410000 30.225000  20.635000 ;
      RECT 11.265000  20.635000 75.000000  27.145000 ;
      RECT 11.265000  27.145000 75.000000  27.360000 ;
      RECT 11.265000  27.340000 75.000000  27.410000 ;
      RECT 11.265000  28.090000 75.000000  31.025000 ;
      RECT 11.265000  31.025000 75.000000  31.420000 ;
      RECT 11.325000   9.725000 29.040000   9.795000 ;
      RECT 11.330000  27.890000 75.000000  27.960000 ;
      RECT 11.335000  27.270000 75.000000  27.340000 ;
      RECT 11.395000   9.795000 29.040000   9.865000 ;
      RECT 11.400000  27.960000 75.000000  28.030000 ;
      RECT 11.405000   9.865000 29.040000   9.875000 ;
      RECT 11.405000   9.875000 14.405000  11.200000 ;
      RECT 11.405000  11.200000 29.040000  11.270000 ;
      RECT 11.405000  11.270000 29.110000  11.340000 ;
      RECT 11.405000  11.340000 29.180000  11.410000 ;
      RECT 11.405000  11.410000 29.250000  11.480000 ;
      RECT 11.405000  11.480000 29.320000  11.550000 ;
      RECT 11.405000  11.550000 29.390000  11.620000 ;
      RECT 11.405000  11.620000 29.460000  11.650000 ;
      RECT 11.405000  11.650000 14.410000  15.870000 ;
      RECT 11.405000  15.870000 29.490000  15.940000 ;
      RECT 11.405000  15.940000 29.560000  16.010000 ;
      RECT 11.405000  16.010000 29.630000  16.080000 ;
      RECT 11.405000  16.080000 29.700000  16.150000 ;
      RECT 11.405000  16.150000 29.770000  16.220000 ;
      RECT 11.405000  16.220000 29.840000  16.290000 ;
      RECT 11.405000  16.290000 29.910000  16.360000 ;
      RECT 11.405000  16.360000 29.980000  16.430000 ;
      RECT 11.405000  16.430000 30.050000  16.465000 ;
      RECT 11.405000  16.465000 14.410000  20.775000 ;
      RECT 11.405000  20.775000 14.805000  27.415000 ;
      RECT 11.405000  27.200000 75.000000  27.270000 ;
      RECT 11.405000  27.820000 14.805000  30.970000 ;
      RECT 11.405000  28.030000 75.000000  28.035000 ;
      RECT 11.475000  30.970000 75.000000  31.040000 ;
      RECT 11.545000  31.040000 75.000000  31.110000 ;
      RECT 11.615000  31.110000 75.000000  31.180000 ;
      RECT 11.660000  31.420000 75.000000  35.880000 ;
      RECT 11.685000  31.180000 75.000000  31.250000 ;
      RECT 11.755000  31.250000 75.000000  31.320000 ;
      RECT 11.800000  30.970000 14.805000  35.740000 ;
      RECT 11.800000  31.320000 75.000000  31.365000 ;
      RECT 12.290000  35.880000 75.000000  36.420000 ;
      RECT 12.430000  20.775000 75.000000  36.560000 ;
      RECT 12.685000   0.000000 14.415000   1.125000 ;
      RECT 12.685000   1.125000 17.105000   1.610000 ;
      RECT 12.795000   1.745000 16.965000   1.750000 ;
      RECT 12.810000   1.730000 16.965000   1.745000 ;
      RECT 12.825000   0.000000 14.275000   1.265000 ;
      RECT 12.825000   1.265000 16.965000   1.715000 ;
      RECT 12.825000   1.715000 16.965000   1.730000 ;
      RECT 13.275000   6.975000 13.415000   7.045000 ;
      RECT 13.275000   6.975000 13.415000   7.045000 ;
      RECT 13.275000   7.045000 13.485000   7.115000 ;
      RECT 13.275000   7.045000 13.485000   7.115000 ;
      RECT 13.275000   7.115000 13.555000   7.185000 ;
      RECT 13.275000   7.115000 13.555000   7.185000 ;
      RECT 13.275000   7.185000 13.625000   7.255000 ;
      RECT 13.275000   7.185000 13.625000   7.255000 ;
      RECT 13.275000   7.255000 13.695000   7.325000 ;
      RECT 13.275000   7.255000 13.695000   7.325000 ;
      RECT 13.275000   7.325000 13.765000   7.395000 ;
      RECT 13.275000   7.325000 13.765000   7.395000 ;
      RECT 13.275000   7.395000 13.835000   7.465000 ;
      RECT 13.275000   7.395000 13.835000   7.465000 ;
      RECT 13.275000   7.465000 13.905000   7.500000 ;
      RECT 13.275000   7.465000 13.905000   7.500000 ;
      RECT 13.345000   7.500000 13.940000   7.570000 ;
      RECT 13.345000   7.500000 13.940000   7.570000 ;
      RECT 13.415000   7.570000 14.010000   7.640000 ;
      RECT 13.415000   7.570000 14.010000   7.640000 ;
      RECT 13.485000   7.640000 14.080000   7.710000 ;
      RECT 13.485000   7.640000 14.080000   7.710000 ;
      RECT 13.555000   7.710000 14.150000   7.780000 ;
      RECT 13.555000   7.710000 14.150000   7.780000 ;
      RECT 13.625000   7.780000 14.220000   7.850000 ;
      RECT 13.625000   7.780000 14.220000   7.850000 ;
      RECT 13.695000   7.850000 14.290000   7.920000 ;
      RECT 13.695000   7.850000 14.290000   7.920000 ;
      RECT 13.765000   7.920000 14.360000   7.990000 ;
      RECT 13.765000   7.920000 14.360000   7.990000 ;
      RECT 13.835000   7.990000 14.430000   8.060000 ;
      RECT 13.835000   7.990000 14.430000   8.060000 ;
      RECT 13.860000   8.060000 14.500000   8.085000 ;
      RECT 13.860000   8.060000 14.500000   8.085000 ;
      RECT 13.930000   8.085000 26.040000   8.155000 ;
      RECT 13.930000   8.085000 26.040000   8.155000 ;
      RECT 14.000000   8.155000 26.040000   8.225000 ;
      RECT 14.000000   8.155000 26.040000   8.225000 ;
      RECT 14.070000   8.225000 26.040000   8.295000 ;
      RECT 14.070000   8.225000 26.040000   8.295000 ;
      RECT 14.140000   8.295000 26.040000   8.365000 ;
      RECT 14.140000   8.295000 26.040000   8.365000 ;
      RECT 14.210000   8.365000 26.040000   8.435000 ;
      RECT 14.210000   8.365000 26.040000   8.435000 ;
      RECT 14.280000   8.435000 26.040000   8.505000 ;
      RECT 14.280000   8.435000 26.040000   8.505000 ;
      RECT 14.350000   8.505000 26.040000   8.575000 ;
      RECT 14.350000   8.505000 26.040000   8.575000 ;
      RECT 14.405000   8.575000 26.040000   8.630000 ;
      RECT 14.405000   8.575000 26.040000   8.630000 ;
      RECT 14.405000   8.630000 26.040000  12.445000 ;
      RECT 14.405000  12.445000 26.040000  12.515000 ;
      RECT 14.405000  12.445000 26.040000  12.515000 ;
      RECT 14.405000  12.515000 26.110000  12.585000 ;
      RECT 14.405000  12.515000 26.110000  12.585000 ;
      RECT 14.405000  12.585000 26.180000  12.655000 ;
      RECT 14.405000  12.585000 26.180000  12.655000 ;
      RECT 14.405000  12.655000 26.250000  12.725000 ;
      RECT 14.405000  12.655000 26.250000  12.725000 ;
      RECT 14.405000  12.725000 26.320000  12.795000 ;
      RECT 14.405000  12.725000 26.320000  12.795000 ;
      RECT 14.405000  12.795000 26.390000  12.865000 ;
      RECT 14.405000  12.795000 26.390000  12.865000 ;
      RECT 14.405000  12.865000 26.455000  12.895000 ;
      RECT 14.405000  12.865000 26.455000  12.895000 ;
      RECT 14.405000  12.895000 26.490000  17.115000 ;
      RECT 14.405000  17.115000 26.490000  17.185000 ;
      RECT 14.405000  17.115000 26.490000  17.185000 ;
      RECT 14.405000  17.185000 26.560000  17.255000 ;
      RECT 14.405000  17.185000 26.560000  17.255000 ;
      RECT 14.405000  17.255000 26.630000  17.325000 ;
      RECT 14.405000  17.255000 26.630000  17.325000 ;
      RECT 14.405000  17.325000 26.700000  17.395000 ;
      RECT 14.405000  17.325000 26.700000  17.395000 ;
      RECT 14.405000  17.395000 26.770000  17.465000 ;
      RECT 14.405000  17.395000 26.770000  17.465000 ;
      RECT 14.405000  17.465000 26.840000  17.535000 ;
      RECT 14.405000  17.465000 26.840000  17.535000 ;
      RECT 14.405000  17.535000 26.910000  17.605000 ;
      RECT 14.405000  17.535000 26.910000  17.605000 ;
      RECT 14.405000  17.605000 26.980000  17.675000 ;
      RECT 14.405000  17.605000 26.980000  17.675000 ;
      RECT 14.405000  17.675000 27.045000  17.710000 ;
      RECT 14.405000  17.675000 27.045000  17.710000 ;
      RECT 14.405000  17.710000 27.080000  23.775000 ;
      RECT 14.405000  23.775000 72.000000  29.725000 ;
      RECT 14.475000  29.725000 72.000000  29.795000 ;
      RECT 14.475000  29.725000 72.000000  29.795000 ;
      RECT 14.545000  29.795000 72.000000  29.865000 ;
      RECT 14.545000  29.795000 72.000000  29.865000 ;
      RECT 14.615000  29.865000 72.000000  29.935000 ;
      RECT 14.615000  29.865000 72.000000  29.935000 ;
      RECT 14.685000  29.935000 72.000000  30.005000 ;
      RECT 14.685000  29.935000 72.000000  30.005000 ;
      RECT 14.755000  30.005000 72.000000  30.075000 ;
      RECT 14.755000  30.005000 72.000000  30.075000 ;
      RECT 14.800000  30.075000 72.000000  30.120000 ;
      RECT 14.800000  30.075000 72.000000  30.120000 ;
      RECT 14.800000  30.120000 72.000000  32.740000 ;
      RECT 14.945000   3.295000 19.935000   3.595000 ;
      RECT 15.070000   3.155000 16.965000   3.225000 ;
      RECT 15.140000   3.225000 16.965000   3.295000 ;
      RECT 15.210000   3.295000 16.965000   3.365000 ;
      RECT 15.245000   3.595000 22.220000   4.185000 ;
      RECT 15.260000   3.365000 16.965000   3.415000 ;
      RECT 15.275000   0.000000 17.105000   1.125000 ;
      RECT 15.330000   3.415000 19.795000   3.485000 ;
      RECT 15.400000   3.485000 19.795000   3.555000 ;
      RECT 15.415000   0.000000 16.965000   1.265000 ;
      RECT 15.430000  32.740000 72.000000  39.560000 ;
      RECT 15.470000   3.555000 19.795000   3.625000 ;
      RECT 15.540000   3.625000 19.795000   3.695000 ;
      RECT 15.580000   3.695000 19.795000   3.735000 ;
      RECT 15.650000   3.735000 22.080000   3.805000 ;
      RECT 15.720000   3.805000 22.080000   3.875000 ;
      RECT 15.790000   3.875000 22.080000   3.945000 ;
      RECT 15.835000   4.185000 22.000000   4.405000 ;
      RECT 15.860000   3.945000 22.080000   4.015000 ;
      RECT 15.930000   4.015000 22.080000   4.085000 ;
      RECT 15.975000   4.085000 22.080000   4.130000 ;
      RECT 16.040000   4.130000 22.015000   4.195000 ;
      RECT 16.110000   4.195000 21.945000   4.265000 ;
      RECT 19.050000   0.000000 19.935000   3.275000 ;
      RECT 19.190000   0.000000 19.795000   3.415000 ;
      RECT 21.365000   0.000000 22.220000   3.595000 ;
      RECT 21.505000   0.000000 22.080000   3.735000 ;
      RECT 22.800000   0.000000 27.440000   0.470000 ;
      RECT 22.800000   0.470000 28.775000   0.475000 ;
      RECT 22.800000   0.475000 32.620000   0.780000 ;
      RECT 22.800000   0.780000 72.075000   0.910000 ;
      RECT 22.800000   0.910000 75.000000   4.200000 ;
      RECT 22.800000   4.200000 75.000000   4.405000 ;
      RECT 22.940000   0.000000 27.300000   0.610000 ;
      RECT 22.940000   0.610000 28.635000   0.615000 ;
      RECT 22.940000   0.615000 32.480000   0.920000 ;
      RECT 22.940000   0.920000 33.300000   3.925000 ;
      RECT 22.940000   3.925000 29.860000   4.145000 ;
      RECT 23.000000   4.145000 75.000000   4.205000 ;
      RECT 23.060000   4.205000 75.000000   4.265000 ;
      RECT 26.035000   8.590000 29.040000   8.745000 ;
      RECT 26.040000   9.875000 29.040000  11.200000 ;
      RECT 26.040000  11.650000 29.490000  14.655000 ;
      RECT 26.485000  14.655000 29.490000  15.870000 ;
      RECT 26.490000  16.465000 30.085000  19.470000 ;
      RECT 27.080000  19.470000 30.085000  20.775000 ;
      RECT 28.370000   0.000000 28.775000   0.470000 ;
      RECT 28.825000   4.405000 75.000000   5.300000 ;
      RECT 28.950000   4.265000 75.000000   4.335000 ;
      RECT 29.020000   4.335000 75.000000   4.405000 ;
      RECT 29.090000   4.405000 75.000000   4.475000 ;
      RECT 29.160000   4.475000 75.000000   4.545000 ;
      RECT 29.230000   4.545000 75.000000   4.615000 ;
      RECT 29.300000   4.615000 75.000000   4.685000 ;
      RECT 29.370000   4.685000 75.000000   4.755000 ;
      RECT 29.440000   4.755000 75.000000   4.825000 ;
      RECT 29.510000   4.825000 75.000000   4.895000 ;
      RECT 29.580000   4.895000 75.000000   4.965000 ;
      RECT 29.650000   4.965000 75.000000   5.035000 ;
      RECT 29.720000   5.035000 75.000000   5.105000 ;
      RECT 29.720000   5.300000 75.000000  10.915000 ;
      RECT 29.720000  10.915000 75.000000  11.365000 ;
      RECT 29.790000   5.105000 75.000000   5.175000 ;
      RECT 29.825000   0.000000 30.365000   0.470000 ;
      RECT 29.825000   0.470000 32.620000   0.475000 ;
      RECT 29.860000   1.050000 75.000000  10.860000 ;
      RECT 29.860000   1.050000 75.000000  10.860000 ;
      RECT 29.860000   5.175000 75.000000   5.245000 ;
      RECT 29.930000  10.860000 75.000000  10.930000 ;
      RECT 29.965000   0.000000 30.225000   0.610000 ;
      RECT 29.965000   0.610000 32.480000   0.615000 ;
      RECT 30.000000  10.930000 75.000000  11.000000 ;
      RECT 30.070000  11.000000 75.000000  11.070000 ;
      RECT 30.140000  11.070000 75.000000  11.140000 ;
      RECT 30.170000  11.365000 75.000000  15.585000 ;
      RECT 30.170000  15.585000 75.000000  16.180000 ;
      RECT 30.210000  11.140000 75.000000  11.210000 ;
      RECT 30.280000  11.210000 75.000000  11.280000 ;
      RECT 30.310000  10.860000 33.315000  12.525000 ;
      RECT 30.310000  11.280000 75.000000  11.310000 ;
      RECT 30.310000  12.525000 33.905000  15.530000 ;
      RECT 30.380000  15.530000 75.000000  15.600000 ;
      RECT 30.450000  15.600000 75.000000  15.670000 ;
      RECT 30.520000  15.670000 75.000000  15.740000 ;
      RECT 30.590000  15.740000 75.000000  15.810000 ;
      RECT 30.660000  15.810000 75.000000  15.880000 ;
      RECT 30.730000  15.880000 75.000000  15.950000 ;
      RECT 30.765000  16.180000 75.000000  20.635000 ;
      RECT 30.800000  15.950000 75.000000  16.020000 ;
      RECT 30.870000  16.020000 75.000000  16.090000 ;
      RECT 30.905000  16.090000 75.000000  16.125000 ;
      RECT 30.905000  16.125000 33.910000  20.775000 ;
      RECT 31.295000   0.000000 32.620000   0.470000 ;
      RECT 31.435000   0.000000 32.480000   0.610000 ;
      RECT 32.820000   3.920000 68.935000   3.960000 ;
      RECT 32.820000   3.920000 68.935000   3.960000 ;
      RECT 32.860000   3.960000 68.935000   4.000000 ;
      RECT 32.860000   3.960000 68.935000   4.000000 ;
      RECT 32.860000   4.000000 68.935000   4.050000 ;
      RECT 32.860000   4.050000 72.000000   9.615000 ;
      RECT 32.930000   9.615000 72.000000   9.685000 ;
      RECT 32.930000   9.615000 72.000000   9.685000 ;
      RECT 33.000000   9.685000 72.000000   9.755000 ;
      RECT 33.000000   9.685000 72.000000   9.755000 ;
      RECT 33.070000   9.755000 72.000000   9.825000 ;
      RECT 33.070000   9.755000 72.000000   9.825000 ;
      RECT 33.140000   9.825000 72.000000   9.895000 ;
      RECT 33.140000   9.825000 72.000000   9.895000 ;
      RECT 33.160000   0.000000 72.075000   0.780000 ;
      RECT 33.210000   9.895000 72.000000   9.965000 ;
      RECT 33.210000   9.895000 72.000000   9.965000 ;
      RECT 33.280000   9.965000 72.000000  10.035000 ;
      RECT 33.280000   9.965000 72.000000  10.035000 ;
      RECT 33.300000   0.000000 71.935000  10.860000 ;
      RECT 33.300000   0.000000 71.935000  10.860000 ;
      RECT 33.310000  10.035000 72.000000  10.065000 ;
      RECT 33.310000  10.035000 72.000000  10.065000 ;
      RECT 33.310000  10.065000 72.000000  14.285000 ;
      RECT 33.380000  14.285000 72.000000  14.355000 ;
      RECT 33.380000  14.285000 72.000000  14.355000 ;
      RECT 33.450000  14.355000 72.000000  14.425000 ;
      RECT 33.450000  14.355000 72.000000  14.425000 ;
      RECT 33.520000  14.425000 72.000000  14.495000 ;
      RECT 33.520000  14.425000 72.000000  14.495000 ;
      RECT 33.590000  14.495000 72.000000  14.565000 ;
      RECT 33.590000  14.495000 72.000000  14.565000 ;
      RECT 33.660000  14.565000 72.000000  14.635000 ;
      RECT 33.660000  14.565000 72.000000  14.635000 ;
      RECT 33.730000  14.635000 72.000000  14.705000 ;
      RECT 33.730000  14.635000 72.000000  14.705000 ;
      RECT 33.800000  14.705000 72.000000  14.775000 ;
      RECT 33.800000  14.705000 72.000000  14.775000 ;
      RECT 33.870000  14.775000 72.000000  14.845000 ;
      RECT 33.870000  14.775000 72.000000  14.845000 ;
      RECT 33.905000  14.845000 72.000000  14.880000 ;
      RECT 33.905000  14.845000 72.000000  14.880000 ;
      RECT 33.905000  14.880000 72.000000  23.775000 ;
      RECT 36.300000   3.000000 68.935000   3.920000 ;
      RECT 71.995000  10.860000 75.000000  15.530000 ;
      RECT 71.995000  16.125000 75.000000  20.775000 ;
      RECT 71.995000  36.560000 75.000000 196.995000 ;
      RECT 73.130000   1.020000 75.000000   1.050000 ;
      RECT 73.375000   0.000000 75.000000   0.910000 ;
      RECT 73.515000   0.000000 75.000000   1.020000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  8.000000   3.005000 ;
      RECT  0.000000   0.000000  8.100000  15.660000 ;
      RECT  0.000000   3.005000  3.005000  17.245000 ;
      RECT  0.000000  15.620000  7.850000  15.770000 ;
      RECT  0.000000  15.660000  6.475000  17.285000 ;
      RECT  0.000000  15.770000  7.700000  15.920000 ;
      RECT  0.000000  15.920000  7.550000  16.070000 ;
      RECT  0.000000  16.070000  7.400000  16.220000 ;
      RECT  0.000000  16.220000  7.250000  16.370000 ;
      RECT  0.000000  16.370000  7.100000  16.520000 ;
      RECT  0.000000  16.520000  6.950000  16.670000 ;
      RECT  0.000000  16.670000  6.800000  16.820000 ;
      RECT  0.000000  16.820000  6.650000  16.970000 ;
      RECT  0.000000  16.970000  6.500000  17.120000 ;
      RECT  0.000000  17.120000  6.375000  17.245000 ;
      RECT  0.000000  17.245000  6.375000  64.435000 ;
      RECT  0.000000  17.285000  6.475000  31.630000 ;
      RECT  0.000000  31.630000  9.270000  34.425000 ;
      RECT  0.000000  31.670000  6.375000  31.820000 ;
      RECT  0.000000  31.820000  6.525000  31.970000 ;
      RECT  0.000000  31.970000  6.675000  32.120000 ;
      RECT  0.000000  32.120000  6.825000  32.270000 ;
      RECT  0.000000  32.270000  6.975000  32.420000 ;
      RECT  0.000000  32.420000  7.125000  32.570000 ;
      RECT  0.000000  32.570000  7.275000  32.720000 ;
      RECT  0.000000  32.720000  7.425000  32.870000 ;
      RECT  0.000000  32.870000  7.575000  33.020000 ;
      RECT  0.000000  33.020000  7.725000  33.170000 ;
      RECT  0.000000  33.170000  7.875000  33.320000 ;
      RECT  0.000000  33.320000  8.025000  33.470000 ;
      RECT  0.000000  33.470000  8.175000  33.620000 ;
      RECT  0.000000  33.620000  8.325000  33.770000 ;
      RECT  0.000000  33.770000  8.475000  33.920000 ;
      RECT  0.000000  33.920000  8.625000  34.070000 ;
      RECT  0.000000  34.070000  8.775000  34.220000 ;
      RECT  0.000000  34.220000  8.925000  34.370000 ;
      RECT  0.000000  34.370000  9.075000  34.520000 ;
      RECT  0.000000  34.425000 71.890000  64.475000 ;
      RECT  0.000000  34.520000  9.225000  34.525000 ;
      RECT  0.000000  64.435000 71.640000  64.585000 ;
      RECT  0.000000  64.475000 64.560000  71.805000 ;
      RECT  0.000000  64.585000 71.490000  64.735000 ;
      RECT  0.000000  64.735000 71.340000  64.885000 ;
      RECT  0.000000  64.885000 71.190000  65.035000 ;
      RECT  0.000000  65.035000 71.040000  65.185000 ;
      RECT  0.000000  65.185000 70.890000  65.335000 ;
      RECT  0.000000  65.335000 70.740000  65.485000 ;
      RECT  0.000000  65.485000 70.590000  65.635000 ;
      RECT  0.000000  65.635000 70.440000  65.785000 ;
      RECT  0.000000  65.785000 70.290000  65.935000 ;
      RECT  0.000000  65.935000 70.140000  66.085000 ;
      RECT  0.000000  66.085000 69.990000  66.235000 ;
      RECT  0.000000  66.235000 69.840000  66.385000 ;
      RECT  0.000000  66.385000 69.690000  66.535000 ;
      RECT  0.000000  66.535000 69.540000  66.685000 ;
      RECT  0.000000  66.685000 69.390000  66.835000 ;
      RECT  0.000000  66.835000 69.240000  66.985000 ;
      RECT  0.000000  66.985000 69.090000  67.135000 ;
      RECT  0.000000  67.135000 68.940000  67.285000 ;
      RECT  0.000000  67.285000 68.790000  67.435000 ;
      RECT  0.000000  67.435000 68.640000  67.585000 ;
      RECT  0.000000  67.585000 68.490000  67.735000 ;
      RECT  0.000000  67.735000 68.340000  67.885000 ;
      RECT  0.000000  67.885000 68.190000  68.035000 ;
      RECT  0.000000  68.035000 68.040000  68.185000 ;
      RECT  0.000000  68.185000 67.890000  68.335000 ;
      RECT  0.000000  68.335000 67.740000  68.485000 ;
      RECT  0.000000  68.485000 67.590000  68.635000 ;
      RECT  0.000000  68.635000 67.440000  68.785000 ;
      RECT  0.000000  68.785000 67.290000  68.935000 ;
      RECT  0.000000  68.935000 67.140000  69.085000 ;
      RECT  0.000000  69.085000 66.990000  69.235000 ;
      RECT  0.000000  69.235000 66.840000  69.385000 ;
      RECT  0.000000  69.385000 66.690000  69.535000 ;
      RECT  0.000000  69.535000 66.540000  69.685000 ;
      RECT  0.000000  69.685000 66.390000  69.835000 ;
      RECT  0.000000  69.835000 66.240000  69.985000 ;
      RECT  0.000000  69.985000 66.090000  70.135000 ;
      RECT  0.000000  70.135000 65.940000  70.285000 ;
      RECT  0.000000  70.285000 65.790000  70.435000 ;
      RECT  0.000000  70.435000 65.640000  70.585000 ;
      RECT  0.000000  70.585000 65.490000  70.735000 ;
      RECT  0.000000  70.735000 65.340000  70.885000 ;
      RECT  0.000000  70.885000 65.190000  71.035000 ;
      RECT  0.000000  71.035000 65.040000  71.185000 ;
      RECT  0.000000  71.185000 64.890000  71.335000 ;
      RECT  0.000000  71.335000 64.740000  71.485000 ;
      RECT  0.000000  71.485000 64.590000  71.635000 ;
      RECT  0.000000  71.635000 64.460000  71.765000 ;
      RECT  0.000000  71.765000  3.005000 196.995000 ;
      RECT  0.000000  71.805000 64.560000  94.945000 ;
      RECT  0.000000  94.945000 75.000000 200.000000 ;
      RECT  0.000000 196.995000 75.000000 200.000000 ;
      RECT  3.000000   3.002000  5.000000  14.375000 ;
      RECT  3.000000  14.375000  4.850000  14.525000 ;
      RECT  3.000000  14.375000  4.850000  14.525000 ;
      RECT  3.000000  14.525000  4.700000  14.675000 ;
      RECT  3.000000  14.525000  4.700000  14.675000 ;
      RECT  3.000000  14.675000  4.550000  14.825000 ;
      RECT  3.000000  14.675000  4.550000  14.825000 ;
      RECT  3.000000  14.825000  4.395000  14.975000 ;
      RECT  3.000000  14.825000  4.395000  14.975000 ;
      RECT  3.000000  14.975000  4.250000  15.125000 ;
      RECT  3.000000  14.975000  4.250000  15.125000 ;
      RECT  3.000000  15.125000  4.100000  15.275000 ;
      RECT  3.000000  15.125000  4.100000  15.275000 ;
      RECT  3.000000  15.275000  3.945000  15.425000 ;
      RECT  3.000000  15.275000  3.945000  15.425000 ;
      RECT  3.000000  15.425000  3.800000  15.575000 ;
      RECT  3.000000  15.425000  3.800000  15.575000 ;
      RECT  3.000000  15.575000  3.650000  15.725000 ;
      RECT  3.000000  15.575000  3.650000  15.725000 ;
      RECT  3.000000  15.725000  3.500000  15.875000 ;
      RECT  3.000000  15.725000  3.500000  15.875000 ;
      RECT  3.000000  15.875000  3.375000  16.000000 ;
      RECT  3.000000  15.875000  3.375000  16.000000 ;
      RECT  3.000000  16.000000  3.375000  32.915000 ;
      RECT  3.000000  32.915000  3.375000  33.065000 ;
      RECT  3.000000  32.915000  3.375000  33.065000 ;
      RECT  3.000000  33.065000  3.525000  33.215000 ;
      RECT  3.000000  33.065000  3.525000  33.215000 ;
      RECT  3.000000  33.215000  3.675000  33.365000 ;
      RECT  3.000000  33.215000  3.675000  33.365000 ;
      RECT  3.000000  33.365000  3.820000  33.515000 ;
      RECT  3.000000  33.365000  3.820000  33.515000 ;
      RECT  3.000000  33.515000  3.970000  33.665000 ;
      RECT  3.000000  33.515000  3.970000  33.665000 ;
      RECT  3.000000  33.665000  4.125000  33.815000 ;
      RECT  3.000000  33.665000  4.125000  33.815000 ;
      RECT  3.000000  33.815000  4.270000  33.965000 ;
      RECT  3.000000  33.815000  4.270000  33.965000 ;
      RECT  3.000000  33.965000  4.425000  34.115000 ;
      RECT  3.000000  33.965000  4.425000  34.115000 ;
      RECT  3.000000  34.115000  4.575000  34.265000 ;
      RECT  3.000000  34.115000  4.575000  34.265000 ;
      RECT  3.000000  34.265000  4.725000  34.415000 ;
      RECT  3.000000  34.265000  4.725000  34.415000 ;
      RECT  3.000000  34.415000  4.875000  34.565000 ;
      RECT  3.000000  34.415000  4.875000  34.565000 ;
      RECT  3.000000  34.565000  5.020000  34.715000 ;
      RECT  3.000000  34.565000  5.020000  34.715000 ;
      RECT  3.000000  34.715000  5.175000  34.865000 ;
      RECT  3.000000  34.715000  5.175000  34.865000 ;
      RECT  3.000000  34.865000  5.325000  35.015000 ;
      RECT  3.000000  34.865000  5.325000  35.015000 ;
      RECT  3.000000  35.015000  5.475000  35.165000 ;
      RECT  3.000000  35.015000  5.475000  35.165000 ;
      RECT  3.000000  35.165000  5.625000  35.315000 ;
      RECT  3.000000  35.165000  5.625000  35.315000 ;
      RECT  3.000000  35.315000  5.770000  35.465000 ;
      RECT  3.000000  35.315000  5.770000  35.465000 ;
      RECT  3.000000  35.465000  5.925000  35.615000 ;
      RECT  3.000000  35.465000  5.925000  35.615000 ;
      RECT  3.000000  35.615000  6.075000  35.765000 ;
      RECT  3.000000  35.615000  6.075000  35.765000 ;
      RECT  3.000000  35.765000  6.225000  35.915000 ;
      RECT  3.000000  35.765000  6.225000  35.915000 ;
      RECT  3.000000  35.915000  6.375000  36.065000 ;
      RECT  3.000000  35.915000  6.375000  36.065000 ;
      RECT  3.000000  36.065000  6.520000  36.215000 ;
      RECT  3.000000  36.065000  6.520000  36.215000 ;
      RECT  3.000000  36.215000  6.675000  36.365000 ;
      RECT  3.000000  36.215000  6.675000  36.365000 ;
      RECT  3.000000  36.365000  6.825000  36.515000 ;
      RECT  3.000000  36.365000  6.825000  36.515000 ;
      RECT  3.000000  36.515000  6.975000  36.665000 ;
      RECT  3.000000  36.515000  6.975000  36.665000 ;
      RECT  3.000000  36.665000  7.125000  36.815000 ;
      RECT  3.000000  36.665000  7.125000  36.815000 ;
      RECT  3.000000  36.815000  7.270000  36.965000 ;
      RECT  3.000000  36.815000  7.270000  36.965000 ;
      RECT  3.000000  36.965000  7.425000  37.115000 ;
      RECT  3.000000  36.965000  7.425000  37.115000 ;
      RECT  3.000000  37.115000  7.575000  37.265000 ;
      RECT  3.000000  37.115000  7.575000  37.265000 ;
      RECT  3.000000  37.265000  7.725000  37.415000 ;
      RECT  3.000000  37.265000  7.725000  37.415000 ;
      RECT  3.000000  37.415000  7.875000  37.525000 ;
      RECT  3.000000  37.415000  7.875000  37.525000 ;
      RECT  3.000000  37.525000 68.785000  63.190000 ;
      RECT  3.000000  63.190000 68.640000  63.340000 ;
      RECT  3.000000  63.190000 68.640000  63.340000 ;
      RECT  3.000000  63.340000 68.490000  63.490000 ;
      RECT  3.000000  63.340000 68.490000  63.490000 ;
      RECT  3.000000  63.490000 68.335000  63.640000 ;
      RECT  3.000000  63.490000 68.335000  63.640000 ;
      RECT  3.000000  63.640000 68.190000  63.790000 ;
      RECT  3.000000  63.640000 68.190000  63.790000 ;
      RECT  3.000000  63.790000 68.035000  63.940000 ;
      RECT  3.000000  63.790000 68.035000  63.940000 ;
      RECT  3.000000  63.940000 67.890000  64.090000 ;
      RECT  3.000000  63.940000 67.890000  64.090000 ;
      RECT  3.000000  64.090000 67.740000  64.240000 ;
      RECT  3.000000  64.090000 67.740000  64.240000 ;
      RECT  3.000000  64.240000 67.585000  64.390000 ;
      RECT  3.000000  64.240000 67.585000  64.390000 ;
      RECT  3.000000  64.390000 67.440000  64.540000 ;
      RECT  3.000000  64.390000 67.440000  64.540000 ;
      RECT  3.000000  64.540000 67.285000  64.690000 ;
      RECT  3.000000  64.540000 67.285000  64.690000 ;
      RECT  3.000000  64.690000 67.140000  64.840000 ;
      RECT  3.000000  64.690000 67.140000  64.840000 ;
      RECT  3.000000  64.840000 66.990000  64.990000 ;
      RECT  3.000000  64.840000 66.990000  64.990000 ;
      RECT  3.000000  64.990000 66.835000  65.140000 ;
      RECT  3.000000  64.990000 66.835000  65.140000 ;
      RECT  3.000000  65.140000 66.690000  65.290000 ;
      RECT  3.000000  65.140000 66.690000  65.290000 ;
      RECT  3.000000  65.290000 66.535000  65.440000 ;
      RECT  3.000000  65.290000 66.535000  65.440000 ;
      RECT  3.000000  65.440000 66.390000  65.590000 ;
      RECT  3.000000  65.440000 66.390000  65.590000 ;
      RECT  3.000000  65.590000 66.240000  65.740000 ;
      RECT  3.000000  65.590000 66.240000  65.740000 ;
      RECT  3.000000  65.740000 66.085000  65.890000 ;
      RECT  3.000000  65.740000 66.085000  65.890000 ;
      RECT  3.000000  65.890000 65.940000  66.040000 ;
      RECT  3.000000  65.890000 65.940000  66.040000 ;
      RECT  3.000000  66.040000 65.785000  66.190000 ;
      RECT  3.000000  66.040000 65.785000  66.190000 ;
      RECT  3.000000  66.190000 65.640000  66.340000 ;
      RECT  3.000000  66.190000 65.640000  66.340000 ;
      RECT  3.000000  66.340000 65.485000  66.490000 ;
      RECT  3.000000  66.340000 65.485000  66.490000 ;
      RECT  3.000000  66.490000 65.335000  66.640000 ;
      RECT  3.000000  66.490000 65.335000  66.640000 ;
      RECT  3.000000  66.640000 65.190000  66.790000 ;
      RECT  3.000000  66.640000 65.190000  66.790000 ;
      RECT  3.000000  66.790000 65.035000  66.940000 ;
      RECT  3.000000  66.790000 65.035000  66.940000 ;
      RECT  3.000000  66.940000 64.890000  67.090000 ;
      RECT  3.000000  66.940000 64.890000  67.090000 ;
      RECT  3.000000  67.090000 64.735000  67.240000 ;
      RECT  3.000000  67.090000 64.735000  67.240000 ;
      RECT  3.000000  67.240000 64.585000  67.390000 ;
      RECT  3.000000  67.240000 64.585000  67.390000 ;
      RECT  3.000000  67.390000 64.440000  67.540000 ;
      RECT  3.000000  67.390000 64.440000  67.540000 ;
      RECT  3.000000  67.540000 64.285000  67.690000 ;
      RECT  3.000000  67.540000 64.285000  67.690000 ;
      RECT  3.000000  67.690000 64.140000  67.840000 ;
      RECT  3.000000  67.690000 64.140000  67.840000 ;
      RECT  3.000000  67.840000 63.990000  67.990000 ;
      RECT  3.000000  67.840000 63.990000  67.990000 ;
      RECT  3.000000  67.990000 63.840000  68.140000 ;
      RECT  3.000000  67.990000 63.840000  68.140000 ;
      RECT  3.000000  68.140000 63.690000  68.290000 ;
      RECT  3.000000  68.140000 63.690000  68.290000 ;
      RECT  3.000000  68.290000 63.540000  68.440000 ;
      RECT  3.000000  68.290000 63.540000  68.440000 ;
      RECT  3.000000  68.440000 63.390000  68.590000 ;
      RECT  3.000000  68.440000 63.390000  68.590000 ;
      RECT  3.000000  68.590000 63.240000  68.740000 ;
      RECT  3.000000  68.590000 63.240000  68.740000 ;
      RECT  3.000000  68.740000 63.090000  68.890000 ;
      RECT  3.000000  68.740000 63.090000  68.890000 ;
      RECT  3.000000  68.890000 62.940000  69.040000 ;
      RECT  3.000000  68.890000 62.940000  69.040000 ;
      RECT  3.000000  69.040000 62.790000  69.190000 ;
      RECT  3.000000  69.040000 62.790000  69.190000 ;
      RECT  3.000000  69.190000 62.640000  69.340000 ;
      RECT  3.000000  69.190000 62.640000  69.340000 ;
      RECT  3.000000  69.340000 62.490000  69.490000 ;
      RECT  3.000000  69.340000 62.490000  69.490000 ;
      RECT  3.000000  69.490000 62.340000  69.640000 ;
      RECT  3.000000  69.490000 62.340000  69.640000 ;
      RECT  3.000000  69.640000 62.190000  69.790000 ;
      RECT  3.000000  69.640000 62.190000  69.790000 ;
      RECT  3.000000  69.790000 62.040000  69.940000 ;
      RECT  3.000000  69.790000 62.040000  69.940000 ;
      RECT  3.000000  69.940000 61.890000  70.090000 ;
      RECT  3.000000  69.940000 61.890000  70.090000 ;
      RECT  3.000000  70.090000 61.740000  70.240000 ;
      RECT  3.000000  70.090000 61.740000  70.240000 ;
      RECT  3.000000  70.240000 61.590000  70.390000 ;
      RECT  3.000000  70.240000 61.590000  70.390000 ;
      RECT  3.000000  70.390000 61.460000  70.520000 ;
      RECT  3.000000  70.390000 61.460000  70.520000 ;
      RECT  3.000000  70.520000 61.460000  98.045000 ;
      RECT  3.000000  98.045000 72.000000 197.000000 ;
      RECT  3.370000   3.005000  8.000000  15.620000 ;
      RECT  3.370000  15.620000  6.375000  17.245000 ;
      RECT  6.375000  34.525000 25.680000  37.525000 ;
      RECT  6.375000  37.525000 25.675000  37.530000 ;
      RECT  7.595000  17.745000 71.890000  31.170000 ;
      RECT  7.595000  31.170000 71.890000  33.095000 ;
      RECT  7.695000  17.785000 12.325000  28.125000 ;
      RECT  7.695000  28.125000 25.675000  29.990000 ;
      RECT  7.695000  29.990000 25.680000  31.130000 ;
      RECT  7.820000  17.660000 71.790000  17.785000 ;
      RECT  7.845000  31.130000 71.790000  31.280000 ;
      RECT  7.970000  17.510000 71.790000  17.660000 ;
      RECT  7.995000  31.280000 71.790000  31.430000 ;
      RECT  8.120000  17.360000 71.790000  17.510000 ;
      RECT  8.145000  31.430000 71.790000  31.580000 ;
      RECT  8.270000  17.210000 71.790000  17.360000 ;
      RECT  8.295000  31.580000 71.790000  31.730000 ;
      RECT  8.420000  17.060000 71.790000  17.210000 ;
      RECT  8.445000  31.730000 71.790000  31.880000 ;
      RECT  8.570000  16.910000 71.790000  17.060000 ;
      RECT  8.595000  31.880000 71.790000  32.030000 ;
      RECT  8.720000  16.760000 71.790000  16.910000 ;
      RECT  8.745000  32.030000 71.790000  32.180000 ;
      RECT  8.870000  16.610000 71.790000  16.760000 ;
      RECT  8.895000  32.180000 71.790000  32.330000 ;
      RECT  9.020000  16.460000 71.790000  16.610000 ;
      RECT  9.045000  32.330000 71.790000  32.480000 ;
      RECT  9.170000  16.310000 71.790000  16.460000 ;
      RECT  9.195000  32.480000 71.790000  32.630000 ;
      RECT  9.220000   0.000000 16.945000   3.435000 ;
      RECT  9.220000   3.435000 19.775000   7.275000 ;
      RECT  9.220000   7.275000 22.605000  10.105000 ;
      RECT  9.220000  10.105000 22.605000  12.565000 ;
      RECT  9.220000  12.565000 27.870000  15.070000 ;
      RECT  9.220000  15.070000 71.890000  16.120000 ;
      RECT  9.220000  16.120000 71.890000  17.745000 ;
      RECT  9.320000   0.000000 16.845000   7.315000 ;
      RECT  9.320000   0.000000 16.845000  10.145000 ;
      RECT  9.320000   3.535000 19.675000  12.665000 ;
      RECT  9.320000   7.315000 19.675000   7.465000 ;
      RECT  9.320000   7.465000 19.825000   7.615000 ;
      RECT  9.320000   7.615000 19.975000   7.765000 ;
      RECT  9.320000   7.765000 20.125000   7.915000 ;
      RECT  9.320000   7.915000 20.275000   8.065000 ;
      RECT  9.320000   8.065000 20.425000   8.215000 ;
      RECT  9.320000   8.215000 20.575000   8.365000 ;
      RECT  9.320000   8.365000 20.725000   8.515000 ;
      RECT  9.320000   8.515000 20.875000   8.665000 ;
      RECT  9.320000   8.665000 21.025000   8.815000 ;
      RECT  9.320000   8.815000 21.175000   8.965000 ;
      RECT  9.320000   8.965000 21.325000   9.115000 ;
      RECT  9.320000   9.115000 21.475000   9.265000 ;
      RECT  9.320000   9.265000 21.625000   9.415000 ;
      RECT  9.320000   9.415000 21.775000   9.565000 ;
      RECT  9.320000   9.565000 21.925000   9.715000 ;
      RECT  9.320000   9.715000 22.075000   9.865000 ;
      RECT  9.320000   9.865000 22.225000  10.015000 ;
      RECT  9.320000  10.015000 22.375000  10.145000 ;
      RECT  9.320000  12.665000 12.325000  17.785000 ;
      RECT  9.320000  16.160000 71.790000  16.310000 ;
      RECT  9.345000  32.630000 71.790000  32.780000 ;
      RECT  9.495000  32.780000 71.790000  32.930000 ;
      RECT  9.560000  32.930000 71.790000  32.995000 ;
      RECT 10.695000  19.030000 68.785000  29.885000 ;
      RECT 10.750000  29.885000 68.785000  29.940000 ;
      RECT 10.750000  29.885000 68.785000  29.940000 ;
      RECT 10.805000  18.920000 68.785000  19.030000 ;
      RECT 10.805000  18.920000 68.785000  19.030000 ;
      RECT 10.805000  29.940000 68.785000  29.995000 ;
      RECT 10.805000  29.940000 68.785000  29.995000 ;
      RECT 10.955000  18.770000 68.785000  18.920000 ;
      RECT 10.955000  18.770000 68.785000  18.920000 ;
      RECT 11.105000  18.620000 68.785000  18.770000 ;
      RECT 11.105000  18.620000 68.785000  18.770000 ;
      RECT 11.255000  18.470000 68.785000  18.620000 ;
      RECT 11.255000  18.470000 68.785000  18.620000 ;
      RECT 11.405000  18.320000 68.785000  18.470000 ;
      RECT 11.405000  18.320000 68.785000  18.470000 ;
      RECT 11.555000  18.170000 68.785000  18.320000 ;
      RECT 11.555000  18.170000 68.785000  18.320000 ;
      RECT 11.570000  18.155000 24.770000  18.170000 ;
      RECT 11.570000  18.155000 24.770000  18.170000 ;
      RECT 11.720000  18.005000 24.770000  18.155000 ;
      RECT 11.720000  18.005000 24.770000  18.155000 ;
      RECT 11.870000  17.855000 24.770000  18.005000 ;
      RECT 11.870000  17.855000 24.770000  18.005000 ;
      RECT 12.020000  17.705000 24.770000  17.855000 ;
      RECT 12.020000  17.705000 24.770000  17.855000 ;
      RECT 12.170000  17.555000 24.770000  17.705000 ;
      RECT 12.170000  17.555000 24.770000  17.705000 ;
      RECT 12.320000   3.000000 13.845000   6.535000 ;
      RECT 12.320000   6.535000 16.670000   8.560000 ;
      RECT 12.320000   8.560000 16.670000   8.710000 ;
      RECT 12.320000   8.560000 16.670000   8.710000 ;
      RECT 12.320000   8.710000 16.825000   8.860000 ;
      RECT 12.320000   8.710000 16.825000   8.860000 ;
      RECT 12.320000   8.860000 16.970000   9.010000 ;
      RECT 12.320000   8.860000 16.970000   9.010000 ;
      RECT 12.320000   9.010000 17.125000   9.160000 ;
      RECT 12.320000   9.010000 17.125000   9.160000 ;
      RECT 12.320000   9.160000 17.275000   9.310000 ;
      RECT 12.320000   9.160000 17.275000   9.310000 ;
      RECT 12.320000   9.310000 17.420000   9.460000 ;
      RECT 12.320000   9.310000 17.420000   9.460000 ;
      RECT 12.320000   9.460000 17.575000   9.610000 ;
      RECT 12.320000   9.460000 17.575000   9.610000 ;
      RECT 12.320000   9.610000 17.720000   9.760000 ;
      RECT 12.320000   9.610000 17.720000   9.760000 ;
      RECT 12.320000   9.760000 17.875000   9.910000 ;
      RECT 12.320000   9.760000 17.875000   9.910000 ;
      RECT 12.320000   9.910000 18.025000  10.060000 ;
      RECT 12.320000   9.910000 18.025000  10.060000 ;
      RECT 12.320000  10.060000 18.170000  10.210000 ;
      RECT 12.320000  10.060000 18.170000  10.210000 ;
      RECT 12.320000  10.210000 18.325000  10.360000 ;
      RECT 12.320000  10.210000 18.325000  10.360000 ;
      RECT 12.320000  10.360000 18.470000  10.510000 ;
      RECT 12.320000  10.360000 18.470000  10.510000 ;
      RECT 12.320000  10.510000 18.625000  10.660000 ;
      RECT 12.320000  10.510000 18.625000  10.660000 ;
      RECT 12.320000  10.660000 18.775000  10.810000 ;
      RECT 12.320000  10.660000 18.775000  10.810000 ;
      RECT 12.320000  10.810000 18.920000  10.960000 ;
      RECT 12.320000  10.810000 18.920000  10.960000 ;
      RECT 12.320000  10.960000 19.075000  11.110000 ;
      RECT 12.320000  10.960000 19.075000  11.110000 ;
      RECT 12.320000  11.110000 19.220000  11.260000 ;
      RECT 12.320000  11.110000 19.220000  11.260000 ;
      RECT 12.320000  11.260000 19.375000  11.390000 ;
      RECT 12.320000  11.260000 19.375000  11.390000 ;
      RECT 12.320000  11.390000 19.505000  15.665000 ;
      RECT 12.320000  15.665000 24.770000  17.405000 ;
      RECT 12.320000  17.405000 24.770000  17.555000 ;
      RECT 12.320000  17.405000 24.770000  17.555000 ;
      RECT 19.210000   0.000000 19.775000   3.435000 ;
      RECT 19.310000   0.000000 19.675000   3.535000 ;
      RECT 19.500000  10.145000 22.505000  12.665000 ;
      RECT 19.500000  12.665000 27.770000  15.170000 ;
      RECT 19.505000  15.170000 32.305000  18.170000 ;
      RECT 19.505000  18.170000 32.300000  18.175000 ;
      RECT 21.525000   0.000000 28.635000   6.545000 ;
      RECT 21.525000   6.545000 28.635000   9.370000 ;
      RECT 21.625000   0.000000 28.535000   3.005000 ;
      RECT 21.625000   3.005000 24.630000   3.500000 ;
      RECT 21.625000   3.500000 28.535000   6.505000 ;
      RECT 21.775000   6.505000 28.535000   6.655000 ;
      RECT 21.925000   6.655000 28.535000   6.805000 ;
      RECT 22.075000   6.805000 28.535000   6.955000 ;
      RECT 22.225000   6.955000 28.535000   7.105000 ;
      RECT 22.375000   7.105000 28.535000   7.255000 ;
      RECT 22.525000   7.255000 28.535000   7.405000 ;
      RECT 22.575000  33.095000 71.890000  34.425000 ;
      RECT 22.675000   7.405000 28.535000   7.555000 ;
      RECT 22.675000  31.130000 25.680000  34.525000 ;
      RECT 22.825000   7.555000 28.535000   7.705000 ;
      RECT 22.975000   7.705000 28.535000   7.855000 ;
      RECT 23.125000   7.855000 28.535000   8.005000 ;
      RECT 23.275000   8.005000 28.535000   8.155000 ;
      RECT 23.425000   8.155000 28.535000   8.305000 ;
      RECT 23.575000   8.305000 28.535000   8.455000 ;
      RECT 23.725000   8.455000 28.535000   8.605000 ;
      RECT 23.875000   8.605000 28.535000   8.755000 ;
      RECT 24.025000   8.755000 28.535000   8.905000 ;
      RECT 24.175000   8.905000 28.535000   9.055000 ;
      RECT 24.325000   9.055000 28.535000   9.205000 ;
      RECT 24.350000   9.370000 28.635000   9.720000 ;
      RECT 24.350000   9.720000 27.870000  10.485000 ;
      RECT 24.350000  10.485000 27.870000  12.565000 ;
      RECT 24.450000   9.205000 28.535000   9.330000 ;
      RECT 24.450000   9.330000 28.535000   9.680000 ;
      RECT 24.450000   9.680000 27.770000  12.665000 ;
      RECT 24.450000   9.680000 28.385000   9.830000 ;
      RECT 24.450000   9.830000 28.235000   9.980000 ;
      RECT 24.450000   9.980000 28.085000  10.130000 ;
      RECT 24.450000  10.130000 27.935000  10.280000 ;
      RECT 24.450000  10.280000 27.785000  10.430000 ;
      RECT 24.450000  10.430000 27.770000  10.445000 ;
      RECT 24.625000   3.000000 25.535000   5.260000 ;
      RECT 24.625000   3.000000 25.535000   5.260000 ;
      RECT 24.770000  18.175000 32.300000  20.790000 ;
      RECT 25.530000   3.005000 28.535000   3.500000 ;
      RECT 25.675000  29.990000 68.785000  37.525000 ;
      RECT 29.200000  11.035000 71.890000  15.070000 ;
      RECT 29.300000  11.075000 33.065000  14.080000 ;
      RECT 29.300000  14.080000 32.305000  15.170000 ;
      RECT 29.315000  11.060000 71.790000  11.075000 ;
      RECT 29.465000  10.910000 71.790000  11.060000 ;
      RECT 29.615000  10.760000 71.790000  10.910000 ;
      RECT 29.765000  10.610000 71.790000  10.760000 ;
      RECT 29.915000  10.460000 71.790000  10.610000 ;
      RECT 29.965000   0.000000 71.890000  10.270000 ;
      RECT 29.965000  10.270000 71.890000  11.035000 ;
      RECT 30.065000   0.000000 71.790000   3.005000 ;
      RECT 30.065000   3.005000 33.070000  11.075000 ;
      RECT 30.065000  10.310000 71.790000  10.460000 ;
      RECT 32.300000  12.320000 68.785000  18.170000 ;
      RECT 32.315000  12.305000 68.785000  12.320000 ;
      RECT 32.315000  12.305000 68.785000  12.320000 ;
      RECT 32.465000  12.155000 68.785000  12.305000 ;
      RECT 32.465000  12.155000 68.785000  12.305000 ;
      RECT 32.615000  12.005000 68.785000  12.155000 ;
      RECT 32.615000  12.005000 68.785000  12.155000 ;
      RECT 32.765000  11.855000 68.785000  12.005000 ;
      RECT 32.765000  11.855000 68.785000  12.005000 ;
      RECT 32.915000  11.705000 68.785000  11.855000 ;
      RECT 32.915000  11.705000 68.785000  11.855000 ;
      RECT 33.065000   3.000000 68.785000  11.555000 ;
      RECT 33.065000  11.555000 68.785000  11.705000 ;
      RECT 33.065000  11.555000 68.785000  11.705000 ;
      RECT 61.455000  71.765000 64.460000  95.045000 ;
      RECT 61.460000  95.045000 69.390000  98.050000 ;
      RECT 66.290000  72.525000 75.000000  94.945000 ;
      RECT 66.390000  72.565000 70.635000  75.570000 ;
      RECT 66.390000  75.570000 69.395000  95.045000 ;
      RECT 66.525000  72.430000 75.000000  72.565000 ;
      RECT 66.675000  72.280000 75.000000  72.430000 ;
      RECT 66.825000  72.130000 75.000000  72.280000 ;
      RECT 66.975000  71.980000 75.000000  72.130000 ;
      RECT 67.125000  71.830000 75.000000  71.980000 ;
      RECT 67.275000  71.680000 75.000000  71.830000 ;
      RECT 67.425000  71.530000 75.000000  71.680000 ;
      RECT 67.545000  61.430000 71.790000  64.435000 ;
      RECT 67.575000  71.380000 75.000000  71.530000 ;
      RECT 67.725000  71.230000 75.000000  71.380000 ;
      RECT 67.875000  71.080000 75.000000  71.230000 ;
      RECT 68.025000  70.930000 75.000000  71.080000 ;
      RECT 68.175000  70.780000 75.000000  70.930000 ;
      RECT 68.325000  70.630000 75.000000  70.780000 ;
      RECT 68.475000  70.480000 75.000000  70.630000 ;
      RECT 68.625000  70.330000 75.000000  70.480000 ;
      RECT 68.775000  70.180000 75.000000  70.330000 ;
      RECT 68.785000   3.005000 71.790000  61.430000 ;
      RECT 68.925000  70.030000 75.000000  70.180000 ;
      RECT 69.075000  69.880000 75.000000  70.030000 ;
      RECT 69.225000  69.730000 75.000000  69.880000 ;
      RECT 69.375000  69.580000 75.000000  69.730000 ;
      RECT 69.390000  73.810000 72.000000  98.045000 ;
      RECT 69.445000  73.755000 72.000000  73.810000 ;
      RECT 69.445000  73.755000 72.000000  73.810000 ;
      RECT 69.525000  69.430000 75.000000  69.580000 ;
      RECT 69.595000  73.605000 72.000000  73.755000 ;
      RECT 69.595000  73.605000 72.000000  73.755000 ;
      RECT 69.675000  69.280000 75.000000  69.430000 ;
      RECT 69.745000  73.455000 72.000000  73.605000 ;
      RECT 69.745000  73.455000 72.000000  73.605000 ;
      RECT 69.825000  69.130000 75.000000  69.280000 ;
      RECT 69.895000  73.305000 72.000000  73.455000 ;
      RECT 69.895000  73.305000 72.000000  73.455000 ;
      RECT 69.975000  68.980000 75.000000  69.130000 ;
      RECT 70.045000  73.155000 72.000000  73.305000 ;
      RECT 70.045000  73.155000 72.000000  73.305000 ;
      RECT 70.125000  68.830000 75.000000  68.980000 ;
      RECT 70.195000  73.005000 72.000000  73.155000 ;
      RECT 70.195000  73.005000 72.000000  73.155000 ;
      RECT 70.275000  68.680000 75.000000  68.830000 ;
      RECT 70.345000  72.855000 72.000000  73.005000 ;
      RECT 70.345000  72.855000 72.000000  73.005000 ;
      RECT 70.425000  68.530000 75.000000  68.680000 ;
      RECT 70.495000  72.705000 72.000000  72.855000 ;
      RECT 70.495000  72.705000 72.000000  72.855000 ;
      RECT 70.575000  68.380000 75.000000  68.530000 ;
      RECT 70.645000  72.555000 72.000000  72.705000 ;
      RECT 70.645000  72.555000 72.000000  72.705000 ;
      RECT 70.725000  68.230000 75.000000  68.380000 ;
      RECT 70.795000  72.405000 72.000000  72.555000 ;
      RECT 70.795000  72.405000 72.000000  72.555000 ;
      RECT 70.875000  68.080000 75.000000  68.230000 ;
      RECT 70.945000  72.255000 72.000000  72.405000 ;
      RECT 70.945000  72.255000 72.000000  72.405000 ;
      RECT 71.025000  67.930000 75.000000  68.080000 ;
      RECT 71.095000  72.105000 72.000000  72.255000 ;
      RECT 71.095000  72.105000 72.000000  72.255000 ;
      RECT 71.175000  67.780000 75.000000  67.930000 ;
      RECT 71.245000  71.955000 72.000000  72.105000 ;
      RECT 71.245000  71.955000 72.000000  72.105000 ;
      RECT 71.325000  67.630000 75.000000  67.780000 ;
      RECT 71.395000  71.805000 72.000000  71.955000 ;
      RECT 71.395000  71.805000 72.000000  71.955000 ;
      RECT 71.475000  67.480000 75.000000  67.630000 ;
      RECT 71.545000  71.655000 72.000000  71.805000 ;
      RECT 71.545000  71.655000 72.000000  71.805000 ;
      RECT 71.625000  67.330000 75.000000  67.480000 ;
      RECT 71.695000  71.505000 72.000000  71.655000 ;
      RECT 71.695000  71.505000 72.000000  71.655000 ;
      RECT 71.775000  67.180000 75.000000  67.330000 ;
      RECT 71.845000  71.355000 72.000000  71.505000 ;
      RECT 71.845000  71.355000 72.000000  71.505000 ;
      RECT 71.925000  67.030000 75.000000  67.180000 ;
      RECT 71.995000  72.565000 75.000000 196.995000 ;
      RECT 72.075000  66.880000 75.000000  67.030000 ;
      RECT 72.225000  66.730000 75.000000  66.880000 ;
      RECT 72.375000  66.580000 75.000000  66.730000 ;
      RECT 72.525000  66.430000 75.000000  66.580000 ;
      RECT 72.675000  66.280000 75.000000  66.430000 ;
      RECT 72.825000  66.130000 75.000000  66.280000 ;
      RECT 72.975000  65.980000 75.000000  66.130000 ;
      RECT 73.125000  65.830000 75.000000  65.980000 ;
      RECT 73.275000  65.680000 75.000000  65.830000 ;
      RECT 73.425000  65.530000 75.000000  65.680000 ;
      RECT 73.560000   0.000000 75.000000  49.195000 ;
      RECT 73.560000  49.195000 75.000000  49.860000 ;
      RECT 73.575000  65.380000 75.000000  65.530000 ;
      RECT 73.660000   0.000000 75.000000  49.155000 ;
      RECT 73.725000  65.230000 75.000000  65.380000 ;
      RECT 73.810000  49.155000 75.000000  49.305000 ;
      RECT 73.875000  65.080000 75.000000  65.230000 ;
      RECT 73.960000  49.305000 75.000000  49.455000 ;
      RECT 74.025000  64.930000 75.000000  65.080000 ;
      RECT 74.110000  49.455000 75.000000  49.605000 ;
      RECT 74.175000  64.780000 75.000000  64.930000 ;
      RECT 74.225000  49.860000 75.000000  64.590000 ;
      RECT 74.225000  64.590000 75.000000  72.525000 ;
      RECT 74.260000  49.605000 75.000000  49.755000 ;
      RECT 74.325000  49.755000 75.000000  49.820000 ;
      RECT 74.325000  49.820000 75.000000  64.630000 ;
      RECT 74.325000  64.630000 75.000000  64.780000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   0.000000 75.000000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000   7.885000 75.000000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  13.935000 75.000000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  18.785000 75.000000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  24.835000 75.000000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  30.885000 75.000000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  35.735000 75.000000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  40.585000 75.000000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  46.635000 75.000000  47.435000 ;
      RECT  0.000000  57.035000 75.000000  57.835000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  63.085000 75.000000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  68.935000 75.000000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.570000  47.435000 73.430000  57.035000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000  19.385000 73.330000  41.230000 ;
      RECT  1.670000  36.335000 73.330000  41.230000 ;
      RECT  1.670000  36.335000 73.330000  41.230000 ;
      RECT  1.670000  41.185000 75.000000  41.255000 ;
      RECT  1.670000  41.230000 73.255000  41.255000 ;
      RECT  1.670000  46.570000 73.255000  46.590000 ;
      RECT  1.670000  46.570000 73.255000  57.135000 ;
      RECT  1.670000  46.570000 75.000000  46.635000 ;
      RECT  1.670000  46.590000 73.330000  57.135000 ;
      RECT  1.670000  46.590000 73.330000  57.135000 ;
      RECT  1.670000  46.590000 73.330000  95.400000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT  4.120000  41.230000 73.255000  46.570000 ;
      RECT  4.120000  41.255000 73.255000  46.570000 ;
      RECT  4.120000  41.255000 73.255000  57.135000 ;
      RECT  4.120000  41.255000 75.000000  41.285000 ;
      RECT  4.120000  41.285000 73.430000  41.330000 ;
      RECT  4.120000  41.330000 73.355000  46.490000 ;
      RECT  4.120000  46.490000 73.430000  46.535000 ;
      RECT  4.120000  46.535000 75.000000  46.570000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000 75.000000   1.335000 ;
      RECT  0.000000  36.035000 75.000000  36.040000 ;
      RECT  0.000000  95.785000 75.000000 126.315000 ;
      RECT  0.000000 126.315000 28.895000 146.425000 ;
      RECT  0.000000 146.425000 75.000000 174.985000 ;
      RECT  1.765000  14.235000 73.235000  19.085000 ;
      RECT  2.070000   1.335000 72.930000  14.235000 ;
      RECT  2.070000  19.085000 72.930000  95.785000 ;
      RECT  2.070000 174.985000 72.930000 200.000000 ;
      RECT 42.790000 126.315000 75.000000 146.425000 ;
  END
END sky130_fd_io__top_xres4v2


MACRO sky130_fd_io__overlay_vssio_lvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.500000 171.195000 12.900000 198.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500000 23.840000 24.400000 28.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 23.840000 74.290000 28.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.045000 171.195000 74.700000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000  1.270000 173.835000 ;
        RECT 0.000000 173.835000 12.900000 197.970000 ;
        RECT 0.000000 197.970000  1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 24.375000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.075000 173.835000 75.000000 197.970000 ;
        RECT 73.730000 173.785000 75.000000 173.835000 ;
        RECT 73.730000 197.970000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.590000  23.910000  0.790000  24.110000 ;
        RECT  0.590000  24.340000  0.790000  24.540000 ;
        RECT  0.590000  24.770000  0.790000  24.970000 ;
        RECT  0.590000  25.200000  0.790000  25.400000 ;
        RECT  0.590000  25.630000  0.790000  25.830000 ;
        RECT  0.590000  26.060000  0.790000  26.260000 ;
        RECT  0.590000  26.490000  0.790000  26.690000 ;
        RECT  0.590000  26.920000  0.790000  27.120000 ;
        RECT  0.590000  27.350000  0.790000  27.550000 ;
        RECT  0.590000  27.780000  0.790000  27.980000 ;
        RECT  0.590000  28.210000  0.790000  28.410000 ;
        RECT  0.615000 173.900000  0.815000 174.100000 ;
        RECT  0.615000 174.300000  0.815000 174.500000 ;
        RECT  0.615000 174.700000  0.815000 174.900000 ;
        RECT  0.615000 175.100000  0.815000 175.300000 ;
        RECT  0.615000 175.500000  0.815000 175.700000 ;
        RECT  0.615000 175.900000  0.815000 176.100000 ;
        RECT  0.615000 176.300000  0.815000 176.500000 ;
        RECT  0.615000 176.700000  0.815000 176.900000 ;
        RECT  0.615000 177.100000  0.815000 177.300000 ;
        RECT  0.615000 177.500000  0.815000 177.700000 ;
        RECT  0.615000 177.900000  0.815000 178.100000 ;
        RECT  0.615000 178.300000  0.815000 178.500000 ;
        RECT  0.615000 178.700000  0.815000 178.900000 ;
        RECT  0.615000 179.100000  0.815000 179.300000 ;
        RECT  0.615000 179.500000  0.815000 179.700000 ;
        RECT  0.615000 179.900000  0.815000 180.100000 ;
        RECT  0.615000 180.300000  0.815000 180.500000 ;
        RECT  0.615000 180.700000  0.815000 180.900000 ;
        RECT  0.615000 181.100000  0.815000 181.300000 ;
        RECT  0.615000 181.505000  0.815000 181.705000 ;
        RECT  0.615000 181.910000  0.815000 182.110000 ;
        RECT  0.615000 182.315000  0.815000 182.515000 ;
        RECT  0.615000 182.720000  0.815000 182.920000 ;
        RECT  0.615000 183.125000  0.815000 183.325000 ;
        RECT  0.615000 183.530000  0.815000 183.730000 ;
        RECT  0.615000 183.935000  0.815000 184.135000 ;
        RECT  0.615000 184.340000  0.815000 184.540000 ;
        RECT  0.615000 184.745000  0.815000 184.945000 ;
        RECT  0.615000 185.150000  0.815000 185.350000 ;
        RECT  0.615000 185.555000  0.815000 185.755000 ;
        RECT  0.615000 185.960000  0.815000 186.160000 ;
        RECT  0.615000 186.365000  0.815000 186.565000 ;
        RECT  0.615000 186.770000  0.815000 186.970000 ;
        RECT  0.615000 187.175000  0.815000 187.375000 ;
        RECT  0.615000 187.580000  0.815000 187.780000 ;
        RECT  0.615000 187.985000  0.815000 188.185000 ;
        RECT  0.615000 188.390000  0.815000 188.590000 ;
        RECT  0.615000 188.795000  0.815000 188.995000 ;
        RECT  0.615000 189.200000  0.815000 189.400000 ;
        RECT  0.615000 189.605000  0.815000 189.805000 ;
        RECT  0.615000 190.010000  0.815000 190.210000 ;
        RECT  0.615000 190.415000  0.815000 190.615000 ;
        RECT  0.615000 190.820000  0.815000 191.020000 ;
        RECT  0.615000 191.225000  0.815000 191.425000 ;
        RECT  0.615000 191.630000  0.815000 191.830000 ;
        RECT  0.615000 192.035000  0.815000 192.235000 ;
        RECT  0.615000 192.440000  0.815000 192.640000 ;
        RECT  0.615000 192.845000  0.815000 193.045000 ;
        RECT  0.615000 193.250000  0.815000 193.450000 ;
        RECT  0.615000 193.655000  0.815000 193.855000 ;
        RECT  0.615000 194.060000  0.815000 194.260000 ;
        RECT  0.615000 194.465000  0.815000 194.665000 ;
        RECT  0.615000 194.870000  0.815000 195.070000 ;
        RECT  0.615000 195.275000  0.815000 195.475000 ;
        RECT  0.615000 195.680000  0.815000 195.880000 ;
        RECT  0.615000 196.085000  0.815000 196.285000 ;
        RECT  0.615000 196.490000  0.815000 196.690000 ;
        RECT  0.615000 196.895000  0.815000 197.095000 ;
        RECT  0.615000 197.300000  0.815000 197.500000 ;
        RECT  0.615000 197.705000  0.815000 197.905000 ;
        RECT  1.000000  23.910000  1.200000  24.110000 ;
        RECT  1.000000  24.340000  1.200000  24.540000 ;
        RECT  1.000000  24.770000  1.200000  24.970000 ;
        RECT  1.000000  25.200000  1.200000  25.400000 ;
        RECT  1.000000  25.630000  1.200000  25.830000 ;
        RECT  1.000000  26.060000  1.200000  26.260000 ;
        RECT  1.000000  26.490000  1.200000  26.690000 ;
        RECT  1.000000  26.920000  1.200000  27.120000 ;
        RECT  1.000000  27.350000  1.200000  27.550000 ;
        RECT  1.000000  27.780000  1.200000  27.980000 ;
        RECT  1.000000  28.210000  1.200000  28.410000 ;
        RECT  1.015000 173.900000  1.215000 174.100000 ;
        RECT  1.015000 174.300000  1.215000 174.500000 ;
        RECT  1.015000 174.700000  1.215000 174.900000 ;
        RECT  1.015000 175.100000  1.215000 175.300000 ;
        RECT  1.015000 175.500000  1.215000 175.700000 ;
        RECT  1.015000 175.900000  1.215000 176.100000 ;
        RECT  1.015000 176.300000  1.215000 176.500000 ;
        RECT  1.015000 176.700000  1.215000 176.900000 ;
        RECT  1.015000 177.100000  1.215000 177.300000 ;
        RECT  1.015000 177.500000  1.215000 177.700000 ;
        RECT  1.015000 177.900000  1.215000 178.100000 ;
        RECT  1.015000 178.300000  1.215000 178.500000 ;
        RECT  1.015000 178.700000  1.215000 178.900000 ;
        RECT  1.015000 179.100000  1.215000 179.300000 ;
        RECT  1.015000 179.500000  1.215000 179.700000 ;
        RECT  1.015000 179.900000  1.215000 180.100000 ;
        RECT  1.015000 180.300000  1.215000 180.500000 ;
        RECT  1.015000 180.700000  1.215000 180.900000 ;
        RECT  1.015000 181.100000  1.215000 181.300000 ;
        RECT  1.015000 181.505000  1.215000 181.705000 ;
        RECT  1.015000 181.910000  1.215000 182.110000 ;
        RECT  1.015000 182.315000  1.215000 182.515000 ;
        RECT  1.015000 182.720000  1.215000 182.920000 ;
        RECT  1.015000 183.125000  1.215000 183.325000 ;
        RECT  1.015000 183.530000  1.215000 183.730000 ;
        RECT  1.015000 183.935000  1.215000 184.135000 ;
        RECT  1.015000 184.340000  1.215000 184.540000 ;
        RECT  1.015000 184.745000  1.215000 184.945000 ;
        RECT  1.015000 185.150000  1.215000 185.350000 ;
        RECT  1.015000 185.555000  1.215000 185.755000 ;
        RECT  1.015000 185.960000  1.215000 186.160000 ;
        RECT  1.015000 186.365000  1.215000 186.565000 ;
        RECT  1.015000 186.770000  1.215000 186.970000 ;
        RECT  1.015000 187.175000  1.215000 187.375000 ;
        RECT  1.015000 187.580000  1.215000 187.780000 ;
        RECT  1.015000 187.985000  1.215000 188.185000 ;
        RECT  1.015000 188.390000  1.215000 188.590000 ;
        RECT  1.015000 188.795000  1.215000 188.995000 ;
        RECT  1.015000 189.200000  1.215000 189.400000 ;
        RECT  1.015000 189.605000  1.215000 189.805000 ;
        RECT  1.015000 190.010000  1.215000 190.210000 ;
        RECT  1.015000 190.415000  1.215000 190.615000 ;
        RECT  1.015000 190.820000  1.215000 191.020000 ;
        RECT  1.015000 191.225000  1.215000 191.425000 ;
        RECT  1.015000 191.630000  1.215000 191.830000 ;
        RECT  1.015000 192.035000  1.215000 192.235000 ;
        RECT  1.015000 192.440000  1.215000 192.640000 ;
        RECT  1.015000 192.845000  1.215000 193.045000 ;
        RECT  1.015000 193.250000  1.215000 193.450000 ;
        RECT  1.015000 193.655000  1.215000 193.855000 ;
        RECT  1.015000 194.060000  1.215000 194.260000 ;
        RECT  1.015000 194.465000  1.215000 194.665000 ;
        RECT  1.015000 194.870000  1.215000 195.070000 ;
        RECT  1.015000 195.275000  1.215000 195.475000 ;
        RECT  1.015000 195.680000  1.215000 195.880000 ;
        RECT  1.015000 196.085000  1.215000 196.285000 ;
        RECT  1.015000 196.490000  1.215000 196.690000 ;
        RECT  1.015000 196.895000  1.215000 197.095000 ;
        RECT  1.015000 197.300000  1.215000 197.500000 ;
        RECT  1.015000 197.705000  1.215000 197.905000 ;
        RECT  1.410000  23.910000  1.610000  24.110000 ;
        RECT  1.410000  24.340000  1.610000  24.540000 ;
        RECT  1.410000  24.770000  1.610000  24.970000 ;
        RECT  1.410000  25.200000  1.610000  25.400000 ;
        RECT  1.410000  25.630000  1.610000  25.830000 ;
        RECT  1.410000  26.060000  1.610000  26.260000 ;
        RECT  1.410000  26.490000  1.610000  26.690000 ;
        RECT  1.410000  26.920000  1.610000  27.120000 ;
        RECT  1.410000  27.350000  1.610000  27.550000 ;
        RECT  1.410000  27.780000  1.610000  27.980000 ;
        RECT  1.410000  28.210000  1.610000  28.410000 ;
        RECT  1.415000 173.900000  1.615000 174.100000 ;
        RECT  1.415000 174.300000  1.615000 174.500000 ;
        RECT  1.415000 174.700000  1.615000 174.900000 ;
        RECT  1.415000 175.100000  1.615000 175.300000 ;
        RECT  1.415000 175.500000  1.615000 175.700000 ;
        RECT  1.415000 175.900000  1.615000 176.100000 ;
        RECT  1.415000 176.300000  1.615000 176.500000 ;
        RECT  1.415000 176.700000  1.615000 176.900000 ;
        RECT  1.415000 177.100000  1.615000 177.300000 ;
        RECT  1.415000 177.500000  1.615000 177.700000 ;
        RECT  1.415000 177.900000  1.615000 178.100000 ;
        RECT  1.415000 178.300000  1.615000 178.500000 ;
        RECT  1.415000 178.700000  1.615000 178.900000 ;
        RECT  1.415000 179.100000  1.615000 179.300000 ;
        RECT  1.415000 179.500000  1.615000 179.700000 ;
        RECT  1.415000 179.900000  1.615000 180.100000 ;
        RECT  1.415000 180.300000  1.615000 180.500000 ;
        RECT  1.415000 180.700000  1.615000 180.900000 ;
        RECT  1.415000 181.100000  1.615000 181.300000 ;
        RECT  1.415000 181.505000  1.615000 181.705000 ;
        RECT  1.415000 181.910000  1.615000 182.110000 ;
        RECT  1.415000 182.315000  1.615000 182.515000 ;
        RECT  1.415000 182.720000  1.615000 182.920000 ;
        RECT  1.415000 183.125000  1.615000 183.325000 ;
        RECT  1.415000 183.530000  1.615000 183.730000 ;
        RECT  1.415000 183.935000  1.615000 184.135000 ;
        RECT  1.415000 184.340000  1.615000 184.540000 ;
        RECT  1.415000 184.745000  1.615000 184.945000 ;
        RECT  1.415000 185.150000  1.615000 185.350000 ;
        RECT  1.415000 185.555000  1.615000 185.755000 ;
        RECT  1.415000 185.960000  1.615000 186.160000 ;
        RECT  1.415000 186.365000  1.615000 186.565000 ;
        RECT  1.415000 186.770000  1.615000 186.970000 ;
        RECT  1.415000 187.175000  1.615000 187.375000 ;
        RECT  1.415000 187.580000  1.615000 187.780000 ;
        RECT  1.415000 187.985000  1.615000 188.185000 ;
        RECT  1.415000 188.390000  1.615000 188.590000 ;
        RECT  1.415000 188.795000  1.615000 188.995000 ;
        RECT  1.415000 189.200000  1.615000 189.400000 ;
        RECT  1.415000 189.605000  1.615000 189.805000 ;
        RECT  1.415000 190.010000  1.615000 190.210000 ;
        RECT  1.415000 190.415000  1.615000 190.615000 ;
        RECT  1.415000 190.820000  1.615000 191.020000 ;
        RECT  1.415000 191.225000  1.615000 191.425000 ;
        RECT  1.415000 191.630000  1.615000 191.830000 ;
        RECT  1.415000 192.035000  1.615000 192.235000 ;
        RECT  1.415000 192.440000  1.615000 192.640000 ;
        RECT  1.415000 192.845000  1.615000 193.045000 ;
        RECT  1.415000 193.250000  1.615000 193.450000 ;
        RECT  1.415000 193.655000  1.615000 193.855000 ;
        RECT  1.415000 194.060000  1.615000 194.260000 ;
        RECT  1.415000 194.465000  1.615000 194.665000 ;
        RECT  1.415000 194.870000  1.615000 195.070000 ;
        RECT  1.415000 195.275000  1.615000 195.475000 ;
        RECT  1.415000 195.680000  1.615000 195.880000 ;
        RECT  1.415000 196.085000  1.615000 196.285000 ;
        RECT  1.415000 196.490000  1.615000 196.690000 ;
        RECT  1.415000 196.895000  1.615000 197.095000 ;
        RECT  1.415000 197.300000  1.615000 197.500000 ;
        RECT  1.415000 197.705000  1.615000 197.905000 ;
        RECT  1.815000 173.900000  2.015000 174.100000 ;
        RECT  1.815000 174.300000  2.015000 174.500000 ;
        RECT  1.815000 174.700000  2.015000 174.900000 ;
        RECT  1.815000 175.100000  2.015000 175.300000 ;
        RECT  1.815000 175.500000  2.015000 175.700000 ;
        RECT  1.815000 175.900000  2.015000 176.100000 ;
        RECT  1.815000 176.300000  2.015000 176.500000 ;
        RECT  1.815000 176.700000  2.015000 176.900000 ;
        RECT  1.815000 177.100000  2.015000 177.300000 ;
        RECT  1.815000 177.500000  2.015000 177.700000 ;
        RECT  1.815000 177.900000  2.015000 178.100000 ;
        RECT  1.815000 178.300000  2.015000 178.500000 ;
        RECT  1.815000 178.700000  2.015000 178.900000 ;
        RECT  1.815000 179.100000  2.015000 179.300000 ;
        RECT  1.815000 179.500000  2.015000 179.700000 ;
        RECT  1.815000 179.900000  2.015000 180.100000 ;
        RECT  1.815000 180.300000  2.015000 180.500000 ;
        RECT  1.815000 180.700000  2.015000 180.900000 ;
        RECT  1.815000 181.100000  2.015000 181.300000 ;
        RECT  1.815000 181.505000  2.015000 181.705000 ;
        RECT  1.815000 181.910000  2.015000 182.110000 ;
        RECT  1.815000 182.315000  2.015000 182.515000 ;
        RECT  1.815000 182.720000  2.015000 182.920000 ;
        RECT  1.815000 183.125000  2.015000 183.325000 ;
        RECT  1.815000 183.530000  2.015000 183.730000 ;
        RECT  1.815000 183.935000  2.015000 184.135000 ;
        RECT  1.815000 184.340000  2.015000 184.540000 ;
        RECT  1.815000 184.745000  2.015000 184.945000 ;
        RECT  1.815000 185.150000  2.015000 185.350000 ;
        RECT  1.815000 185.555000  2.015000 185.755000 ;
        RECT  1.815000 185.960000  2.015000 186.160000 ;
        RECT  1.815000 186.365000  2.015000 186.565000 ;
        RECT  1.815000 186.770000  2.015000 186.970000 ;
        RECT  1.815000 187.175000  2.015000 187.375000 ;
        RECT  1.815000 187.580000  2.015000 187.780000 ;
        RECT  1.815000 187.985000  2.015000 188.185000 ;
        RECT  1.815000 188.390000  2.015000 188.590000 ;
        RECT  1.815000 188.795000  2.015000 188.995000 ;
        RECT  1.815000 189.200000  2.015000 189.400000 ;
        RECT  1.815000 189.605000  2.015000 189.805000 ;
        RECT  1.815000 190.010000  2.015000 190.210000 ;
        RECT  1.815000 190.415000  2.015000 190.615000 ;
        RECT  1.815000 190.820000  2.015000 191.020000 ;
        RECT  1.815000 191.225000  2.015000 191.425000 ;
        RECT  1.815000 191.630000  2.015000 191.830000 ;
        RECT  1.815000 192.035000  2.015000 192.235000 ;
        RECT  1.815000 192.440000  2.015000 192.640000 ;
        RECT  1.815000 192.845000  2.015000 193.045000 ;
        RECT  1.815000 193.250000  2.015000 193.450000 ;
        RECT  1.815000 193.655000  2.015000 193.855000 ;
        RECT  1.815000 194.060000  2.015000 194.260000 ;
        RECT  1.815000 194.465000  2.015000 194.665000 ;
        RECT  1.815000 194.870000  2.015000 195.070000 ;
        RECT  1.815000 195.275000  2.015000 195.475000 ;
        RECT  1.815000 195.680000  2.015000 195.880000 ;
        RECT  1.815000 196.085000  2.015000 196.285000 ;
        RECT  1.815000 196.490000  2.015000 196.690000 ;
        RECT  1.815000 196.895000  2.015000 197.095000 ;
        RECT  1.815000 197.300000  2.015000 197.500000 ;
        RECT  1.815000 197.705000  2.015000 197.905000 ;
        RECT  1.820000  23.910000  2.020000  24.110000 ;
        RECT  1.820000  24.340000  2.020000  24.540000 ;
        RECT  1.820000  24.770000  2.020000  24.970000 ;
        RECT  1.820000  25.200000  2.020000  25.400000 ;
        RECT  1.820000  25.630000  2.020000  25.830000 ;
        RECT  1.820000  26.060000  2.020000  26.260000 ;
        RECT  1.820000  26.490000  2.020000  26.690000 ;
        RECT  1.820000  26.920000  2.020000  27.120000 ;
        RECT  1.820000  27.350000  2.020000  27.550000 ;
        RECT  1.820000  27.780000  2.020000  27.980000 ;
        RECT  1.820000  28.210000  2.020000  28.410000 ;
        RECT  2.215000 173.900000  2.415000 174.100000 ;
        RECT  2.215000 174.300000  2.415000 174.500000 ;
        RECT  2.215000 174.700000  2.415000 174.900000 ;
        RECT  2.215000 175.100000  2.415000 175.300000 ;
        RECT  2.215000 175.500000  2.415000 175.700000 ;
        RECT  2.215000 175.900000  2.415000 176.100000 ;
        RECT  2.215000 176.300000  2.415000 176.500000 ;
        RECT  2.215000 176.700000  2.415000 176.900000 ;
        RECT  2.215000 177.100000  2.415000 177.300000 ;
        RECT  2.215000 177.500000  2.415000 177.700000 ;
        RECT  2.215000 177.900000  2.415000 178.100000 ;
        RECT  2.215000 178.300000  2.415000 178.500000 ;
        RECT  2.215000 178.700000  2.415000 178.900000 ;
        RECT  2.215000 179.100000  2.415000 179.300000 ;
        RECT  2.215000 179.500000  2.415000 179.700000 ;
        RECT  2.215000 179.900000  2.415000 180.100000 ;
        RECT  2.215000 180.300000  2.415000 180.500000 ;
        RECT  2.215000 180.700000  2.415000 180.900000 ;
        RECT  2.215000 181.100000  2.415000 181.300000 ;
        RECT  2.215000 181.505000  2.415000 181.705000 ;
        RECT  2.215000 181.910000  2.415000 182.110000 ;
        RECT  2.215000 182.315000  2.415000 182.515000 ;
        RECT  2.215000 182.720000  2.415000 182.920000 ;
        RECT  2.215000 183.125000  2.415000 183.325000 ;
        RECT  2.215000 183.530000  2.415000 183.730000 ;
        RECT  2.215000 183.935000  2.415000 184.135000 ;
        RECT  2.215000 184.340000  2.415000 184.540000 ;
        RECT  2.215000 184.745000  2.415000 184.945000 ;
        RECT  2.215000 185.150000  2.415000 185.350000 ;
        RECT  2.215000 185.555000  2.415000 185.755000 ;
        RECT  2.215000 185.960000  2.415000 186.160000 ;
        RECT  2.215000 186.365000  2.415000 186.565000 ;
        RECT  2.215000 186.770000  2.415000 186.970000 ;
        RECT  2.215000 187.175000  2.415000 187.375000 ;
        RECT  2.215000 187.580000  2.415000 187.780000 ;
        RECT  2.215000 187.985000  2.415000 188.185000 ;
        RECT  2.215000 188.390000  2.415000 188.590000 ;
        RECT  2.215000 188.795000  2.415000 188.995000 ;
        RECT  2.215000 189.200000  2.415000 189.400000 ;
        RECT  2.215000 189.605000  2.415000 189.805000 ;
        RECT  2.215000 190.010000  2.415000 190.210000 ;
        RECT  2.215000 190.415000  2.415000 190.615000 ;
        RECT  2.215000 190.820000  2.415000 191.020000 ;
        RECT  2.215000 191.225000  2.415000 191.425000 ;
        RECT  2.215000 191.630000  2.415000 191.830000 ;
        RECT  2.215000 192.035000  2.415000 192.235000 ;
        RECT  2.215000 192.440000  2.415000 192.640000 ;
        RECT  2.215000 192.845000  2.415000 193.045000 ;
        RECT  2.215000 193.250000  2.415000 193.450000 ;
        RECT  2.215000 193.655000  2.415000 193.855000 ;
        RECT  2.215000 194.060000  2.415000 194.260000 ;
        RECT  2.215000 194.465000  2.415000 194.665000 ;
        RECT  2.215000 194.870000  2.415000 195.070000 ;
        RECT  2.215000 195.275000  2.415000 195.475000 ;
        RECT  2.215000 195.680000  2.415000 195.880000 ;
        RECT  2.215000 196.085000  2.415000 196.285000 ;
        RECT  2.215000 196.490000  2.415000 196.690000 ;
        RECT  2.215000 196.895000  2.415000 197.095000 ;
        RECT  2.215000 197.300000  2.415000 197.500000 ;
        RECT  2.215000 197.705000  2.415000 197.905000 ;
        RECT  2.230000  23.910000  2.430000  24.110000 ;
        RECT  2.230000  24.340000  2.430000  24.540000 ;
        RECT  2.230000  24.770000  2.430000  24.970000 ;
        RECT  2.230000  25.200000  2.430000  25.400000 ;
        RECT  2.230000  25.630000  2.430000  25.830000 ;
        RECT  2.230000  26.060000  2.430000  26.260000 ;
        RECT  2.230000  26.490000  2.430000  26.690000 ;
        RECT  2.230000  26.920000  2.430000  27.120000 ;
        RECT  2.230000  27.350000  2.430000  27.550000 ;
        RECT  2.230000  27.780000  2.430000  27.980000 ;
        RECT  2.230000  28.210000  2.430000  28.410000 ;
        RECT  2.615000 173.900000  2.815000 174.100000 ;
        RECT  2.615000 174.300000  2.815000 174.500000 ;
        RECT  2.615000 174.700000  2.815000 174.900000 ;
        RECT  2.615000 175.100000  2.815000 175.300000 ;
        RECT  2.615000 175.500000  2.815000 175.700000 ;
        RECT  2.615000 175.900000  2.815000 176.100000 ;
        RECT  2.615000 176.300000  2.815000 176.500000 ;
        RECT  2.615000 176.700000  2.815000 176.900000 ;
        RECT  2.615000 177.100000  2.815000 177.300000 ;
        RECT  2.615000 177.500000  2.815000 177.700000 ;
        RECT  2.615000 177.900000  2.815000 178.100000 ;
        RECT  2.615000 178.300000  2.815000 178.500000 ;
        RECT  2.615000 178.700000  2.815000 178.900000 ;
        RECT  2.615000 179.100000  2.815000 179.300000 ;
        RECT  2.615000 179.500000  2.815000 179.700000 ;
        RECT  2.615000 179.900000  2.815000 180.100000 ;
        RECT  2.615000 180.300000  2.815000 180.500000 ;
        RECT  2.615000 180.700000  2.815000 180.900000 ;
        RECT  2.615000 181.100000  2.815000 181.300000 ;
        RECT  2.615000 181.505000  2.815000 181.705000 ;
        RECT  2.615000 181.910000  2.815000 182.110000 ;
        RECT  2.615000 182.315000  2.815000 182.515000 ;
        RECT  2.615000 182.720000  2.815000 182.920000 ;
        RECT  2.615000 183.125000  2.815000 183.325000 ;
        RECT  2.615000 183.530000  2.815000 183.730000 ;
        RECT  2.615000 183.935000  2.815000 184.135000 ;
        RECT  2.615000 184.340000  2.815000 184.540000 ;
        RECT  2.615000 184.745000  2.815000 184.945000 ;
        RECT  2.615000 185.150000  2.815000 185.350000 ;
        RECT  2.615000 185.555000  2.815000 185.755000 ;
        RECT  2.615000 185.960000  2.815000 186.160000 ;
        RECT  2.615000 186.365000  2.815000 186.565000 ;
        RECT  2.615000 186.770000  2.815000 186.970000 ;
        RECT  2.615000 187.175000  2.815000 187.375000 ;
        RECT  2.615000 187.580000  2.815000 187.780000 ;
        RECT  2.615000 187.985000  2.815000 188.185000 ;
        RECT  2.615000 188.390000  2.815000 188.590000 ;
        RECT  2.615000 188.795000  2.815000 188.995000 ;
        RECT  2.615000 189.200000  2.815000 189.400000 ;
        RECT  2.615000 189.605000  2.815000 189.805000 ;
        RECT  2.615000 190.010000  2.815000 190.210000 ;
        RECT  2.615000 190.415000  2.815000 190.615000 ;
        RECT  2.615000 190.820000  2.815000 191.020000 ;
        RECT  2.615000 191.225000  2.815000 191.425000 ;
        RECT  2.615000 191.630000  2.815000 191.830000 ;
        RECT  2.615000 192.035000  2.815000 192.235000 ;
        RECT  2.615000 192.440000  2.815000 192.640000 ;
        RECT  2.615000 192.845000  2.815000 193.045000 ;
        RECT  2.615000 193.250000  2.815000 193.450000 ;
        RECT  2.615000 193.655000  2.815000 193.855000 ;
        RECT  2.615000 194.060000  2.815000 194.260000 ;
        RECT  2.615000 194.465000  2.815000 194.665000 ;
        RECT  2.615000 194.870000  2.815000 195.070000 ;
        RECT  2.615000 195.275000  2.815000 195.475000 ;
        RECT  2.615000 195.680000  2.815000 195.880000 ;
        RECT  2.615000 196.085000  2.815000 196.285000 ;
        RECT  2.615000 196.490000  2.815000 196.690000 ;
        RECT  2.615000 196.895000  2.815000 197.095000 ;
        RECT  2.615000 197.300000  2.815000 197.500000 ;
        RECT  2.615000 197.705000  2.815000 197.905000 ;
        RECT  2.640000  23.910000  2.840000  24.110000 ;
        RECT  2.640000  24.340000  2.840000  24.540000 ;
        RECT  2.640000  24.770000  2.840000  24.970000 ;
        RECT  2.640000  25.200000  2.840000  25.400000 ;
        RECT  2.640000  25.630000  2.840000  25.830000 ;
        RECT  2.640000  26.060000  2.840000  26.260000 ;
        RECT  2.640000  26.490000  2.840000  26.690000 ;
        RECT  2.640000  26.920000  2.840000  27.120000 ;
        RECT  2.640000  27.350000  2.840000  27.550000 ;
        RECT  2.640000  27.780000  2.840000  27.980000 ;
        RECT  2.640000  28.210000  2.840000  28.410000 ;
        RECT  3.015000 173.900000  3.215000 174.100000 ;
        RECT  3.015000 174.300000  3.215000 174.500000 ;
        RECT  3.015000 174.700000  3.215000 174.900000 ;
        RECT  3.015000 175.100000  3.215000 175.300000 ;
        RECT  3.015000 175.500000  3.215000 175.700000 ;
        RECT  3.015000 175.900000  3.215000 176.100000 ;
        RECT  3.015000 176.300000  3.215000 176.500000 ;
        RECT  3.015000 176.700000  3.215000 176.900000 ;
        RECT  3.015000 177.100000  3.215000 177.300000 ;
        RECT  3.015000 177.500000  3.215000 177.700000 ;
        RECT  3.015000 177.900000  3.215000 178.100000 ;
        RECT  3.015000 178.300000  3.215000 178.500000 ;
        RECT  3.015000 178.700000  3.215000 178.900000 ;
        RECT  3.015000 179.100000  3.215000 179.300000 ;
        RECT  3.015000 179.500000  3.215000 179.700000 ;
        RECT  3.015000 179.900000  3.215000 180.100000 ;
        RECT  3.015000 180.300000  3.215000 180.500000 ;
        RECT  3.015000 180.700000  3.215000 180.900000 ;
        RECT  3.015000 181.100000  3.215000 181.300000 ;
        RECT  3.015000 181.505000  3.215000 181.705000 ;
        RECT  3.015000 181.910000  3.215000 182.110000 ;
        RECT  3.015000 182.315000  3.215000 182.515000 ;
        RECT  3.015000 182.720000  3.215000 182.920000 ;
        RECT  3.015000 183.125000  3.215000 183.325000 ;
        RECT  3.015000 183.530000  3.215000 183.730000 ;
        RECT  3.015000 183.935000  3.215000 184.135000 ;
        RECT  3.015000 184.340000  3.215000 184.540000 ;
        RECT  3.015000 184.745000  3.215000 184.945000 ;
        RECT  3.015000 185.150000  3.215000 185.350000 ;
        RECT  3.015000 185.555000  3.215000 185.755000 ;
        RECT  3.015000 185.960000  3.215000 186.160000 ;
        RECT  3.015000 186.365000  3.215000 186.565000 ;
        RECT  3.015000 186.770000  3.215000 186.970000 ;
        RECT  3.015000 187.175000  3.215000 187.375000 ;
        RECT  3.015000 187.580000  3.215000 187.780000 ;
        RECT  3.015000 187.985000  3.215000 188.185000 ;
        RECT  3.015000 188.390000  3.215000 188.590000 ;
        RECT  3.015000 188.795000  3.215000 188.995000 ;
        RECT  3.015000 189.200000  3.215000 189.400000 ;
        RECT  3.015000 189.605000  3.215000 189.805000 ;
        RECT  3.015000 190.010000  3.215000 190.210000 ;
        RECT  3.015000 190.415000  3.215000 190.615000 ;
        RECT  3.015000 190.820000  3.215000 191.020000 ;
        RECT  3.015000 191.225000  3.215000 191.425000 ;
        RECT  3.015000 191.630000  3.215000 191.830000 ;
        RECT  3.015000 192.035000  3.215000 192.235000 ;
        RECT  3.015000 192.440000  3.215000 192.640000 ;
        RECT  3.015000 192.845000  3.215000 193.045000 ;
        RECT  3.015000 193.250000  3.215000 193.450000 ;
        RECT  3.015000 193.655000  3.215000 193.855000 ;
        RECT  3.015000 194.060000  3.215000 194.260000 ;
        RECT  3.015000 194.465000  3.215000 194.665000 ;
        RECT  3.015000 194.870000  3.215000 195.070000 ;
        RECT  3.015000 195.275000  3.215000 195.475000 ;
        RECT  3.015000 195.680000  3.215000 195.880000 ;
        RECT  3.015000 196.085000  3.215000 196.285000 ;
        RECT  3.015000 196.490000  3.215000 196.690000 ;
        RECT  3.015000 196.895000  3.215000 197.095000 ;
        RECT  3.015000 197.300000  3.215000 197.500000 ;
        RECT  3.015000 197.705000  3.215000 197.905000 ;
        RECT  3.050000  23.910000  3.250000  24.110000 ;
        RECT  3.050000  24.340000  3.250000  24.540000 ;
        RECT  3.050000  24.770000  3.250000  24.970000 ;
        RECT  3.050000  25.200000  3.250000  25.400000 ;
        RECT  3.050000  25.630000  3.250000  25.830000 ;
        RECT  3.050000  26.060000  3.250000  26.260000 ;
        RECT  3.050000  26.490000  3.250000  26.690000 ;
        RECT  3.050000  26.920000  3.250000  27.120000 ;
        RECT  3.050000  27.350000  3.250000  27.550000 ;
        RECT  3.050000  27.780000  3.250000  27.980000 ;
        RECT  3.050000  28.210000  3.250000  28.410000 ;
        RECT  3.415000 173.900000  3.615000 174.100000 ;
        RECT  3.415000 174.300000  3.615000 174.500000 ;
        RECT  3.415000 174.700000  3.615000 174.900000 ;
        RECT  3.415000 175.100000  3.615000 175.300000 ;
        RECT  3.415000 175.500000  3.615000 175.700000 ;
        RECT  3.415000 175.900000  3.615000 176.100000 ;
        RECT  3.415000 176.300000  3.615000 176.500000 ;
        RECT  3.415000 176.700000  3.615000 176.900000 ;
        RECT  3.415000 177.100000  3.615000 177.300000 ;
        RECT  3.415000 177.500000  3.615000 177.700000 ;
        RECT  3.415000 177.900000  3.615000 178.100000 ;
        RECT  3.415000 178.300000  3.615000 178.500000 ;
        RECT  3.415000 178.700000  3.615000 178.900000 ;
        RECT  3.415000 179.100000  3.615000 179.300000 ;
        RECT  3.415000 179.500000  3.615000 179.700000 ;
        RECT  3.415000 179.900000  3.615000 180.100000 ;
        RECT  3.415000 180.300000  3.615000 180.500000 ;
        RECT  3.415000 180.700000  3.615000 180.900000 ;
        RECT  3.415000 181.100000  3.615000 181.300000 ;
        RECT  3.415000 181.505000  3.615000 181.705000 ;
        RECT  3.415000 181.910000  3.615000 182.110000 ;
        RECT  3.415000 182.315000  3.615000 182.515000 ;
        RECT  3.415000 182.720000  3.615000 182.920000 ;
        RECT  3.415000 183.125000  3.615000 183.325000 ;
        RECT  3.415000 183.530000  3.615000 183.730000 ;
        RECT  3.415000 183.935000  3.615000 184.135000 ;
        RECT  3.415000 184.340000  3.615000 184.540000 ;
        RECT  3.415000 184.745000  3.615000 184.945000 ;
        RECT  3.415000 185.150000  3.615000 185.350000 ;
        RECT  3.415000 185.555000  3.615000 185.755000 ;
        RECT  3.415000 185.960000  3.615000 186.160000 ;
        RECT  3.415000 186.365000  3.615000 186.565000 ;
        RECT  3.415000 186.770000  3.615000 186.970000 ;
        RECT  3.415000 187.175000  3.615000 187.375000 ;
        RECT  3.415000 187.580000  3.615000 187.780000 ;
        RECT  3.415000 187.985000  3.615000 188.185000 ;
        RECT  3.415000 188.390000  3.615000 188.590000 ;
        RECT  3.415000 188.795000  3.615000 188.995000 ;
        RECT  3.415000 189.200000  3.615000 189.400000 ;
        RECT  3.415000 189.605000  3.615000 189.805000 ;
        RECT  3.415000 190.010000  3.615000 190.210000 ;
        RECT  3.415000 190.415000  3.615000 190.615000 ;
        RECT  3.415000 190.820000  3.615000 191.020000 ;
        RECT  3.415000 191.225000  3.615000 191.425000 ;
        RECT  3.415000 191.630000  3.615000 191.830000 ;
        RECT  3.415000 192.035000  3.615000 192.235000 ;
        RECT  3.415000 192.440000  3.615000 192.640000 ;
        RECT  3.415000 192.845000  3.615000 193.045000 ;
        RECT  3.415000 193.250000  3.615000 193.450000 ;
        RECT  3.415000 193.655000  3.615000 193.855000 ;
        RECT  3.415000 194.060000  3.615000 194.260000 ;
        RECT  3.415000 194.465000  3.615000 194.665000 ;
        RECT  3.415000 194.870000  3.615000 195.070000 ;
        RECT  3.415000 195.275000  3.615000 195.475000 ;
        RECT  3.415000 195.680000  3.615000 195.880000 ;
        RECT  3.415000 196.085000  3.615000 196.285000 ;
        RECT  3.415000 196.490000  3.615000 196.690000 ;
        RECT  3.415000 196.895000  3.615000 197.095000 ;
        RECT  3.415000 197.300000  3.615000 197.500000 ;
        RECT  3.415000 197.705000  3.615000 197.905000 ;
        RECT  3.455000  23.910000  3.655000  24.110000 ;
        RECT  3.455000  24.340000  3.655000  24.540000 ;
        RECT  3.455000  24.770000  3.655000  24.970000 ;
        RECT  3.455000  25.200000  3.655000  25.400000 ;
        RECT  3.455000  25.630000  3.655000  25.830000 ;
        RECT  3.455000  26.060000  3.655000  26.260000 ;
        RECT  3.455000  26.490000  3.655000  26.690000 ;
        RECT  3.455000  26.920000  3.655000  27.120000 ;
        RECT  3.455000  27.350000  3.655000  27.550000 ;
        RECT  3.455000  27.780000  3.655000  27.980000 ;
        RECT  3.455000  28.210000  3.655000  28.410000 ;
        RECT  3.815000 173.900000  4.015000 174.100000 ;
        RECT  3.815000 174.300000  4.015000 174.500000 ;
        RECT  3.815000 174.700000  4.015000 174.900000 ;
        RECT  3.815000 175.100000  4.015000 175.300000 ;
        RECT  3.815000 175.500000  4.015000 175.700000 ;
        RECT  3.815000 175.900000  4.015000 176.100000 ;
        RECT  3.815000 176.300000  4.015000 176.500000 ;
        RECT  3.815000 176.700000  4.015000 176.900000 ;
        RECT  3.815000 177.100000  4.015000 177.300000 ;
        RECT  3.815000 177.500000  4.015000 177.700000 ;
        RECT  3.815000 177.900000  4.015000 178.100000 ;
        RECT  3.815000 178.300000  4.015000 178.500000 ;
        RECT  3.815000 178.700000  4.015000 178.900000 ;
        RECT  3.815000 179.100000  4.015000 179.300000 ;
        RECT  3.815000 179.500000  4.015000 179.700000 ;
        RECT  3.815000 179.900000  4.015000 180.100000 ;
        RECT  3.815000 180.300000  4.015000 180.500000 ;
        RECT  3.815000 180.700000  4.015000 180.900000 ;
        RECT  3.815000 181.100000  4.015000 181.300000 ;
        RECT  3.815000 181.505000  4.015000 181.705000 ;
        RECT  3.815000 181.910000  4.015000 182.110000 ;
        RECT  3.815000 182.315000  4.015000 182.515000 ;
        RECT  3.815000 182.720000  4.015000 182.920000 ;
        RECT  3.815000 183.125000  4.015000 183.325000 ;
        RECT  3.815000 183.530000  4.015000 183.730000 ;
        RECT  3.815000 183.935000  4.015000 184.135000 ;
        RECT  3.815000 184.340000  4.015000 184.540000 ;
        RECT  3.815000 184.745000  4.015000 184.945000 ;
        RECT  3.815000 185.150000  4.015000 185.350000 ;
        RECT  3.815000 185.555000  4.015000 185.755000 ;
        RECT  3.815000 185.960000  4.015000 186.160000 ;
        RECT  3.815000 186.365000  4.015000 186.565000 ;
        RECT  3.815000 186.770000  4.015000 186.970000 ;
        RECT  3.815000 187.175000  4.015000 187.375000 ;
        RECT  3.815000 187.580000  4.015000 187.780000 ;
        RECT  3.815000 187.985000  4.015000 188.185000 ;
        RECT  3.815000 188.390000  4.015000 188.590000 ;
        RECT  3.815000 188.795000  4.015000 188.995000 ;
        RECT  3.815000 189.200000  4.015000 189.400000 ;
        RECT  3.815000 189.605000  4.015000 189.805000 ;
        RECT  3.815000 190.010000  4.015000 190.210000 ;
        RECT  3.815000 190.415000  4.015000 190.615000 ;
        RECT  3.815000 190.820000  4.015000 191.020000 ;
        RECT  3.815000 191.225000  4.015000 191.425000 ;
        RECT  3.815000 191.630000  4.015000 191.830000 ;
        RECT  3.815000 192.035000  4.015000 192.235000 ;
        RECT  3.815000 192.440000  4.015000 192.640000 ;
        RECT  3.815000 192.845000  4.015000 193.045000 ;
        RECT  3.815000 193.250000  4.015000 193.450000 ;
        RECT  3.815000 193.655000  4.015000 193.855000 ;
        RECT  3.815000 194.060000  4.015000 194.260000 ;
        RECT  3.815000 194.465000  4.015000 194.665000 ;
        RECT  3.815000 194.870000  4.015000 195.070000 ;
        RECT  3.815000 195.275000  4.015000 195.475000 ;
        RECT  3.815000 195.680000  4.015000 195.880000 ;
        RECT  3.815000 196.085000  4.015000 196.285000 ;
        RECT  3.815000 196.490000  4.015000 196.690000 ;
        RECT  3.815000 196.895000  4.015000 197.095000 ;
        RECT  3.815000 197.300000  4.015000 197.500000 ;
        RECT  3.815000 197.705000  4.015000 197.905000 ;
        RECT  3.860000  23.910000  4.060000  24.110000 ;
        RECT  3.860000  24.340000  4.060000  24.540000 ;
        RECT  3.860000  24.770000  4.060000  24.970000 ;
        RECT  3.860000  25.200000  4.060000  25.400000 ;
        RECT  3.860000  25.630000  4.060000  25.830000 ;
        RECT  3.860000  26.060000  4.060000  26.260000 ;
        RECT  3.860000  26.490000  4.060000  26.690000 ;
        RECT  3.860000  26.920000  4.060000  27.120000 ;
        RECT  3.860000  27.350000  4.060000  27.550000 ;
        RECT  3.860000  27.780000  4.060000  27.980000 ;
        RECT  3.860000  28.210000  4.060000  28.410000 ;
        RECT  4.215000 173.900000  4.415000 174.100000 ;
        RECT  4.215000 174.300000  4.415000 174.500000 ;
        RECT  4.215000 174.700000  4.415000 174.900000 ;
        RECT  4.215000 175.100000  4.415000 175.300000 ;
        RECT  4.215000 175.500000  4.415000 175.700000 ;
        RECT  4.215000 175.900000  4.415000 176.100000 ;
        RECT  4.215000 176.300000  4.415000 176.500000 ;
        RECT  4.215000 176.700000  4.415000 176.900000 ;
        RECT  4.215000 177.100000  4.415000 177.300000 ;
        RECT  4.215000 177.500000  4.415000 177.700000 ;
        RECT  4.215000 177.900000  4.415000 178.100000 ;
        RECT  4.215000 178.300000  4.415000 178.500000 ;
        RECT  4.215000 178.700000  4.415000 178.900000 ;
        RECT  4.215000 179.100000  4.415000 179.300000 ;
        RECT  4.215000 179.500000  4.415000 179.700000 ;
        RECT  4.215000 179.900000  4.415000 180.100000 ;
        RECT  4.215000 180.300000  4.415000 180.500000 ;
        RECT  4.215000 180.700000  4.415000 180.900000 ;
        RECT  4.215000 181.100000  4.415000 181.300000 ;
        RECT  4.215000 181.505000  4.415000 181.705000 ;
        RECT  4.215000 181.910000  4.415000 182.110000 ;
        RECT  4.215000 182.315000  4.415000 182.515000 ;
        RECT  4.215000 182.720000  4.415000 182.920000 ;
        RECT  4.215000 183.125000  4.415000 183.325000 ;
        RECT  4.215000 183.530000  4.415000 183.730000 ;
        RECT  4.215000 183.935000  4.415000 184.135000 ;
        RECT  4.215000 184.340000  4.415000 184.540000 ;
        RECT  4.215000 184.745000  4.415000 184.945000 ;
        RECT  4.215000 185.150000  4.415000 185.350000 ;
        RECT  4.215000 185.555000  4.415000 185.755000 ;
        RECT  4.215000 185.960000  4.415000 186.160000 ;
        RECT  4.215000 186.365000  4.415000 186.565000 ;
        RECT  4.215000 186.770000  4.415000 186.970000 ;
        RECT  4.215000 187.175000  4.415000 187.375000 ;
        RECT  4.215000 187.580000  4.415000 187.780000 ;
        RECT  4.215000 187.985000  4.415000 188.185000 ;
        RECT  4.215000 188.390000  4.415000 188.590000 ;
        RECT  4.215000 188.795000  4.415000 188.995000 ;
        RECT  4.215000 189.200000  4.415000 189.400000 ;
        RECT  4.215000 189.605000  4.415000 189.805000 ;
        RECT  4.215000 190.010000  4.415000 190.210000 ;
        RECT  4.215000 190.415000  4.415000 190.615000 ;
        RECT  4.215000 190.820000  4.415000 191.020000 ;
        RECT  4.215000 191.225000  4.415000 191.425000 ;
        RECT  4.215000 191.630000  4.415000 191.830000 ;
        RECT  4.215000 192.035000  4.415000 192.235000 ;
        RECT  4.215000 192.440000  4.415000 192.640000 ;
        RECT  4.215000 192.845000  4.415000 193.045000 ;
        RECT  4.215000 193.250000  4.415000 193.450000 ;
        RECT  4.215000 193.655000  4.415000 193.855000 ;
        RECT  4.215000 194.060000  4.415000 194.260000 ;
        RECT  4.215000 194.465000  4.415000 194.665000 ;
        RECT  4.215000 194.870000  4.415000 195.070000 ;
        RECT  4.215000 195.275000  4.415000 195.475000 ;
        RECT  4.215000 195.680000  4.415000 195.880000 ;
        RECT  4.215000 196.085000  4.415000 196.285000 ;
        RECT  4.215000 196.490000  4.415000 196.690000 ;
        RECT  4.215000 196.895000  4.415000 197.095000 ;
        RECT  4.215000 197.300000  4.415000 197.500000 ;
        RECT  4.215000 197.705000  4.415000 197.905000 ;
        RECT  4.265000  23.910000  4.465000  24.110000 ;
        RECT  4.265000  24.340000  4.465000  24.540000 ;
        RECT  4.265000  24.770000  4.465000  24.970000 ;
        RECT  4.265000  25.200000  4.465000  25.400000 ;
        RECT  4.265000  25.630000  4.465000  25.830000 ;
        RECT  4.265000  26.060000  4.465000  26.260000 ;
        RECT  4.265000  26.490000  4.465000  26.690000 ;
        RECT  4.265000  26.920000  4.465000  27.120000 ;
        RECT  4.265000  27.350000  4.465000  27.550000 ;
        RECT  4.265000  27.780000  4.465000  27.980000 ;
        RECT  4.265000  28.210000  4.465000  28.410000 ;
        RECT  4.615000 173.900000  4.815000 174.100000 ;
        RECT  4.615000 174.300000  4.815000 174.500000 ;
        RECT  4.615000 174.700000  4.815000 174.900000 ;
        RECT  4.615000 175.100000  4.815000 175.300000 ;
        RECT  4.615000 175.500000  4.815000 175.700000 ;
        RECT  4.615000 175.900000  4.815000 176.100000 ;
        RECT  4.615000 176.300000  4.815000 176.500000 ;
        RECT  4.615000 176.700000  4.815000 176.900000 ;
        RECT  4.615000 177.100000  4.815000 177.300000 ;
        RECT  4.615000 177.500000  4.815000 177.700000 ;
        RECT  4.615000 177.900000  4.815000 178.100000 ;
        RECT  4.615000 178.300000  4.815000 178.500000 ;
        RECT  4.615000 178.700000  4.815000 178.900000 ;
        RECT  4.615000 179.100000  4.815000 179.300000 ;
        RECT  4.615000 179.500000  4.815000 179.700000 ;
        RECT  4.615000 179.900000  4.815000 180.100000 ;
        RECT  4.615000 180.300000  4.815000 180.500000 ;
        RECT  4.615000 180.700000  4.815000 180.900000 ;
        RECT  4.615000 181.100000  4.815000 181.300000 ;
        RECT  4.615000 181.505000  4.815000 181.705000 ;
        RECT  4.615000 181.910000  4.815000 182.110000 ;
        RECT  4.615000 182.315000  4.815000 182.515000 ;
        RECT  4.615000 182.720000  4.815000 182.920000 ;
        RECT  4.615000 183.125000  4.815000 183.325000 ;
        RECT  4.615000 183.530000  4.815000 183.730000 ;
        RECT  4.615000 183.935000  4.815000 184.135000 ;
        RECT  4.615000 184.340000  4.815000 184.540000 ;
        RECT  4.615000 184.745000  4.815000 184.945000 ;
        RECT  4.615000 185.150000  4.815000 185.350000 ;
        RECT  4.615000 185.555000  4.815000 185.755000 ;
        RECT  4.615000 185.960000  4.815000 186.160000 ;
        RECT  4.615000 186.365000  4.815000 186.565000 ;
        RECT  4.615000 186.770000  4.815000 186.970000 ;
        RECT  4.615000 187.175000  4.815000 187.375000 ;
        RECT  4.615000 187.580000  4.815000 187.780000 ;
        RECT  4.615000 187.985000  4.815000 188.185000 ;
        RECT  4.615000 188.390000  4.815000 188.590000 ;
        RECT  4.615000 188.795000  4.815000 188.995000 ;
        RECT  4.615000 189.200000  4.815000 189.400000 ;
        RECT  4.615000 189.605000  4.815000 189.805000 ;
        RECT  4.615000 190.010000  4.815000 190.210000 ;
        RECT  4.615000 190.415000  4.815000 190.615000 ;
        RECT  4.615000 190.820000  4.815000 191.020000 ;
        RECT  4.615000 191.225000  4.815000 191.425000 ;
        RECT  4.615000 191.630000  4.815000 191.830000 ;
        RECT  4.615000 192.035000  4.815000 192.235000 ;
        RECT  4.615000 192.440000  4.815000 192.640000 ;
        RECT  4.615000 192.845000  4.815000 193.045000 ;
        RECT  4.615000 193.250000  4.815000 193.450000 ;
        RECT  4.615000 193.655000  4.815000 193.855000 ;
        RECT  4.615000 194.060000  4.815000 194.260000 ;
        RECT  4.615000 194.465000  4.815000 194.665000 ;
        RECT  4.615000 194.870000  4.815000 195.070000 ;
        RECT  4.615000 195.275000  4.815000 195.475000 ;
        RECT  4.615000 195.680000  4.815000 195.880000 ;
        RECT  4.615000 196.085000  4.815000 196.285000 ;
        RECT  4.615000 196.490000  4.815000 196.690000 ;
        RECT  4.615000 196.895000  4.815000 197.095000 ;
        RECT  4.615000 197.300000  4.815000 197.500000 ;
        RECT  4.615000 197.705000  4.815000 197.905000 ;
        RECT  4.670000  23.910000  4.870000  24.110000 ;
        RECT  4.670000  24.340000  4.870000  24.540000 ;
        RECT  4.670000  24.770000  4.870000  24.970000 ;
        RECT  4.670000  25.200000  4.870000  25.400000 ;
        RECT  4.670000  25.630000  4.870000  25.830000 ;
        RECT  4.670000  26.060000  4.870000  26.260000 ;
        RECT  4.670000  26.490000  4.870000  26.690000 ;
        RECT  4.670000  26.920000  4.870000  27.120000 ;
        RECT  4.670000  27.350000  4.870000  27.550000 ;
        RECT  4.670000  27.780000  4.870000  27.980000 ;
        RECT  4.670000  28.210000  4.870000  28.410000 ;
        RECT  5.015000 173.900000  5.215000 174.100000 ;
        RECT  5.015000 174.300000  5.215000 174.500000 ;
        RECT  5.015000 174.700000  5.215000 174.900000 ;
        RECT  5.015000 175.100000  5.215000 175.300000 ;
        RECT  5.015000 175.500000  5.215000 175.700000 ;
        RECT  5.015000 175.900000  5.215000 176.100000 ;
        RECT  5.015000 176.300000  5.215000 176.500000 ;
        RECT  5.015000 176.700000  5.215000 176.900000 ;
        RECT  5.015000 177.100000  5.215000 177.300000 ;
        RECT  5.015000 177.500000  5.215000 177.700000 ;
        RECT  5.015000 177.900000  5.215000 178.100000 ;
        RECT  5.015000 178.300000  5.215000 178.500000 ;
        RECT  5.015000 178.700000  5.215000 178.900000 ;
        RECT  5.015000 179.100000  5.215000 179.300000 ;
        RECT  5.015000 179.500000  5.215000 179.700000 ;
        RECT  5.015000 179.900000  5.215000 180.100000 ;
        RECT  5.015000 180.300000  5.215000 180.500000 ;
        RECT  5.015000 180.700000  5.215000 180.900000 ;
        RECT  5.015000 181.100000  5.215000 181.300000 ;
        RECT  5.015000 181.505000  5.215000 181.705000 ;
        RECT  5.015000 181.910000  5.215000 182.110000 ;
        RECT  5.015000 182.315000  5.215000 182.515000 ;
        RECT  5.015000 182.720000  5.215000 182.920000 ;
        RECT  5.015000 183.125000  5.215000 183.325000 ;
        RECT  5.015000 183.530000  5.215000 183.730000 ;
        RECT  5.015000 183.935000  5.215000 184.135000 ;
        RECT  5.015000 184.340000  5.215000 184.540000 ;
        RECT  5.015000 184.745000  5.215000 184.945000 ;
        RECT  5.015000 185.150000  5.215000 185.350000 ;
        RECT  5.015000 185.555000  5.215000 185.755000 ;
        RECT  5.015000 185.960000  5.215000 186.160000 ;
        RECT  5.015000 186.365000  5.215000 186.565000 ;
        RECT  5.015000 186.770000  5.215000 186.970000 ;
        RECT  5.015000 187.175000  5.215000 187.375000 ;
        RECT  5.015000 187.580000  5.215000 187.780000 ;
        RECT  5.015000 187.985000  5.215000 188.185000 ;
        RECT  5.015000 188.390000  5.215000 188.590000 ;
        RECT  5.015000 188.795000  5.215000 188.995000 ;
        RECT  5.015000 189.200000  5.215000 189.400000 ;
        RECT  5.015000 189.605000  5.215000 189.805000 ;
        RECT  5.015000 190.010000  5.215000 190.210000 ;
        RECT  5.015000 190.415000  5.215000 190.615000 ;
        RECT  5.015000 190.820000  5.215000 191.020000 ;
        RECT  5.015000 191.225000  5.215000 191.425000 ;
        RECT  5.015000 191.630000  5.215000 191.830000 ;
        RECT  5.015000 192.035000  5.215000 192.235000 ;
        RECT  5.015000 192.440000  5.215000 192.640000 ;
        RECT  5.015000 192.845000  5.215000 193.045000 ;
        RECT  5.015000 193.250000  5.215000 193.450000 ;
        RECT  5.015000 193.655000  5.215000 193.855000 ;
        RECT  5.015000 194.060000  5.215000 194.260000 ;
        RECT  5.015000 194.465000  5.215000 194.665000 ;
        RECT  5.015000 194.870000  5.215000 195.070000 ;
        RECT  5.015000 195.275000  5.215000 195.475000 ;
        RECT  5.015000 195.680000  5.215000 195.880000 ;
        RECT  5.015000 196.085000  5.215000 196.285000 ;
        RECT  5.015000 196.490000  5.215000 196.690000 ;
        RECT  5.015000 196.895000  5.215000 197.095000 ;
        RECT  5.015000 197.300000  5.215000 197.500000 ;
        RECT  5.015000 197.705000  5.215000 197.905000 ;
        RECT  5.075000  23.910000  5.275000  24.110000 ;
        RECT  5.075000  24.340000  5.275000  24.540000 ;
        RECT  5.075000  24.770000  5.275000  24.970000 ;
        RECT  5.075000  25.200000  5.275000  25.400000 ;
        RECT  5.075000  25.630000  5.275000  25.830000 ;
        RECT  5.075000  26.060000  5.275000  26.260000 ;
        RECT  5.075000  26.490000  5.275000  26.690000 ;
        RECT  5.075000  26.920000  5.275000  27.120000 ;
        RECT  5.075000  27.350000  5.275000  27.550000 ;
        RECT  5.075000  27.780000  5.275000  27.980000 ;
        RECT  5.075000  28.210000  5.275000  28.410000 ;
        RECT  5.415000 173.900000  5.615000 174.100000 ;
        RECT  5.415000 174.300000  5.615000 174.500000 ;
        RECT  5.415000 174.700000  5.615000 174.900000 ;
        RECT  5.415000 175.100000  5.615000 175.300000 ;
        RECT  5.415000 175.500000  5.615000 175.700000 ;
        RECT  5.415000 175.900000  5.615000 176.100000 ;
        RECT  5.415000 176.300000  5.615000 176.500000 ;
        RECT  5.415000 176.700000  5.615000 176.900000 ;
        RECT  5.415000 177.100000  5.615000 177.300000 ;
        RECT  5.415000 177.500000  5.615000 177.700000 ;
        RECT  5.415000 177.900000  5.615000 178.100000 ;
        RECT  5.415000 178.300000  5.615000 178.500000 ;
        RECT  5.415000 178.700000  5.615000 178.900000 ;
        RECT  5.415000 179.100000  5.615000 179.300000 ;
        RECT  5.415000 179.500000  5.615000 179.700000 ;
        RECT  5.415000 179.900000  5.615000 180.100000 ;
        RECT  5.415000 180.300000  5.615000 180.500000 ;
        RECT  5.415000 180.700000  5.615000 180.900000 ;
        RECT  5.415000 181.100000  5.615000 181.300000 ;
        RECT  5.415000 181.505000  5.615000 181.705000 ;
        RECT  5.415000 181.910000  5.615000 182.110000 ;
        RECT  5.415000 182.315000  5.615000 182.515000 ;
        RECT  5.415000 182.720000  5.615000 182.920000 ;
        RECT  5.415000 183.125000  5.615000 183.325000 ;
        RECT  5.415000 183.530000  5.615000 183.730000 ;
        RECT  5.415000 183.935000  5.615000 184.135000 ;
        RECT  5.415000 184.340000  5.615000 184.540000 ;
        RECT  5.415000 184.745000  5.615000 184.945000 ;
        RECT  5.415000 185.150000  5.615000 185.350000 ;
        RECT  5.415000 185.555000  5.615000 185.755000 ;
        RECT  5.415000 185.960000  5.615000 186.160000 ;
        RECT  5.415000 186.365000  5.615000 186.565000 ;
        RECT  5.415000 186.770000  5.615000 186.970000 ;
        RECT  5.415000 187.175000  5.615000 187.375000 ;
        RECT  5.415000 187.580000  5.615000 187.780000 ;
        RECT  5.415000 187.985000  5.615000 188.185000 ;
        RECT  5.415000 188.390000  5.615000 188.590000 ;
        RECT  5.415000 188.795000  5.615000 188.995000 ;
        RECT  5.415000 189.200000  5.615000 189.400000 ;
        RECT  5.415000 189.605000  5.615000 189.805000 ;
        RECT  5.415000 190.010000  5.615000 190.210000 ;
        RECT  5.415000 190.415000  5.615000 190.615000 ;
        RECT  5.415000 190.820000  5.615000 191.020000 ;
        RECT  5.415000 191.225000  5.615000 191.425000 ;
        RECT  5.415000 191.630000  5.615000 191.830000 ;
        RECT  5.415000 192.035000  5.615000 192.235000 ;
        RECT  5.415000 192.440000  5.615000 192.640000 ;
        RECT  5.415000 192.845000  5.615000 193.045000 ;
        RECT  5.415000 193.250000  5.615000 193.450000 ;
        RECT  5.415000 193.655000  5.615000 193.855000 ;
        RECT  5.415000 194.060000  5.615000 194.260000 ;
        RECT  5.415000 194.465000  5.615000 194.665000 ;
        RECT  5.415000 194.870000  5.615000 195.070000 ;
        RECT  5.415000 195.275000  5.615000 195.475000 ;
        RECT  5.415000 195.680000  5.615000 195.880000 ;
        RECT  5.415000 196.085000  5.615000 196.285000 ;
        RECT  5.415000 196.490000  5.615000 196.690000 ;
        RECT  5.415000 196.895000  5.615000 197.095000 ;
        RECT  5.415000 197.300000  5.615000 197.500000 ;
        RECT  5.415000 197.705000  5.615000 197.905000 ;
        RECT  5.480000  23.910000  5.680000  24.110000 ;
        RECT  5.480000  24.340000  5.680000  24.540000 ;
        RECT  5.480000  24.770000  5.680000  24.970000 ;
        RECT  5.480000  25.200000  5.680000  25.400000 ;
        RECT  5.480000  25.630000  5.680000  25.830000 ;
        RECT  5.480000  26.060000  5.680000  26.260000 ;
        RECT  5.480000  26.490000  5.680000  26.690000 ;
        RECT  5.480000  26.920000  5.680000  27.120000 ;
        RECT  5.480000  27.350000  5.680000  27.550000 ;
        RECT  5.480000  27.780000  5.680000  27.980000 ;
        RECT  5.480000  28.210000  5.680000  28.410000 ;
        RECT  5.815000 173.900000  6.015000 174.100000 ;
        RECT  5.815000 174.300000  6.015000 174.500000 ;
        RECT  5.815000 174.700000  6.015000 174.900000 ;
        RECT  5.815000 175.100000  6.015000 175.300000 ;
        RECT  5.815000 175.500000  6.015000 175.700000 ;
        RECT  5.815000 175.900000  6.015000 176.100000 ;
        RECT  5.815000 176.300000  6.015000 176.500000 ;
        RECT  5.815000 176.700000  6.015000 176.900000 ;
        RECT  5.815000 177.100000  6.015000 177.300000 ;
        RECT  5.815000 177.500000  6.015000 177.700000 ;
        RECT  5.815000 177.900000  6.015000 178.100000 ;
        RECT  5.815000 178.300000  6.015000 178.500000 ;
        RECT  5.815000 178.700000  6.015000 178.900000 ;
        RECT  5.815000 179.100000  6.015000 179.300000 ;
        RECT  5.815000 179.500000  6.015000 179.700000 ;
        RECT  5.815000 179.900000  6.015000 180.100000 ;
        RECT  5.815000 180.300000  6.015000 180.500000 ;
        RECT  5.815000 180.700000  6.015000 180.900000 ;
        RECT  5.815000 181.100000  6.015000 181.300000 ;
        RECT  5.815000 181.505000  6.015000 181.705000 ;
        RECT  5.815000 181.910000  6.015000 182.110000 ;
        RECT  5.815000 182.315000  6.015000 182.515000 ;
        RECT  5.815000 182.720000  6.015000 182.920000 ;
        RECT  5.815000 183.125000  6.015000 183.325000 ;
        RECT  5.815000 183.530000  6.015000 183.730000 ;
        RECT  5.815000 183.935000  6.015000 184.135000 ;
        RECT  5.815000 184.340000  6.015000 184.540000 ;
        RECT  5.815000 184.745000  6.015000 184.945000 ;
        RECT  5.815000 185.150000  6.015000 185.350000 ;
        RECT  5.815000 185.555000  6.015000 185.755000 ;
        RECT  5.815000 185.960000  6.015000 186.160000 ;
        RECT  5.815000 186.365000  6.015000 186.565000 ;
        RECT  5.815000 186.770000  6.015000 186.970000 ;
        RECT  5.815000 187.175000  6.015000 187.375000 ;
        RECT  5.815000 187.580000  6.015000 187.780000 ;
        RECT  5.815000 187.985000  6.015000 188.185000 ;
        RECT  5.815000 188.390000  6.015000 188.590000 ;
        RECT  5.815000 188.795000  6.015000 188.995000 ;
        RECT  5.815000 189.200000  6.015000 189.400000 ;
        RECT  5.815000 189.605000  6.015000 189.805000 ;
        RECT  5.815000 190.010000  6.015000 190.210000 ;
        RECT  5.815000 190.415000  6.015000 190.615000 ;
        RECT  5.815000 190.820000  6.015000 191.020000 ;
        RECT  5.815000 191.225000  6.015000 191.425000 ;
        RECT  5.815000 191.630000  6.015000 191.830000 ;
        RECT  5.815000 192.035000  6.015000 192.235000 ;
        RECT  5.815000 192.440000  6.015000 192.640000 ;
        RECT  5.815000 192.845000  6.015000 193.045000 ;
        RECT  5.815000 193.250000  6.015000 193.450000 ;
        RECT  5.815000 193.655000  6.015000 193.855000 ;
        RECT  5.815000 194.060000  6.015000 194.260000 ;
        RECT  5.815000 194.465000  6.015000 194.665000 ;
        RECT  5.815000 194.870000  6.015000 195.070000 ;
        RECT  5.815000 195.275000  6.015000 195.475000 ;
        RECT  5.815000 195.680000  6.015000 195.880000 ;
        RECT  5.815000 196.085000  6.015000 196.285000 ;
        RECT  5.815000 196.490000  6.015000 196.690000 ;
        RECT  5.815000 196.895000  6.015000 197.095000 ;
        RECT  5.815000 197.300000  6.015000 197.500000 ;
        RECT  5.815000 197.705000  6.015000 197.905000 ;
        RECT  5.885000  23.910000  6.085000  24.110000 ;
        RECT  5.885000  24.340000  6.085000  24.540000 ;
        RECT  5.885000  24.770000  6.085000  24.970000 ;
        RECT  5.885000  25.200000  6.085000  25.400000 ;
        RECT  5.885000  25.630000  6.085000  25.830000 ;
        RECT  5.885000  26.060000  6.085000  26.260000 ;
        RECT  5.885000  26.490000  6.085000  26.690000 ;
        RECT  5.885000  26.920000  6.085000  27.120000 ;
        RECT  5.885000  27.350000  6.085000  27.550000 ;
        RECT  5.885000  27.780000  6.085000  27.980000 ;
        RECT  5.885000  28.210000  6.085000  28.410000 ;
        RECT  6.215000 173.900000  6.415000 174.100000 ;
        RECT  6.215000 174.300000  6.415000 174.500000 ;
        RECT  6.215000 174.700000  6.415000 174.900000 ;
        RECT  6.215000 175.100000  6.415000 175.300000 ;
        RECT  6.215000 175.500000  6.415000 175.700000 ;
        RECT  6.215000 175.900000  6.415000 176.100000 ;
        RECT  6.215000 176.300000  6.415000 176.500000 ;
        RECT  6.215000 176.700000  6.415000 176.900000 ;
        RECT  6.215000 177.100000  6.415000 177.300000 ;
        RECT  6.215000 177.500000  6.415000 177.700000 ;
        RECT  6.215000 177.900000  6.415000 178.100000 ;
        RECT  6.215000 178.300000  6.415000 178.500000 ;
        RECT  6.215000 178.700000  6.415000 178.900000 ;
        RECT  6.215000 179.100000  6.415000 179.300000 ;
        RECT  6.215000 179.500000  6.415000 179.700000 ;
        RECT  6.215000 179.900000  6.415000 180.100000 ;
        RECT  6.215000 180.300000  6.415000 180.500000 ;
        RECT  6.215000 180.700000  6.415000 180.900000 ;
        RECT  6.215000 181.100000  6.415000 181.300000 ;
        RECT  6.215000 181.505000  6.415000 181.705000 ;
        RECT  6.215000 181.910000  6.415000 182.110000 ;
        RECT  6.215000 182.315000  6.415000 182.515000 ;
        RECT  6.215000 182.720000  6.415000 182.920000 ;
        RECT  6.215000 183.125000  6.415000 183.325000 ;
        RECT  6.215000 183.530000  6.415000 183.730000 ;
        RECT  6.215000 183.935000  6.415000 184.135000 ;
        RECT  6.215000 184.340000  6.415000 184.540000 ;
        RECT  6.215000 184.745000  6.415000 184.945000 ;
        RECT  6.215000 185.150000  6.415000 185.350000 ;
        RECT  6.215000 185.555000  6.415000 185.755000 ;
        RECT  6.215000 185.960000  6.415000 186.160000 ;
        RECT  6.215000 186.365000  6.415000 186.565000 ;
        RECT  6.215000 186.770000  6.415000 186.970000 ;
        RECT  6.215000 187.175000  6.415000 187.375000 ;
        RECT  6.215000 187.580000  6.415000 187.780000 ;
        RECT  6.215000 187.985000  6.415000 188.185000 ;
        RECT  6.215000 188.390000  6.415000 188.590000 ;
        RECT  6.215000 188.795000  6.415000 188.995000 ;
        RECT  6.215000 189.200000  6.415000 189.400000 ;
        RECT  6.215000 189.605000  6.415000 189.805000 ;
        RECT  6.215000 190.010000  6.415000 190.210000 ;
        RECT  6.215000 190.415000  6.415000 190.615000 ;
        RECT  6.215000 190.820000  6.415000 191.020000 ;
        RECT  6.215000 191.225000  6.415000 191.425000 ;
        RECT  6.215000 191.630000  6.415000 191.830000 ;
        RECT  6.215000 192.035000  6.415000 192.235000 ;
        RECT  6.215000 192.440000  6.415000 192.640000 ;
        RECT  6.215000 192.845000  6.415000 193.045000 ;
        RECT  6.215000 193.250000  6.415000 193.450000 ;
        RECT  6.215000 193.655000  6.415000 193.855000 ;
        RECT  6.215000 194.060000  6.415000 194.260000 ;
        RECT  6.215000 194.465000  6.415000 194.665000 ;
        RECT  6.215000 194.870000  6.415000 195.070000 ;
        RECT  6.215000 195.275000  6.415000 195.475000 ;
        RECT  6.215000 195.680000  6.415000 195.880000 ;
        RECT  6.215000 196.085000  6.415000 196.285000 ;
        RECT  6.215000 196.490000  6.415000 196.690000 ;
        RECT  6.215000 196.895000  6.415000 197.095000 ;
        RECT  6.215000 197.300000  6.415000 197.500000 ;
        RECT  6.215000 197.705000  6.415000 197.905000 ;
        RECT  6.290000  23.910000  6.490000  24.110000 ;
        RECT  6.290000  24.340000  6.490000  24.540000 ;
        RECT  6.290000  24.770000  6.490000  24.970000 ;
        RECT  6.290000  25.200000  6.490000  25.400000 ;
        RECT  6.290000  25.630000  6.490000  25.830000 ;
        RECT  6.290000  26.060000  6.490000  26.260000 ;
        RECT  6.290000  26.490000  6.490000  26.690000 ;
        RECT  6.290000  26.920000  6.490000  27.120000 ;
        RECT  6.290000  27.350000  6.490000  27.550000 ;
        RECT  6.290000  27.780000  6.490000  27.980000 ;
        RECT  6.290000  28.210000  6.490000  28.410000 ;
        RECT  6.615000 173.900000  6.815000 174.100000 ;
        RECT  6.615000 174.300000  6.815000 174.500000 ;
        RECT  6.615000 174.700000  6.815000 174.900000 ;
        RECT  6.615000 175.100000  6.815000 175.300000 ;
        RECT  6.615000 175.500000  6.815000 175.700000 ;
        RECT  6.615000 175.900000  6.815000 176.100000 ;
        RECT  6.615000 176.300000  6.815000 176.500000 ;
        RECT  6.615000 176.700000  6.815000 176.900000 ;
        RECT  6.615000 177.100000  6.815000 177.300000 ;
        RECT  6.615000 177.500000  6.815000 177.700000 ;
        RECT  6.615000 177.900000  6.815000 178.100000 ;
        RECT  6.615000 178.300000  6.815000 178.500000 ;
        RECT  6.615000 178.700000  6.815000 178.900000 ;
        RECT  6.615000 179.100000  6.815000 179.300000 ;
        RECT  6.615000 179.500000  6.815000 179.700000 ;
        RECT  6.615000 179.900000  6.815000 180.100000 ;
        RECT  6.615000 180.300000  6.815000 180.500000 ;
        RECT  6.615000 180.700000  6.815000 180.900000 ;
        RECT  6.615000 181.100000  6.815000 181.300000 ;
        RECT  6.615000 181.505000  6.815000 181.705000 ;
        RECT  6.615000 181.910000  6.815000 182.110000 ;
        RECT  6.615000 182.315000  6.815000 182.515000 ;
        RECT  6.615000 182.720000  6.815000 182.920000 ;
        RECT  6.615000 183.125000  6.815000 183.325000 ;
        RECT  6.615000 183.530000  6.815000 183.730000 ;
        RECT  6.615000 183.935000  6.815000 184.135000 ;
        RECT  6.615000 184.340000  6.815000 184.540000 ;
        RECT  6.615000 184.745000  6.815000 184.945000 ;
        RECT  6.615000 185.150000  6.815000 185.350000 ;
        RECT  6.615000 185.555000  6.815000 185.755000 ;
        RECT  6.615000 185.960000  6.815000 186.160000 ;
        RECT  6.615000 186.365000  6.815000 186.565000 ;
        RECT  6.615000 186.770000  6.815000 186.970000 ;
        RECT  6.615000 187.175000  6.815000 187.375000 ;
        RECT  6.615000 187.580000  6.815000 187.780000 ;
        RECT  6.615000 187.985000  6.815000 188.185000 ;
        RECT  6.615000 188.390000  6.815000 188.590000 ;
        RECT  6.615000 188.795000  6.815000 188.995000 ;
        RECT  6.615000 189.200000  6.815000 189.400000 ;
        RECT  6.615000 189.605000  6.815000 189.805000 ;
        RECT  6.615000 190.010000  6.815000 190.210000 ;
        RECT  6.615000 190.415000  6.815000 190.615000 ;
        RECT  6.615000 190.820000  6.815000 191.020000 ;
        RECT  6.615000 191.225000  6.815000 191.425000 ;
        RECT  6.615000 191.630000  6.815000 191.830000 ;
        RECT  6.615000 192.035000  6.815000 192.235000 ;
        RECT  6.615000 192.440000  6.815000 192.640000 ;
        RECT  6.615000 192.845000  6.815000 193.045000 ;
        RECT  6.615000 193.250000  6.815000 193.450000 ;
        RECT  6.615000 193.655000  6.815000 193.855000 ;
        RECT  6.615000 194.060000  6.815000 194.260000 ;
        RECT  6.615000 194.465000  6.815000 194.665000 ;
        RECT  6.615000 194.870000  6.815000 195.070000 ;
        RECT  6.615000 195.275000  6.815000 195.475000 ;
        RECT  6.615000 195.680000  6.815000 195.880000 ;
        RECT  6.615000 196.085000  6.815000 196.285000 ;
        RECT  6.615000 196.490000  6.815000 196.690000 ;
        RECT  6.615000 196.895000  6.815000 197.095000 ;
        RECT  6.615000 197.300000  6.815000 197.500000 ;
        RECT  6.615000 197.705000  6.815000 197.905000 ;
        RECT  6.695000  23.910000  6.895000  24.110000 ;
        RECT  6.695000  24.340000  6.895000  24.540000 ;
        RECT  6.695000  24.770000  6.895000  24.970000 ;
        RECT  6.695000  25.200000  6.895000  25.400000 ;
        RECT  6.695000  25.630000  6.895000  25.830000 ;
        RECT  6.695000  26.060000  6.895000  26.260000 ;
        RECT  6.695000  26.490000  6.895000  26.690000 ;
        RECT  6.695000  26.920000  6.895000  27.120000 ;
        RECT  6.695000  27.350000  6.895000  27.550000 ;
        RECT  6.695000  27.780000  6.895000  27.980000 ;
        RECT  6.695000  28.210000  6.895000  28.410000 ;
        RECT  7.015000 173.900000  7.215000 174.100000 ;
        RECT  7.015000 174.300000  7.215000 174.500000 ;
        RECT  7.015000 174.700000  7.215000 174.900000 ;
        RECT  7.015000 175.100000  7.215000 175.300000 ;
        RECT  7.015000 175.500000  7.215000 175.700000 ;
        RECT  7.015000 175.900000  7.215000 176.100000 ;
        RECT  7.015000 176.300000  7.215000 176.500000 ;
        RECT  7.015000 176.700000  7.215000 176.900000 ;
        RECT  7.015000 177.100000  7.215000 177.300000 ;
        RECT  7.015000 177.500000  7.215000 177.700000 ;
        RECT  7.015000 177.900000  7.215000 178.100000 ;
        RECT  7.015000 178.300000  7.215000 178.500000 ;
        RECT  7.015000 178.700000  7.215000 178.900000 ;
        RECT  7.015000 179.100000  7.215000 179.300000 ;
        RECT  7.015000 179.500000  7.215000 179.700000 ;
        RECT  7.015000 179.900000  7.215000 180.100000 ;
        RECT  7.015000 180.300000  7.215000 180.500000 ;
        RECT  7.015000 180.700000  7.215000 180.900000 ;
        RECT  7.015000 181.100000  7.215000 181.300000 ;
        RECT  7.015000 181.505000  7.215000 181.705000 ;
        RECT  7.015000 181.910000  7.215000 182.110000 ;
        RECT  7.015000 182.315000  7.215000 182.515000 ;
        RECT  7.015000 182.720000  7.215000 182.920000 ;
        RECT  7.015000 183.125000  7.215000 183.325000 ;
        RECT  7.015000 183.530000  7.215000 183.730000 ;
        RECT  7.015000 183.935000  7.215000 184.135000 ;
        RECT  7.015000 184.340000  7.215000 184.540000 ;
        RECT  7.015000 184.745000  7.215000 184.945000 ;
        RECT  7.015000 185.150000  7.215000 185.350000 ;
        RECT  7.015000 185.555000  7.215000 185.755000 ;
        RECT  7.015000 185.960000  7.215000 186.160000 ;
        RECT  7.015000 186.365000  7.215000 186.565000 ;
        RECT  7.015000 186.770000  7.215000 186.970000 ;
        RECT  7.015000 187.175000  7.215000 187.375000 ;
        RECT  7.015000 187.580000  7.215000 187.780000 ;
        RECT  7.015000 187.985000  7.215000 188.185000 ;
        RECT  7.015000 188.390000  7.215000 188.590000 ;
        RECT  7.015000 188.795000  7.215000 188.995000 ;
        RECT  7.015000 189.200000  7.215000 189.400000 ;
        RECT  7.015000 189.605000  7.215000 189.805000 ;
        RECT  7.015000 190.010000  7.215000 190.210000 ;
        RECT  7.015000 190.415000  7.215000 190.615000 ;
        RECT  7.015000 190.820000  7.215000 191.020000 ;
        RECT  7.015000 191.225000  7.215000 191.425000 ;
        RECT  7.015000 191.630000  7.215000 191.830000 ;
        RECT  7.015000 192.035000  7.215000 192.235000 ;
        RECT  7.015000 192.440000  7.215000 192.640000 ;
        RECT  7.015000 192.845000  7.215000 193.045000 ;
        RECT  7.015000 193.250000  7.215000 193.450000 ;
        RECT  7.015000 193.655000  7.215000 193.855000 ;
        RECT  7.015000 194.060000  7.215000 194.260000 ;
        RECT  7.015000 194.465000  7.215000 194.665000 ;
        RECT  7.015000 194.870000  7.215000 195.070000 ;
        RECT  7.015000 195.275000  7.215000 195.475000 ;
        RECT  7.015000 195.680000  7.215000 195.880000 ;
        RECT  7.015000 196.085000  7.215000 196.285000 ;
        RECT  7.015000 196.490000  7.215000 196.690000 ;
        RECT  7.015000 196.895000  7.215000 197.095000 ;
        RECT  7.015000 197.300000  7.215000 197.500000 ;
        RECT  7.015000 197.705000  7.215000 197.905000 ;
        RECT  7.100000  23.910000  7.300000  24.110000 ;
        RECT  7.100000  24.340000  7.300000  24.540000 ;
        RECT  7.100000  24.770000  7.300000  24.970000 ;
        RECT  7.100000  25.200000  7.300000  25.400000 ;
        RECT  7.100000  25.630000  7.300000  25.830000 ;
        RECT  7.100000  26.060000  7.300000  26.260000 ;
        RECT  7.100000  26.490000  7.300000  26.690000 ;
        RECT  7.100000  26.920000  7.300000  27.120000 ;
        RECT  7.100000  27.350000  7.300000  27.550000 ;
        RECT  7.100000  27.780000  7.300000  27.980000 ;
        RECT  7.100000  28.210000  7.300000  28.410000 ;
        RECT  7.415000 173.900000  7.615000 174.100000 ;
        RECT  7.415000 174.300000  7.615000 174.500000 ;
        RECT  7.415000 174.700000  7.615000 174.900000 ;
        RECT  7.415000 175.100000  7.615000 175.300000 ;
        RECT  7.415000 175.500000  7.615000 175.700000 ;
        RECT  7.415000 175.900000  7.615000 176.100000 ;
        RECT  7.415000 176.300000  7.615000 176.500000 ;
        RECT  7.415000 176.700000  7.615000 176.900000 ;
        RECT  7.415000 177.100000  7.615000 177.300000 ;
        RECT  7.415000 177.500000  7.615000 177.700000 ;
        RECT  7.415000 177.900000  7.615000 178.100000 ;
        RECT  7.415000 178.300000  7.615000 178.500000 ;
        RECT  7.415000 178.700000  7.615000 178.900000 ;
        RECT  7.415000 179.100000  7.615000 179.300000 ;
        RECT  7.415000 179.500000  7.615000 179.700000 ;
        RECT  7.415000 179.900000  7.615000 180.100000 ;
        RECT  7.415000 180.300000  7.615000 180.500000 ;
        RECT  7.415000 180.700000  7.615000 180.900000 ;
        RECT  7.415000 181.100000  7.615000 181.300000 ;
        RECT  7.415000 181.505000  7.615000 181.705000 ;
        RECT  7.415000 181.910000  7.615000 182.110000 ;
        RECT  7.415000 182.315000  7.615000 182.515000 ;
        RECT  7.415000 182.720000  7.615000 182.920000 ;
        RECT  7.415000 183.125000  7.615000 183.325000 ;
        RECT  7.415000 183.530000  7.615000 183.730000 ;
        RECT  7.415000 183.935000  7.615000 184.135000 ;
        RECT  7.415000 184.340000  7.615000 184.540000 ;
        RECT  7.415000 184.745000  7.615000 184.945000 ;
        RECT  7.415000 185.150000  7.615000 185.350000 ;
        RECT  7.415000 185.555000  7.615000 185.755000 ;
        RECT  7.415000 185.960000  7.615000 186.160000 ;
        RECT  7.415000 186.365000  7.615000 186.565000 ;
        RECT  7.415000 186.770000  7.615000 186.970000 ;
        RECT  7.415000 187.175000  7.615000 187.375000 ;
        RECT  7.415000 187.580000  7.615000 187.780000 ;
        RECT  7.415000 187.985000  7.615000 188.185000 ;
        RECT  7.415000 188.390000  7.615000 188.590000 ;
        RECT  7.415000 188.795000  7.615000 188.995000 ;
        RECT  7.415000 189.200000  7.615000 189.400000 ;
        RECT  7.415000 189.605000  7.615000 189.805000 ;
        RECT  7.415000 190.010000  7.615000 190.210000 ;
        RECT  7.415000 190.415000  7.615000 190.615000 ;
        RECT  7.415000 190.820000  7.615000 191.020000 ;
        RECT  7.415000 191.225000  7.615000 191.425000 ;
        RECT  7.415000 191.630000  7.615000 191.830000 ;
        RECT  7.415000 192.035000  7.615000 192.235000 ;
        RECT  7.415000 192.440000  7.615000 192.640000 ;
        RECT  7.415000 192.845000  7.615000 193.045000 ;
        RECT  7.415000 193.250000  7.615000 193.450000 ;
        RECT  7.415000 193.655000  7.615000 193.855000 ;
        RECT  7.415000 194.060000  7.615000 194.260000 ;
        RECT  7.415000 194.465000  7.615000 194.665000 ;
        RECT  7.415000 194.870000  7.615000 195.070000 ;
        RECT  7.415000 195.275000  7.615000 195.475000 ;
        RECT  7.415000 195.680000  7.615000 195.880000 ;
        RECT  7.415000 196.085000  7.615000 196.285000 ;
        RECT  7.415000 196.490000  7.615000 196.690000 ;
        RECT  7.415000 196.895000  7.615000 197.095000 ;
        RECT  7.415000 197.300000  7.615000 197.500000 ;
        RECT  7.415000 197.705000  7.615000 197.905000 ;
        RECT  7.505000  23.910000  7.705000  24.110000 ;
        RECT  7.505000  24.340000  7.705000  24.540000 ;
        RECT  7.505000  24.770000  7.705000  24.970000 ;
        RECT  7.505000  25.200000  7.705000  25.400000 ;
        RECT  7.505000  25.630000  7.705000  25.830000 ;
        RECT  7.505000  26.060000  7.705000  26.260000 ;
        RECT  7.505000  26.490000  7.705000  26.690000 ;
        RECT  7.505000  26.920000  7.705000  27.120000 ;
        RECT  7.505000  27.350000  7.705000  27.550000 ;
        RECT  7.505000  27.780000  7.705000  27.980000 ;
        RECT  7.505000  28.210000  7.705000  28.410000 ;
        RECT  7.815000 173.900000  8.015000 174.100000 ;
        RECT  7.815000 174.300000  8.015000 174.500000 ;
        RECT  7.815000 174.700000  8.015000 174.900000 ;
        RECT  7.815000 175.100000  8.015000 175.300000 ;
        RECT  7.815000 175.500000  8.015000 175.700000 ;
        RECT  7.815000 175.900000  8.015000 176.100000 ;
        RECT  7.815000 176.300000  8.015000 176.500000 ;
        RECT  7.815000 176.700000  8.015000 176.900000 ;
        RECT  7.815000 177.100000  8.015000 177.300000 ;
        RECT  7.815000 177.500000  8.015000 177.700000 ;
        RECT  7.815000 177.900000  8.015000 178.100000 ;
        RECT  7.815000 178.300000  8.015000 178.500000 ;
        RECT  7.815000 178.700000  8.015000 178.900000 ;
        RECT  7.815000 179.100000  8.015000 179.300000 ;
        RECT  7.815000 179.500000  8.015000 179.700000 ;
        RECT  7.815000 179.900000  8.015000 180.100000 ;
        RECT  7.815000 180.300000  8.015000 180.500000 ;
        RECT  7.815000 180.700000  8.015000 180.900000 ;
        RECT  7.815000 181.100000  8.015000 181.300000 ;
        RECT  7.815000 181.505000  8.015000 181.705000 ;
        RECT  7.815000 181.910000  8.015000 182.110000 ;
        RECT  7.815000 182.315000  8.015000 182.515000 ;
        RECT  7.815000 182.720000  8.015000 182.920000 ;
        RECT  7.815000 183.125000  8.015000 183.325000 ;
        RECT  7.815000 183.530000  8.015000 183.730000 ;
        RECT  7.815000 183.935000  8.015000 184.135000 ;
        RECT  7.815000 184.340000  8.015000 184.540000 ;
        RECT  7.815000 184.745000  8.015000 184.945000 ;
        RECT  7.815000 185.150000  8.015000 185.350000 ;
        RECT  7.815000 185.555000  8.015000 185.755000 ;
        RECT  7.815000 185.960000  8.015000 186.160000 ;
        RECT  7.815000 186.365000  8.015000 186.565000 ;
        RECT  7.815000 186.770000  8.015000 186.970000 ;
        RECT  7.815000 187.175000  8.015000 187.375000 ;
        RECT  7.815000 187.580000  8.015000 187.780000 ;
        RECT  7.815000 187.985000  8.015000 188.185000 ;
        RECT  7.815000 188.390000  8.015000 188.590000 ;
        RECT  7.815000 188.795000  8.015000 188.995000 ;
        RECT  7.815000 189.200000  8.015000 189.400000 ;
        RECT  7.815000 189.605000  8.015000 189.805000 ;
        RECT  7.815000 190.010000  8.015000 190.210000 ;
        RECT  7.815000 190.415000  8.015000 190.615000 ;
        RECT  7.815000 190.820000  8.015000 191.020000 ;
        RECT  7.815000 191.225000  8.015000 191.425000 ;
        RECT  7.815000 191.630000  8.015000 191.830000 ;
        RECT  7.815000 192.035000  8.015000 192.235000 ;
        RECT  7.815000 192.440000  8.015000 192.640000 ;
        RECT  7.815000 192.845000  8.015000 193.045000 ;
        RECT  7.815000 193.250000  8.015000 193.450000 ;
        RECT  7.815000 193.655000  8.015000 193.855000 ;
        RECT  7.815000 194.060000  8.015000 194.260000 ;
        RECT  7.815000 194.465000  8.015000 194.665000 ;
        RECT  7.815000 194.870000  8.015000 195.070000 ;
        RECT  7.815000 195.275000  8.015000 195.475000 ;
        RECT  7.815000 195.680000  8.015000 195.880000 ;
        RECT  7.815000 196.085000  8.015000 196.285000 ;
        RECT  7.815000 196.490000  8.015000 196.690000 ;
        RECT  7.815000 196.895000  8.015000 197.095000 ;
        RECT  7.815000 197.300000  8.015000 197.500000 ;
        RECT  7.815000 197.705000  8.015000 197.905000 ;
        RECT  7.910000  23.910000  8.110000  24.110000 ;
        RECT  7.910000  24.340000  8.110000  24.540000 ;
        RECT  7.910000  24.770000  8.110000  24.970000 ;
        RECT  7.910000  25.200000  8.110000  25.400000 ;
        RECT  7.910000  25.630000  8.110000  25.830000 ;
        RECT  7.910000  26.060000  8.110000  26.260000 ;
        RECT  7.910000  26.490000  8.110000  26.690000 ;
        RECT  7.910000  26.920000  8.110000  27.120000 ;
        RECT  7.910000  27.350000  8.110000  27.550000 ;
        RECT  7.910000  27.780000  8.110000  27.980000 ;
        RECT  7.910000  28.210000  8.110000  28.410000 ;
        RECT  8.215000 173.900000  8.415000 174.100000 ;
        RECT  8.215000 174.300000  8.415000 174.500000 ;
        RECT  8.215000 174.700000  8.415000 174.900000 ;
        RECT  8.215000 175.100000  8.415000 175.300000 ;
        RECT  8.215000 175.500000  8.415000 175.700000 ;
        RECT  8.215000 175.900000  8.415000 176.100000 ;
        RECT  8.215000 176.300000  8.415000 176.500000 ;
        RECT  8.215000 176.700000  8.415000 176.900000 ;
        RECT  8.215000 177.100000  8.415000 177.300000 ;
        RECT  8.215000 177.500000  8.415000 177.700000 ;
        RECT  8.215000 177.900000  8.415000 178.100000 ;
        RECT  8.215000 178.300000  8.415000 178.500000 ;
        RECT  8.215000 178.700000  8.415000 178.900000 ;
        RECT  8.215000 179.100000  8.415000 179.300000 ;
        RECT  8.215000 179.500000  8.415000 179.700000 ;
        RECT  8.215000 179.900000  8.415000 180.100000 ;
        RECT  8.215000 180.300000  8.415000 180.500000 ;
        RECT  8.215000 180.700000  8.415000 180.900000 ;
        RECT  8.215000 181.100000  8.415000 181.300000 ;
        RECT  8.215000 181.505000  8.415000 181.705000 ;
        RECT  8.215000 181.910000  8.415000 182.110000 ;
        RECT  8.215000 182.315000  8.415000 182.515000 ;
        RECT  8.215000 182.720000  8.415000 182.920000 ;
        RECT  8.215000 183.125000  8.415000 183.325000 ;
        RECT  8.215000 183.530000  8.415000 183.730000 ;
        RECT  8.215000 183.935000  8.415000 184.135000 ;
        RECT  8.215000 184.340000  8.415000 184.540000 ;
        RECT  8.215000 184.745000  8.415000 184.945000 ;
        RECT  8.215000 185.150000  8.415000 185.350000 ;
        RECT  8.215000 185.555000  8.415000 185.755000 ;
        RECT  8.215000 185.960000  8.415000 186.160000 ;
        RECT  8.215000 186.365000  8.415000 186.565000 ;
        RECT  8.215000 186.770000  8.415000 186.970000 ;
        RECT  8.215000 187.175000  8.415000 187.375000 ;
        RECT  8.215000 187.580000  8.415000 187.780000 ;
        RECT  8.215000 187.985000  8.415000 188.185000 ;
        RECT  8.215000 188.390000  8.415000 188.590000 ;
        RECT  8.215000 188.795000  8.415000 188.995000 ;
        RECT  8.215000 189.200000  8.415000 189.400000 ;
        RECT  8.215000 189.605000  8.415000 189.805000 ;
        RECT  8.215000 190.010000  8.415000 190.210000 ;
        RECT  8.215000 190.415000  8.415000 190.615000 ;
        RECT  8.215000 190.820000  8.415000 191.020000 ;
        RECT  8.215000 191.225000  8.415000 191.425000 ;
        RECT  8.215000 191.630000  8.415000 191.830000 ;
        RECT  8.215000 192.035000  8.415000 192.235000 ;
        RECT  8.215000 192.440000  8.415000 192.640000 ;
        RECT  8.215000 192.845000  8.415000 193.045000 ;
        RECT  8.215000 193.250000  8.415000 193.450000 ;
        RECT  8.215000 193.655000  8.415000 193.855000 ;
        RECT  8.215000 194.060000  8.415000 194.260000 ;
        RECT  8.215000 194.465000  8.415000 194.665000 ;
        RECT  8.215000 194.870000  8.415000 195.070000 ;
        RECT  8.215000 195.275000  8.415000 195.475000 ;
        RECT  8.215000 195.680000  8.415000 195.880000 ;
        RECT  8.215000 196.085000  8.415000 196.285000 ;
        RECT  8.215000 196.490000  8.415000 196.690000 ;
        RECT  8.215000 196.895000  8.415000 197.095000 ;
        RECT  8.215000 197.300000  8.415000 197.500000 ;
        RECT  8.215000 197.705000  8.415000 197.905000 ;
        RECT  8.315000  23.910000  8.515000  24.110000 ;
        RECT  8.315000  24.340000  8.515000  24.540000 ;
        RECT  8.315000  24.770000  8.515000  24.970000 ;
        RECT  8.315000  25.200000  8.515000  25.400000 ;
        RECT  8.315000  25.630000  8.515000  25.830000 ;
        RECT  8.315000  26.060000  8.515000  26.260000 ;
        RECT  8.315000  26.490000  8.515000  26.690000 ;
        RECT  8.315000  26.920000  8.515000  27.120000 ;
        RECT  8.315000  27.350000  8.515000  27.550000 ;
        RECT  8.315000  27.780000  8.515000  27.980000 ;
        RECT  8.315000  28.210000  8.515000  28.410000 ;
        RECT  8.615000 173.900000  8.815000 174.100000 ;
        RECT  8.615000 174.300000  8.815000 174.500000 ;
        RECT  8.615000 174.700000  8.815000 174.900000 ;
        RECT  8.615000 175.100000  8.815000 175.300000 ;
        RECT  8.615000 175.500000  8.815000 175.700000 ;
        RECT  8.615000 175.900000  8.815000 176.100000 ;
        RECT  8.615000 176.300000  8.815000 176.500000 ;
        RECT  8.615000 176.700000  8.815000 176.900000 ;
        RECT  8.615000 177.100000  8.815000 177.300000 ;
        RECT  8.615000 177.500000  8.815000 177.700000 ;
        RECT  8.615000 177.900000  8.815000 178.100000 ;
        RECT  8.615000 178.300000  8.815000 178.500000 ;
        RECT  8.615000 178.700000  8.815000 178.900000 ;
        RECT  8.615000 179.100000  8.815000 179.300000 ;
        RECT  8.615000 179.500000  8.815000 179.700000 ;
        RECT  8.615000 179.900000  8.815000 180.100000 ;
        RECT  8.615000 180.300000  8.815000 180.500000 ;
        RECT  8.615000 180.700000  8.815000 180.900000 ;
        RECT  8.615000 181.100000  8.815000 181.300000 ;
        RECT  8.615000 181.505000  8.815000 181.705000 ;
        RECT  8.615000 181.910000  8.815000 182.110000 ;
        RECT  8.615000 182.315000  8.815000 182.515000 ;
        RECT  8.615000 182.720000  8.815000 182.920000 ;
        RECT  8.615000 183.125000  8.815000 183.325000 ;
        RECT  8.615000 183.530000  8.815000 183.730000 ;
        RECT  8.615000 183.935000  8.815000 184.135000 ;
        RECT  8.615000 184.340000  8.815000 184.540000 ;
        RECT  8.615000 184.745000  8.815000 184.945000 ;
        RECT  8.615000 185.150000  8.815000 185.350000 ;
        RECT  8.615000 185.555000  8.815000 185.755000 ;
        RECT  8.615000 185.960000  8.815000 186.160000 ;
        RECT  8.615000 186.365000  8.815000 186.565000 ;
        RECT  8.615000 186.770000  8.815000 186.970000 ;
        RECT  8.615000 187.175000  8.815000 187.375000 ;
        RECT  8.615000 187.580000  8.815000 187.780000 ;
        RECT  8.615000 187.985000  8.815000 188.185000 ;
        RECT  8.615000 188.390000  8.815000 188.590000 ;
        RECT  8.615000 188.795000  8.815000 188.995000 ;
        RECT  8.615000 189.200000  8.815000 189.400000 ;
        RECT  8.615000 189.605000  8.815000 189.805000 ;
        RECT  8.615000 190.010000  8.815000 190.210000 ;
        RECT  8.615000 190.415000  8.815000 190.615000 ;
        RECT  8.615000 190.820000  8.815000 191.020000 ;
        RECT  8.615000 191.225000  8.815000 191.425000 ;
        RECT  8.615000 191.630000  8.815000 191.830000 ;
        RECT  8.615000 192.035000  8.815000 192.235000 ;
        RECT  8.615000 192.440000  8.815000 192.640000 ;
        RECT  8.615000 192.845000  8.815000 193.045000 ;
        RECT  8.615000 193.250000  8.815000 193.450000 ;
        RECT  8.615000 193.655000  8.815000 193.855000 ;
        RECT  8.615000 194.060000  8.815000 194.260000 ;
        RECT  8.615000 194.465000  8.815000 194.665000 ;
        RECT  8.615000 194.870000  8.815000 195.070000 ;
        RECT  8.615000 195.275000  8.815000 195.475000 ;
        RECT  8.615000 195.680000  8.815000 195.880000 ;
        RECT  8.615000 196.085000  8.815000 196.285000 ;
        RECT  8.615000 196.490000  8.815000 196.690000 ;
        RECT  8.615000 196.895000  8.815000 197.095000 ;
        RECT  8.615000 197.300000  8.815000 197.500000 ;
        RECT  8.615000 197.705000  8.815000 197.905000 ;
        RECT  8.720000  23.910000  8.920000  24.110000 ;
        RECT  8.720000  24.340000  8.920000  24.540000 ;
        RECT  8.720000  24.770000  8.920000  24.970000 ;
        RECT  8.720000  25.200000  8.920000  25.400000 ;
        RECT  8.720000  25.630000  8.920000  25.830000 ;
        RECT  8.720000  26.060000  8.920000  26.260000 ;
        RECT  8.720000  26.490000  8.920000  26.690000 ;
        RECT  8.720000  26.920000  8.920000  27.120000 ;
        RECT  8.720000  27.350000  8.920000  27.550000 ;
        RECT  8.720000  27.780000  8.920000  27.980000 ;
        RECT  8.720000  28.210000  8.920000  28.410000 ;
        RECT  9.015000 173.900000  9.215000 174.100000 ;
        RECT  9.015000 174.300000  9.215000 174.500000 ;
        RECT  9.015000 174.700000  9.215000 174.900000 ;
        RECT  9.015000 175.100000  9.215000 175.300000 ;
        RECT  9.015000 175.500000  9.215000 175.700000 ;
        RECT  9.015000 175.900000  9.215000 176.100000 ;
        RECT  9.015000 176.300000  9.215000 176.500000 ;
        RECT  9.015000 176.700000  9.215000 176.900000 ;
        RECT  9.015000 177.100000  9.215000 177.300000 ;
        RECT  9.015000 177.500000  9.215000 177.700000 ;
        RECT  9.015000 177.900000  9.215000 178.100000 ;
        RECT  9.015000 178.300000  9.215000 178.500000 ;
        RECT  9.015000 178.700000  9.215000 178.900000 ;
        RECT  9.015000 179.100000  9.215000 179.300000 ;
        RECT  9.015000 179.500000  9.215000 179.700000 ;
        RECT  9.015000 179.900000  9.215000 180.100000 ;
        RECT  9.015000 180.300000  9.215000 180.500000 ;
        RECT  9.015000 180.700000  9.215000 180.900000 ;
        RECT  9.015000 181.100000  9.215000 181.300000 ;
        RECT  9.015000 181.505000  9.215000 181.705000 ;
        RECT  9.015000 181.910000  9.215000 182.110000 ;
        RECT  9.015000 182.315000  9.215000 182.515000 ;
        RECT  9.015000 182.720000  9.215000 182.920000 ;
        RECT  9.015000 183.125000  9.215000 183.325000 ;
        RECT  9.015000 183.530000  9.215000 183.730000 ;
        RECT  9.015000 183.935000  9.215000 184.135000 ;
        RECT  9.015000 184.340000  9.215000 184.540000 ;
        RECT  9.015000 184.745000  9.215000 184.945000 ;
        RECT  9.015000 185.150000  9.215000 185.350000 ;
        RECT  9.015000 185.555000  9.215000 185.755000 ;
        RECT  9.015000 185.960000  9.215000 186.160000 ;
        RECT  9.015000 186.365000  9.215000 186.565000 ;
        RECT  9.015000 186.770000  9.215000 186.970000 ;
        RECT  9.015000 187.175000  9.215000 187.375000 ;
        RECT  9.015000 187.580000  9.215000 187.780000 ;
        RECT  9.015000 187.985000  9.215000 188.185000 ;
        RECT  9.015000 188.390000  9.215000 188.590000 ;
        RECT  9.015000 188.795000  9.215000 188.995000 ;
        RECT  9.015000 189.200000  9.215000 189.400000 ;
        RECT  9.015000 189.605000  9.215000 189.805000 ;
        RECT  9.015000 190.010000  9.215000 190.210000 ;
        RECT  9.015000 190.415000  9.215000 190.615000 ;
        RECT  9.015000 190.820000  9.215000 191.020000 ;
        RECT  9.015000 191.225000  9.215000 191.425000 ;
        RECT  9.015000 191.630000  9.215000 191.830000 ;
        RECT  9.015000 192.035000  9.215000 192.235000 ;
        RECT  9.015000 192.440000  9.215000 192.640000 ;
        RECT  9.015000 192.845000  9.215000 193.045000 ;
        RECT  9.015000 193.250000  9.215000 193.450000 ;
        RECT  9.015000 193.655000  9.215000 193.855000 ;
        RECT  9.015000 194.060000  9.215000 194.260000 ;
        RECT  9.015000 194.465000  9.215000 194.665000 ;
        RECT  9.015000 194.870000  9.215000 195.070000 ;
        RECT  9.015000 195.275000  9.215000 195.475000 ;
        RECT  9.015000 195.680000  9.215000 195.880000 ;
        RECT  9.015000 196.085000  9.215000 196.285000 ;
        RECT  9.015000 196.490000  9.215000 196.690000 ;
        RECT  9.015000 196.895000  9.215000 197.095000 ;
        RECT  9.015000 197.300000  9.215000 197.500000 ;
        RECT  9.015000 197.705000  9.215000 197.905000 ;
        RECT  9.125000  23.910000  9.325000  24.110000 ;
        RECT  9.125000  24.340000  9.325000  24.540000 ;
        RECT  9.125000  24.770000  9.325000  24.970000 ;
        RECT  9.125000  25.200000  9.325000  25.400000 ;
        RECT  9.125000  25.630000  9.325000  25.830000 ;
        RECT  9.125000  26.060000  9.325000  26.260000 ;
        RECT  9.125000  26.490000  9.325000  26.690000 ;
        RECT  9.125000  26.920000  9.325000  27.120000 ;
        RECT  9.125000  27.350000  9.325000  27.550000 ;
        RECT  9.125000  27.780000  9.325000  27.980000 ;
        RECT  9.125000  28.210000  9.325000  28.410000 ;
        RECT  9.415000 173.900000  9.615000 174.100000 ;
        RECT  9.415000 174.300000  9.615000 174.500000 ;
        RECT  9.415000 174.700000  9.615000 174.900000 ;
        RECT  9.415000 175.100000  9.615000 175.300000 ;
        RECT  9.415000 175.500000  9.615000 175.700000 ;
        RECT  9.415000 175.900000  9.615000 176.100000 ;
        RECT  9.415000 176.300000  9.615000 176.500000 ;
        RECT  9.415000 176.700000  9.615000 176.900000 ;
        RECT  9.415000 177.100000  9.615000 177.300000 ;
        RECT  9.415000 177.500000  9.615000 177.700000 ;
        RECT  9.415000 177.900000  9.615000 178.100000 ;
        RECT  9.415000 178.300000  9.615000 178.500000 ;
        RECT  9.415000 178.700000  9.615000 178.900000 ;
        RECT  9.415000 179.100000  9.615000 179.300000 ;
        RECT  9.415000 179.500000  9.615000 179.700000 ;
        RECT  9.415000 179.900000  9.615000 180.100000 ;
        RECT  9.415000 180.300000  9.615000 180.500000 ;
        RECT  9.415000 180.700000  9.615000 180.900000 ;
        RECT  9.415000 181.100000  9.615000 181.300000 ;
        RECT  9.415000 181.505000  9.615000 181.705000 ;
        RECT  9.415000 181.910000  9.615000 182.110000 ;
        RECT  9.415000 182.315000  9.615000 182.515000 ;
        RECT  9.415000 182.720000  9.615000 182.920000 ;
        RECT  9.415000 183.125000  9.615000 183.325000 ;
        RECT  9.415000 183.530000  9.615000 183.730000 ;
        RECT  9.415000 183.935000  9.615000 184.135000 ;
        RECT  9.415000 184.340000  9.615000 184.540000 ;
        RECT  9.415000 184.745000  9.615000 184.945000 ;
        RECT  9.415000 185.150000  9.615000 185.350000 ;
        RECT  9.415000 185.555000  9.615000 185.755000 ;
        RECT  9.415000 185.960000  9.615000 186.160000 ;
        RECT  9.415000 186.365000  9.615000 186.565000 ;
        RECT  9.415000 186.770000  9.615000 186.970000 ;
        RECT  9.415000 187.175000  9.615000 187.375000 ;
        RECT  9.415000 187.580000  9.615000 187.780000 ;
        RECT  9.415000 187.985000  9.615000 188.185000 ;
        RECT  9.415000 188.390000  9.615000 188.590000 ;
        RECT  9.415000 188.795000  9.615000 188.995000 ;
        RECT  9.415000 189.200000  9.615000 189.400000 ;
        RECT  9.415000 189.605000  9.615000 189.805000 ;
        RECT  9.415000 190.010000  9.615000 190.210000 ;
        RECT  9.415000 190.415000  9.615000 190.615000 ;
        RECT  9.415000 190.820000  9.615000 191.020000 ;
        RECT  9.415000 191.225000  9.615000 191.425000 ;
        RECT  9.415000 191.630000  9.615000 191.830000 ;
        RECT  9.415000 192.035000  9.615000 192.235000 ;
        RECT  9.415000 192.440000  9.615000 192.640000 ;
        RECT  9.415000 192.845000  9.615000 193.045000 ;
        RECT  9.415000 193.250000  9.615000 193.450000 ;
        RECT  9.415000 193.655000  9.615000 193.855000 ;
        RECT  9.415000 194.060000  9.615000 194.260000 ;
        RECT  9.415000 194.465000  9.615000 194.665000 ;
        RECT  9.415000 194.870000  9.615000 195.070000 ;
        RECT  9.415000 195.275000  9.615000 195.475000 ;
        RECT  9.415000 195.680000  9.615000 195.880000 ;
        RECT  9.415000 196.085000  9.615000 196.285000 ;
        RECT  9.415000 196.490000  9.615000 196.690000 ;
        RECT  9.415000 196.895000  9.615000 197.095000 ;
        RECT  9.415000 197.300000  9.615000 197.500000 ;
        RECT  9.415000 197.705000  9.615000 197.905000 ;
        RECT  9.530000  23.910000  9.730000  24.110000 ;
        RECT  9.530000  24.340000  9.730000  24.540000 ;
        RECT  9.530000  24.770000  9.730000  24.970000 ;
        RECT  9.530000  25.200000  9.730000  25.400000 ;
        RECT  9.530000  25.630000  9.730000  25.830000 ;
        RECT  9.530000  26.060000  9.730000  26.260000 ;
        RECT  9.530000  26.490000  9.730000  26.690000 ;
        RECT  9.530000  26.920000  9.730000  27.120000 ;
        RECT  9.530000  27.350000  9.730000  27.550000 ;
        RECT  9.530000  27.780000  9.730000  27.980000 ;
        RECT  9.530000  28.210000  9.730000  28.410000 ;
        RECT  9.815000 173.900000 10.015000 174.100000 ;
        RECT  9.815000 174.300000 10.015000 174.500000 ;
        RECT  9.815000 174.700000 10.015000 174.900000 ;
        RECT  9.815000 175.100000 10.015000 175.300000 ;
        RECT  9.815000 175.500000 10.015000 175.700000 ;
        RECT  9.815000 175.900000 10.015000 176.100000 ;
        RECT  9.815000 176.300000 10.015000 176.500000 ;
        RECT  9.815000 176.700000 10.015000 176.900000 ;
        RECT  9.815000 177.100000 10.015000 177.300000 ;
        RECT  9.815000 177.500000 10.015000 177.700000 ;
        RECT  9.815000 177.900000 10.015000 178.100000 ;
        RECT  9.815000 178.300000 10.015000 178.500000 ;
        RECT  9.815000 178.700000 10.015000 178.900000 ;
        RECT  9.815000 179.100000 10.015000 179.300000 ;
        RECT  9.815000 179.500000 10.015000 179.700000 ;
        RECT  9.815000 179.900000 10.015000 180.100000 ;
        RECT  9.815000 180.300000 10.015000 180.500000 ;
        RECT  9.815000 180.700000 10.015000 180.900000 ;
        RECT  9.815000 181.100000 10.015000 181.300000 ;
        RECT  9.815000 181.505000 10.015000 181.705000 ;
        RECT  9.815000 181.910000 10.015000 182.110000 ;
        RECT  9.815000 182.315000 10.015000 182.515000 ;
        RECT  9.815000 182.720000 10.015000 182.920000 ;
        RECT  9.815000 183.125000 10.015000 183.325000 ;
        RECT  9.815000 183.530000 10.015000 183.730000 ;
        RECT  9.815000 183.935000 10.015000 184.135000 ;
        RECT  9.815000 184.340000 10.015000 184.540000 ;
        RECT  9.815000 184.745000 10.015000 184.945000 ;
        RECT  9.815000 185.150000 10.015000 185.350000 ;
        RECT  9.815000 185.555000 10.015000 185.755000 ;
        RECT  9.815000 185.960000 10.015000 186.160000 ;
        RECT  9.815000 186.365000 10.015000 186.565000 ;
        RECT  9.815000 186.770000 10.015000 186.970000 ;
        RECT  9.815000 187.175000 10.015000 187.375000 ;
        RECT  9.815000 187.580000 10.015000 187.780000 ;
        RECT  9.815000 187.985000 10.015000 188.185000 ;
        RECT  9.815000 188.390000 10.015000 188.590000 ;
        RECT  9.815000 188.795000 10.015000 188.995000 ;
        RECT  9.815000 189.200000 10.015000 189.400000 ;
        RECT  9.815000 189.605000 10.015000 189.805000 ;
        RECT  9.815000 190.010000 10.015000 190.210000 ;
        RECT  9.815000 190.415000 10.015000 190.615000 ;
        RECT  9.815000 190.820000 10.015000 191.020000 ;
        RECT  9.815000 191.225000 10.015000 191.425000 ;
        RECT  9.815000 191.630000 10.015000 191.830000 ;
        RECT  9.815000 192.035000 10.015000 192.235000 ;
        RECT  9.815000 192.440000 10.015000 192.640000 ;
        RECT  9.815000 192.845000 10.015000 193.045000 ;
        RECT  9.815000 193.250000 10.015000 193.450000 ;
        RECT  9.815000 193.655000 10.015000 193.855000 ;
        RECT  9.815000 194.060000 10.015000 194.260000 ;
        RECT  9.815000 194.465000 10.015000 194.665000 ;
        RECT  9.815000 194.870000 10.015000 195.070000 ;
        RECT  9.815000 195.275000 10.015000 195.475000 ;
        RECT  9.815000 195.680000 10.015000 195.880000 ;
        RECT  9.815000 196.085000 10.015000 196.285000 ;
        RECT  9.815000 196.490000 10.015000 196.690000 ;
        RECT  9.815000 196.895000 10.015000 197.095000 ;
        RECT  9.815000 197.300000 10.015000 197.500000 ;
        RECT  9.815000 197.705000 10.015000 197.905000 ;
        RECT  9.935000  23.910000 10.135000  24.110000 ;
        RECT  9.935000  24.340000 10.135000  24.540000 ;
        RECT  9.935000  24.770000 10.135000  24.970000 ;
        RECT  9.935000  25.200000 10.135000  25.400000 ;
        RECT  9.935000  25.630000 10.135000  25.830000 ;
        RECT  9.935000  26.060000 10.135000  26.260000 ;
        RECT  9.935000  26.490000 10.135000  26.690000 ;
        RECT  9.935000  26.920000 10.135000  27.120000 ;
        RECT  9.935000  27.350000 10.135000  27.550000 ;
        RECT  9.935000  27.780000 10.135000  27.980000 ;
        RECT  9.935000  28.210000 10.135000  28.410000 ;
        RECT 10.215000 173.900000 10.415000 174.100000 ;
        RECT 10.215000 174.300000 10.415000 174.500000 ;
        RECT 10.215000 174.700000 10.415000 174.900000 ;
        RECT 10.215000 175.100000 10.415000 175.300000 ;
        RECT 10.215000 175.500000 10.415000 175.700000 ;
        RECT 10.215000 175.900000 10.415000 176.100000 ;
        RECT 10.215000 176.300000 10.415000 176.500000 ;
        RECT 10.215000 176.700000 10.415000 176.900000 ;
        RECT 10.215000 177.100000 10.415000 177.300000 ;
        RECT 10.215000 177.500000 10.415000 177.700000 ;
        RECT 10.215000 177.900000 10.415000 178.100000 ;
        RECT 10.215000 178.300000 10.415000 178.500000 ;
        RECT 10.215000 178.700000 10.415000 178.900000 ;
        RECT 10.215000 179.100000 10.415000 179.300000 ;
        RECT 10.215000 179.500000 10.415000 179.700000 ;
        RECT 10.215000 179.900000 10.415000 180.100000 ;
        RECT 10.215000 180.300000 10.415000 180.500000 ;
        RECT 10.215000 180.700000 10.415000 180.900000 ;
        RECT 10.215000 181.100000 10.415000 181.300000 ;
        RECT 10.215000 181.505000 10.415000 181.705000 ;
        RECT 10.215000 181.910000 10.415000 182.110000 ;
        RECT 10.215000 182.315000 10.415000 182.515000 ;
        RECT 10.215000 182.720000 10.415000 182.920000 ;
        RECT 10.215000 183.125000 10.415000 183.325000 ;
        RECT 10.215000 183.530000 10.415000 183.730000 ;
        RECT 10.215000 183.935000 10.415000 184.135000 ;
        RECT 10.215000 184.340000 10.415000 184.540000 ;
        RECT 10.215000 184.745000 10.415000 184.945000 ;
        RECT 10.215000 185.150000 10.415000 185.350000 ;
        RECT 10.215000 185.555000 10.415000 185.755000 ;
        RECT 10.215000 185.960000 10.415000 186.160000 ;
        RECT 10.215000 186.365000 10.415000 186.565000 ;
        RECT 10.215000 186.770000 10.415000 186.970000 ;
        RECT 10.215000 187.175000 10.415000 187.375000 ;
        RECT 10.215000 187.580000 10.415000 187.780000 ;
        RECT 10.215000 187.985000 10.415000 188.185000 ;
        RECT 10.215000 188.390000 10.415000 188.590000 ;
        RECT 10.215000 188.795000 10.415000 188.995000 ;
        RECT 10.215000 189.200000 10.415000 189.400000 ;
        RECT 10.215000 189.605000 10.415000 189.805000 ;
        RECT 10.215000 190.010000 10.415000 190.210000 ;
        RECT 10.215000 190.415000 10.415000 190.615000 ;
        RECT 10.215000 190.820000 10.415000 191.020000 ;
        RECT 10.215000 191.225000 10.415000 191.425000 ;
        RECT 10.215000 191.630000 10.415000 191.830000 ;
        RECT 10.215000 192.035000 10.415000 192.235000 ;
        RECT 10.215000 192.440000 10.415000 192.640000 ;
        RECT 10.215000 192.845000 10.415000 193.045000 ;
        RECT 10.215000 193.250000 10.415000 193.450000 ;
        RECT 10.215000 193.655000 10.415000 193.855000 ;
        RECT 10.215000 194.060000 10.415000 194.260000 ;
        RECT 10.215000 194.465000 10.415000 194.665000 ;
        RECT 10.215000 194.870000 10.415000 195.070000 ;
        RECT 10.215000 195.275000 10.415000 195.475000 ;
        RECT 10.215000 195.680000 10.415000 195.880000 ;
        RECT 10.215000 196.085000 10.415000 196.285000 ;
        RECT 10.215000 196.490000 10.415000 196.690000 ;
        RECT 10.215000 196.895000 10.415000 197.095000 ;
        RECT 10.215000 197.300000 10.415000 197.500000 ;
        RECT 10.215000 197.705000 10.415000 197.905000 ;
        RECT 10.340000  23.910000 10.540000  24.110000 ;
        RECT 10.340000  24.340000 10.540000  24.540000 ;
        RECT 10.340000  24.770000 10.540000  24.970000 ;
        RECT 10.340000  25.200000 10.540000  25.400000 ;
        RECT 10.340000  25.630000 10.540000  25.830000 ;
        RECT 10.340000  26.060000 10.540000  26.260000 ;
        RECT 10.340000  26.490000 10.540000  26.690000 ;
        RECT 10.340000  26.920000 10.540000  27.120000 ;
        RECT 10.340000  27.350000 10.540000  27.550000 ;
        RECT 10.340000  27.780000 10.540000  27.980000 ;
        RECT 10.340000  28.210000 10.540000  28.410000 ;
        RECT 10.615000 173.900000 10.815000 174.100000 ;
        RECT 10.615000 174.300000 10.815000 174.500000 ;
        RECT 10.615000 174.700000 10.815000 174.900000 ;
        RECT 10.615000 175.100000 10.815000 175.300000 ;
        RECT 10.615000 175.500000 10.815000 175.700000 ;
        RECT 10.615000 175.900000 10.815000 176.100000 ;
        RECT 10.615000 176.300000 10.815000 176.500000 ;
        RECT 10.615000 176.700000 10.815000 176.900000 ;
        RECT 10.615000 177.100000 10.815000 177.300000 ;
        RECT 10.615000 177.500000 10.815000 177.700000 ;
        RECT 10.615000 177.900000 10.815000 178.100000 ;
        RECT 10.615000 178.300000 10.815000 178.500000 ;
        RECT 10.615000 178.700000 10.815000 178.900000 ;
        RECT 10.615000 179.100000 10.815000 179.300000 ;
        RECT 10.615000 179.500000 10.815000 179.700000 ;
        RECT 10.615000 179.900000 10.815000 180.100000 ;
        RECT 10.615000 180.300000 10.815000 180.500000 ;
        RECT 10.615000 180.700000 10.815000 180.900000 ;
        RECT 10.615000 181.100000 10.815000 181.300000 ;
        RECT 10.615000 181.505000 10.815000 181.705000 ;
        RECT 10.615000 181.910000 10.815000 182.110000 ;
        RECT 10.615000 182.315000 10.815000 182.515000 ;
        RECT 10.615000 182.720000 10.815000 182.920000 ;
        RECT 10.615000 183.125000 10.815000 183.325000 ;
        RECT 10.615000 183.530000 10.815000 183.730000 ;
        RECT 10.615000 183.935000 10.815000 184.135000 ;
        RECT 10.615000 184.340000 10.815000 184.540000 ;
        RECT 10.615000 184.745000 10.815000 184.945000 ;
        RECT 10.615000 185.150000 10.815000 185.350000 ;
        RECT 10.615000 185.555000 10.815000 185.755000 ;
        RECT 10.615000 185.960000 10.815000 186.160000 ;
        RECT 10.615000 186.365000 10.815000 186.565000 ;
        RECT 10.615000 186.770000 10.815000 186.970000 ;
        RECT 10.615000 187.175000 10.815000 187.375000 ;
        RECT 10.615000 187.580000 10.815000 187.780000 ;
        RECT 10.615000 187.985000 10.815000 188.185000 ;
        RECT 10.615000 188.390000 10.815000 188.590000 ;
        RECT 10.615000 188.795000 10.815000 188.995000 ;
        RECT 10.615000 189.200000 10.815000 189.400000 ;
        RECT 10.615000 189.605000 10.815000 189.805000 ;
        RECT 10.615000 190.010000 10.815000 190.210000 ;
        RECT 10.615000 190.415000 10.815000 190.615000 ;
        RECT 10.615000 190.820000 10.815000 191.020000 ;
        RECT 10.615000 191.225000 10.815000 191.425000 ;
        RECT 10.615000 191.630000 10.815000 191.830000 ;
        RECT 10.615000 192.035000 10.815000 192.235000 ;
        RECT 10.615000 192.440000 10.815000 192.640000 ;
        RECT 10.615000 192.845000 10.815000 193.045000 ;
        RECT 10.615000 193.250000 10.815000 193.450000 ;
        RECT 10.615000 193.655000 10.815000 193.855000 ;
        RECT 10.615000 194.060000 10.815000 194.260000 ;
        RECT 10.615000 194.465000 10.815000 194.665000 ;
        RECT 10.615000 194.870000 10.815000 195.070000 ;
        RECT 10.615000 195.275000 10.815000 195.475000 ;
        RECT 10.615000 195.680000 10.815000 195.880000 ;
        RECT 10.615000 196.085000 10.815000 196.285000 ;
        RECT 10.615000 196.490000 10.815000 196.690000 ;
        RECT 10.615000 196.895000 10.815000 197.095000 ;
        RECT 10.615000 197.300000 10.815000 197.500000 ;
        RECT 10.615000 197.705000 10.815000 197.905000 ;
        RECT 10.745000  23.910000 10.945000  24.110000 ;
        RECT 10.745000  24.340000 10.945000  24.540000 ;
        RECT 10.745000  24.770000 10.945000  24.970000 ;
        RECT 10.745000  25.200000 10.945000  25.400000 ;
        RECT 10.745000  25.630000 10.945000  25.830000 ;
        RECT 10.745000  26.060000 10.945000  26.260000 ;
        RECT 10.745000  26.490000 10.945000  26.690000 ;
        RECT 10.745000  26.920000 10.945000  27.120000 ;
        RECT 10.745000  27.350000 10.945000  27.550000 ;
        RECT 10.745000  27.780000 10.945000  27.980000 ;
        RECT 10.745000  28.210000 10.945000  28.410000 ;
        RECT 11.015000 173.900000 11.215000 174.100000 ;
        RECT 11.015000 174.300000 11.215000 174.500000 ;
        RECT 11.015000 174.700000 11.215000 174.900000 ;
        RECT 11.015000 175.100000 11.215000 175.300000 ;
        RECT 11.015000 175.500000 11.215000 175.700000 ;
        RECT 11.015000 175.900000 11.215000 176.100000 ;
        RECT 11.015000 176.300000 11.215000 176.500000 ;
        RECT 11.015000 176.700000 11.215000 176.900000 ;
        RECT 11.015000 177.100000 11.215000 177.300000 ;
        RECT 11.015000 177.500000 11.215000 177.700000 ;
        RECT 11.015000 177.900000 11.215000 178.100000 ;
        RECT 11.015000 178.300000 11.215000 178.500000 ;
        RECT 11.015000 178.700000 11.215000 178.900000 ;
        RECT 11.015000 179.100000 11.215000 179.300000 ;
        RECT 11.015000 179.500000 11.215000 179.700000 ;
        RECT 11.015000 179.900000 11.215000 180.100000 ;
        RECT 11.015000 180.300000 11.215000 180.500000 ;
        RECT 11.015000 180.700000 11.215000 180.900000 ;
        RECT 11.015000 181.100000 11.215000 181.300000 ;
        RECT 11.015000 181.505000 11.215000 181.705000 ;
        RECT 11.015000 181.910000 11.215000 182.110000 ;
        RECT 11.015000 182.315000 11.215000 182.515000 ;
        RECT 11.015000 182.720000 11.215000 182.920000 ;
        RECT 11.015000 183.125000 11.215000 183.325000 ;
        RECT 11.015000 183.530000 11.215000 183.730000 ;
        RECT 11.015000 183.935000 11.215000 184.135000 ;
        RECT 11.015000 184.340000 11.215000 184.540000 ;
        RECT 11.015000 184.745000 11.215000 184.945000 ;
        RECT 11.015000 185.150000 11.215000 185.350000 ;
        RECT 11.015000 185.555000 11.215000 185.755000 ;
        RECT 11.015000 185.960000 11.215000 186.160000 ;
        RECT 11.015000 186.365000 11.215000 186.565000 ;
        RECT 11.015000 186.770000 11.215000 186.970000 ;
        RECT 11.015000 187.175000 11.215000 187.375000 ;
        RECT 11.015000 187.580000 11.215000 187.780000 ;
        RECT 11.015000 187.985000 11.215000 188.185000 ;
        RECT 11.015000 188.390000 11.215000 188.590000 ;
        RECT 11.015000 188.795000 11.215000 188.995000 ;
        RECT 11.015000 189.200000 11.215000 189.400000 ;
        RECT 11.015000 189.605000 11.215000 189.805000 ;
        RECT 11.015000 190.010000 11.215000 190.210000 ;
        RECT 11.015000 190.415000 11.215000 190.615000 ;
        RECT 11.015000 190.820000 11.215000 191.020000 ;
        RECT 11.015000 191.225000 11.215000 191.425000 ;
        RECT 11.015000 191.630000 11.215000 191.830000 ;
        RECT 11.015000 192.035000 11.215000 192.235000 ;
        RECT 11.015000 192.440000 11.215000 192.640000 ;
        RECT 11.015000 192.845000 11.215000 193.045000 ;
        RECT 11.015000 193.250000 11.215000 193.450000 ;
        RECT 11.015000 193.655000 11.215000 193.855000 ;
        RECT 11.015000 194.060000 11.215000 194.260000 ;
        RECT 11.015000 194.465000 11.215000 194.665000 ;
        RECT 11.015000 194.870000 11.215000 195.070000 ;
        RECT 11.015000 195.275000 11.215000 195.475000 ;
        RECT 11.015000 195.680000 11.215000 195.880000 ;
        RECT 11.015000 196.085000 11.215000 196.285000 ;
        RECT 11.015000 196.490000 11.215000 196.690000 ;
        RECT 11.015000 196.895000 11.215000 197.095000 ;
        RECT 11.015000 197.300000 11.215000 197.500000 ;
        RECT 11.015000 197.705000 11.215000 197.905000 ;
        RECT 11.150000  23.910000 11.350000  24.110000 ;
        RECT 11.150000  24.340000 11.350000  24.540000 ;
        RECT 11.150000  24.770000 11.350000  24.970000 ;
        RECT 11.150000  25.200000 11.350000  25.400000 ;
        RECT 11.150000  25.630000 11.350000  25.830000 ;
        RECT 11.150000  26.060000 11.350000  26.260000 ;
        RECT 11.150000  26.490000 11.350000  26.690000 ;
        RECT 11.150000  26.920000 11.350000  27.120000 ;
        RECT 11.150000  27.350000 11.350000  27.550000 ;
        RECT 11.150000  27.780000 11.350000  27.980000 ;
        RECT 11.150000  28.210000 11.350000  28.410000 ;
        RECT 11.415000 173.900000 11.615000 174.100000 ;
        RECT 11.415000 174.300000 11.615000 174.500000 ;
        RECT 11.415000 174.700000 11.615000 174.900000 ;
        RECT 11.415000 175.100000 11.615000 175.300000 ;
        RECT 11.415000 175.500000 11.615000 175.700000 ;
        RECT 11.415000 175.900000 11.615000 176.100000 ;
        RECT 11.415000 176.300000 11.615000 176.500000 ;
        RECT 11.415000 176.700000 11.615000 176.900000 ;
        RECT 11.415000 177.100000 11.615000 177.300000 ;
        RECT 11.415000 177.500000 11.615000 177.700000 ;
        RECT 11.415000 177.900000 11.615000 178.100000 ;
        RECT 11.415000 178.300000 11.615000 178.500000 ;
        RECT 11.415000 178.700000 11.615000 178.900000 ;
        RECT 11.415000 179.100000 11.615000 179.300000 ;
        RECT 11.415000 179.500000 11.615000 179.700000 ;
        RECT 11.415000 179.900000 11.615000 180.100000 ;
        RECT 11.415000 180.300000 11.615000 180.500000 ;
        RECT 11.415000 180.700000 11.615000 180.900000 ;
        RECT 11.415000 181.100000 11.615000 181.300000 ;
        RECT 11.415000 181.505000 11.615000 181.705000 ;
        RECT 11.415000 181.910000 11.615000 182.110000 ;
        RECT 11.415000 182.315000 11.615000 182.515000 ;
        RECT 11.415000 182.720000 11.615000 182.920000 ;
        RECT 11.415000 183.125000 11.615000 183.325000 ;
        RECT 11.415000 183.530000 11.615000 183.730000 ;
        RECT 11.415000 183.935000 11.615000 184.135000 ;
        RECT 11.415000 184.340000 11.615000 184.540000 ;
        RECT 11.415000 184.745000 11.615000 184.945000 ;
        RECT 11.415000 185.150000 11.615000 185.350000 ;
        RECT 11.415000 185.555000 11.615000 185.755000 ;
        RECT 11.415000 185.960000 11.615000 186.160000 ;
        RECT 11.415000 186.365000 11.615000 186.565000 ;
        RECT 11.415000 186.770000 11.615000 186.970000 ;
        RECT 11.415000 187.175000 11.615000 187.375000 ;
        RECT 11.415000 187.580000 11.615000 187.780000 ;
        RECT 11.415000 187.985000 11.615000 188.185000 ;
        RECT 11.415000 188.390000 11.615000 188.590000 ;
        RECT 11.415000 188.795000 11.615000 188.995000 ;
        RECT 11.415000 189.200000 11.615000 189.400000 ;
        RECT 11.415000 189.605000 11.615000 189.805000 ;
        RECT 11.415000 190.010000 11.615000 190.210000 ;
        RECT 11.415000 190.415000 11.615000 190.615000 ;
        RECT 11.415000 190.820000 11.615000 191.020000 ;
        RECT 11.415000 191.225000 11.615000 191.425000 ;
        RECT 11.415000 191.630000 11.615000 191.830000 ;
        RECT 11.415000 192.035000 11.615000 192.235000 ;
        RECT 11.415000 192.440000 11.615000 192.640000 ;
        RECT 11.415000 192.845000 11.615000 193.045000 ;
        RECT 11.415000 193.250000 11.615000 193.450000 ;
        RECT 11.415000 193.655000 11.615000 193.855000 ;
        RECT 11.415000 194.060000 11.615000 194.260000 ;
        RECT 11.415000 194.465000 11.615000 194.665000 ;
        RECT 11.415000 194.870000 11.615000 195.070000 ;
        RECT 11.415000 195.275000 11.615000 195.475000 ;
        RECT 11.415000 195.680000 11.615000 195.880000 ;
        RECT 11.415000 196.085000 11.615000 196.285000 ;
        RECT 11.415000 196.490000 11.615000 196.690000 ;
        RECT 11.415000 196.895000 11.615000 197.095000 ;
        RECT 11.415000 197.300000 11.615000 197.500000 ;
        RECT 11.415000 197.705000 11.615000 197.905000 ;
        RECT 11.555000  23.910000 11.755000  24.110000 ;
        RECT 11.555000  24.340000 11.755000  24.540000 ;
        RECT 11.555000  24.770000 11.755000  24.970000 ;
        RECT 11.555000  25.200000 11.755000  25.400000 ;
        RECT 11.555000  25.630000 11.755000  25.830000 ;
        RECT 11.555000  26.060000 11.755000  26.260000 ;
        RECT 11.555000  26.490000 11.755000  26.690000 ;
        RECT 11.555000  26.920000 11.755000  27.120000 ;
        RECT 11.555000  27.350000 11.755000  27.550000 ;
        RECT 11.555000  27.780000 11.755000  27.980000 ;
        RECT 11.555000  28.210000 11.755000  28.410000 ;
        RECT 11.815000 173.900000 12.015000 174.100000 ;
        RECT 11.815000 174.300000 12.015000 174.500000 ;
        RECT 11.815000 174.700000 12.015000 174.900000 ;
        RECT 11.815000 175.100000 12.015000 175.300000 ;
        RECT 11.815000 175.500000 12.015000 175.700000 ;
        RECT 11.815000 175.900000 12.015000 176.100000 ;
        RECT 11.815000 176.300000 12.015000 176.500000 ;
        RECT 11.815000 176.700000 12.015000 176.900000 ;
        RECT 11.815000 177.100000 12.015000 177.300000 ;
        RECT 11.815000 177.500000 12.015000 177.700000 ;
        RECT 11.815000 177.900000 12.015000 178.100000 ;
        RECT 11.815000 178.300000 12.015000 178.500000 ;
        RECT 11.815000 178.700000 12.015000 178.900000 ;
        RECT 11.815000 179.100000 12.015000 179.300000 ;
        RECT 11.815000 179.500000 12.015000 179.700000 ;
        RECT 11.815000 179.900000 12.015000 180.100000 ;
        RECT 11.815000 180.300000 12.015000 180.500000 ;
        RECT 11.815000 180.700000 12.015000 180.900000 ;
        RECT 11.815000 181.100000 12.015000 181.300000 ;
        RECT 11.815000 181.505000 12.015000 181.705000 ;
        RECT 11.815000 181.910000 12.015000 182.110000 ;
        RECT 11.815000 182.315000 12.015000 182.515000 ;
        RECT 11.815000 182.720000 12.015000 182.920000 ;
        RECT 11.815000 183.125000 12.015000 183.325000 ;
        RECT 11.815000 183.530000 12.015000 183.730000 ;
        RECT 11.815000 183.935000 12.015000 184.135000 ;
        RECT 11.815000 184.340000 12.015000 184.540000 ;
        RECT 11.815000 184.745000 12.015000 184.945000 ;
        RECT 11.815000 185.150000 12.015000 185.350000 ;
        RECT 11.815000 185.555000 12.015000 185.755000 ;
        RECT 11.815000 185.960000 12.015000 186.160000 ;
        RECT 11.815000 186.365000 12.015000 186.565000 ;
        RECT 11.815000 186.770000 12.015000 186.970000 ;
        RECT 11.815000 187.175000 12.015000 187.375000 ;
        RECT 11.815000 187.580000 12.015000 187.780000 ;
        RECT 11.815000 187.985000 12.015000 188.185000 ;
        RECT 11.815000 188.390000 12.015000 188.590000 ;
        RECT 11.815000 188.795000 12.015000 188.995000 ;
        RECT 11.815000 189.200000 12.015000 189.400000 ;
        RECT 11.815000 189.605000 12.015000 189.805000 ;
        RECT 11.815000 190.010000 12.015000 190.210000 ;
        RECT 11.815000 190.415000 12.015000 190.615000 ;
        RECT 11.815000 190.820000 12.015000 191.020000 ;
        RECT 11.815000 191.225000 12.015000 191.425000 ;
        RECT 11.815000 191.630000 12.015000 191.830000 ;
        RECT 11.815000 192.035000 12.015000 192.235000 ;
        RECT 11.815000 192.440000 12.015000 192.640000 ;
        RECT 11.815000 192.845000 12.015000 193.045000 ;
        RECT 11.815000 193.250000 12.015000 193.450000 ;
        RECT 11.815000 193.655000 12.015000 193.855000 ;
        RECT 11.815000 194.060000 12.015000 194.260000 ;
        RECT 11.815000 194.465000 12.015000 194.665000 ;
        RECT 11.815000 194.870000 12.015000 195.070000 ;
        RECT 11.815000 195.275000 12.015000 195.475000 ;
        RECT 11.815000 195.680000 12.015000 195.880000 ;
        RECT 11.815000 196.085000 12.015000 196.285000 ;
        RECT 11.815000 196.490000 12.015000 196.690000 ;
        RECT 11.815000 196.895000 12.015000 197.095000 ;
        RECT 11.815000 197.300000 12.015000 197.500000 ;
        RECT 11.815000 197.705000 12.015000 197.905000 ;
        RECT 11.960000  23.910000 12.160000  24.110000 ;
        RECT 11.960000  24.340000 12.160000  24.540000 ;
        RECT 11.960000  24.770000 12.160000  24.970000 ;
        RECT 11.960000  25.200000 12.160000  25.400000 ;
        RECT 11.960000  25.630000 12.160000  25.830000 ;
        RECT 11.960000  26.060000 12.160000  26.260000 ;
        RECT 11.960000  26.490000 12.160000  26.690000 ;
        RECT 11.960000  26.920000 12.160000  27.120000 ;
        RECT 11.960000  27.350000 12.160000  27.550000 ;
        RECT 11.960000  27.780000 12.160000  27.980000 ;
        RECT 11.960000  28.210000 12.160000  28.410000 ;
        RECT 12.215000 173.900000 12.415000 174.100000 ;
        RECT 12.215000 174.300000 12.415000 174.500000 ;
        RECT 12.215000 174.700000 12.415000 174.900000 ;
        RECT 12.215000 175.100000 12.415000 175.300000 ;
        RECT 12.215000 175.500000 12.415000 175.700000 ;
        RECT 12.215000 175.900000 12.415000 176.100000 ;
        RECT 12.215000 176.300000 12.415000 176.500000 ;
        RECT 12.215000 176.700000 12.415000 176.900000 ;
        RECT 12.215000 177.100000 12.415000 177.300000 ;
        RECT 12.215000 177.500000 12.415000 177.700000 ;
        RECT 12.215000 177.900000 12.415000 178.100000 ;
        RECT 12.215000 178.300000 12.415000 178.500000 ;
        RECT 12.215000 178.700000 12.415000 178.900000 ;
        RECT 12.215000 179.100000 12.415000 179.300000 ;
        RECT 12.215000 179.500000 12.415000 179.700000 ;
        RECT 12.215000 179.900000 12.415000 180.100000 ;
        RECT 12.215000 180.300000 12.415000 180.500000 ;
        RECT 12.215000 180.700000 12.415000 180.900000 ;
        RECT 12.215000 181.100000 12.415000 181.300000 ;
        RECT 12.215000 181.505000 12.415000 181.705000 ;
        RECT 12.215000 181.910000 12.415000 182.110000 ;
        RECT 12.215000 182.315000 12.415000 182.515000 ;
        RECT 12.215000 182.720000 12.415000 182.920000 ;
        RECT 12.215000 183.125000 12.415000 183.325000 ;
        RECT 12.215000 183.530000 12.415000 183.730000 ;
        RECT 12.215000 183.935000 12.415000 184.135000 ;
        RECT 12.215000 184.340000 12.415000 184.540000 ;
        RECT 12.215000 184.745000 12.415000 184.945000 ;
        RECT 12.215000 185.150000 12.415000 185.350000 ;
        RECT 12.215000 185.555000 12.415000 185.755000 ;
        RECT 12.215000 185.960000 12.415000 186.160000 ;
        RECT 12.215000 186.365000 12.415000 186.565000 ;
        RECT 12.215000 186.770000 12.415000 186.970000 ;
        RECT 12.215000 187.175000 12.415000 187.375000 ;
        RECT 12.215000 187.580000 12.415000 187.780000 ;
        RECT 12.215000 187.985000 12.415000 188.185000 ;
        RECT 12.215000 188.390000 12.415000 188.590000 ;
        RECT 12.215000 188.795000 12.415000 188.995000 ;
        RECT 12.215000 189.200000 12.415000 189.400000 ;
        RECT 12.215000 189.605000 12.415000 189.805000 ;
        RECT 12.215000 190.010000 12.415000 190.210000 ;
        RECT 12.215000 190.415000 12.415000 190.615000 ;
        RECT 12.215000 190.820000 12.415000 191.020000 ;
        RECT 12.215000 191.225000 12.415000 191.425000 ;
        RECT 12.215000 191.630000 12.415000 191.830000 ;
        RECT 12.215000 192.035000 12.415000 192.235000 ;
        RECT 12.215000 192.440000 12.415000 192.640000 ;
        RECT 12.215000 192.845000 12.415000 193.045000 ;
        RECT 12.215000 193.250000 12.415000 193.450000 ;
        RECT 12.215000 193.655000 12.415000 193.855000 ;
        RECT 12.215000 194.060000 12.415000 194.260000 ;
        RECT 12.215000 194.465000 12.415000 194.665000 ;
        RECT 12.215000 194.870000 12.415000 195.070000 ;
        RECT 12.215000 195.275000 12.415000 195.475000 ;
        RECT 12.215000 195.680000 12.415000 195.880000 ;
        RECT 12.215000 196.085000 12.415000 196.285000 ;
        RECT 12.215000 196.490000 12.415000 196.690000 ;
        RECT 12.215000 196.895000 12.415000 197.095000 ;
        RECT 12.215000 197.300000 12.415000 197.500000 ;
        RECT 12.215000 197.705000 12.415000 197.905000 ;
        RECT 12.365000  23.910000 12.565000  24.110000 ;
        RECT 12.365000  24.340000 12.565000  24.540000 ;
        RECT 12.365000  24.770000 12.565000  24.970000 ;
        RECT 12.365000  25.200000 12.565000  25.400000 ;
        RECT 12.365000  25.630000 12.565000  25.830000 ;
        RECT 12.365000  26.060000 12.565000  26.260000 ;
        RECT 12.365000  26.490000 12.565000  26.690000 ;
        RECT 12.365000  26.920000 12.565000  27.120000 ;
        RECT 12.365000  27.350000 12.565000  27.550000 ;
        RECT 12.365000  27.780000 12.565000  27.980000 ;
        RECT 12.365000  28.210000 12.565000  28.410000 ;
        RECT 12.615000 173.900000 12.815000 174.100000 ;
        RECT 12.615000 174.300000 12.815000 174.500000 ;
        RECT 12.615000 174.700000 12.815000 174.900000 ;
        RECT 12.615000 175.100000 12.815000 175.300000 ;
        RECT 12.615000 175.500000 12.815000 175.700000 ;
        RECT 12.615000 175.900000 12.815000 176.100000 ;
        RECT 12.615000 176.300000 12.815000 176.500000 ;
        RECT 12.615000 176.700000 12.815000 176.900000 ;
        RECT 12.615000 177.100000 12.815000 177.300000 ;
        RECT 12.615000 177.500000 12.815000 177.700000 ;
        RECT 12.615000 177.900000 12.815000 178.100000 ;
        RECT 12.615000 178.300000 12.815000 178.500000 ;
        RECT 12.615000 178.700000 12.815000 178.900000 ;
        RECT 12.615000 179.100000 12.815000 179.300000 ;
        RECT 12.615000 179.500000 12.815000 179.700000 ;
        RECT 12.615000 179.900000 12.815000 180.100000 ;
        RECT 12.615000 180.300000 12.815000 180.500000 ;
        RECT 12.615000 180.700000 12.815000 180.900000 ;
        RECT 12.615000 181.100000 12.815000 181.300000 ;
        RECT 12.615000 181.505000 12.815000 181.705000 ;
        RECT 12.615000 181.910000 12.815000 182.110000 ;
        RECT 12.615000 182.315000 12.815000 182.515000 ;
        RECT 12.615000 182.720000 12.815000 182.920000 ;
        RECT 12.615000 183.125000 12.815000 183.325000 ;
        RECT 12.615000 183.530000 12.815000 183.730000 ;
        RECT 12.615000 183.935000 12.815000 184.135000 ;
        RECT 12.615000 184.340000 12.815000 184.540000 ;
        RECT 12.615000 184.745000 12.815000 184.945000 ;
        RECT 12.615000 185.150000 12.815000 185.350000 ;
        RECT 12.615000 185.555000 12.815000 185.755000 ;
        RECT 12.615000 185.960000 12.815000 186.160000 ;
        RECT 12.615000 186.365000 12.815000 186.565000 ;
        RECT 12.615000 186.770000 12.815000 186.970000 ;
        RECT 12.615000 187.175000 12.815000 187.375000 ;
        RECT 12.615000 187.580000 12.815000 187.780000 ;
        RECT 12.615000 187.985000 12.815000 188.185000 ;
        RECT 12.615000 188.390000 12.815000 188.590000 ;
        RECT 12.615000 188.795000 12.815000 188.995000 ;
        RECT 12.615000 189.200000 12.815000 189.400000 ;
        RECT 12.615000 189.605000 12.815000 189.805000 ;
        RECT 12.615000 190.010000 12.815000 190.210000 ;
        RECT 12.615000 190.415000 12.815000 190.615000 ;
        RECT 12.615000 190.820000 12.815000 191.020000 ;
        RECT 12.615000 191.225000 12.815000 191.425000 ;
        RECT 12.615000 191.630000 12.815000 191.830000 ;
        RECT 12.615000 192.035000 12.815000 192.235000 ;
        RECT 12.615000 192.440000 12.815000 192.640000 ;
        RECT 12.615000 192.845000 12.815000 193.045000 ;
        RECT 12.615000 193.250000 12.815000 193.450000 ;
        RECT 12.615000 193.655000 12.815000 193.855000 ;
        RECT 12.615000 194.060000 12.815000 194.260000 ;
        RECT 12.615000 194.465000 12.815000 194.665000 ;
        RECT 12.615000 194.870000 12.815000 195.070000 ;
        RECT 12.615000 195.275000 12.815000 195.475000 ;
        RECT 12.615000 195.680000 12.815000 195.880000 ;
        RECT 12.615000 196.085000 12.815000 196.285000 ;
        RECT 12.615000 196.490000 12.815000 196.690000 ;
        RECT 12.615000 196.895000 12.815000 197.095000 ;
        RECT 12.615000 197.300000 12.815000 197.500000 ;
        RECT 12.615000 197.705000 12.815000 197.905000 ;
        RECT 12.770000  23.910000 12.970000  24.110000 ;
        RECT 12.770000  24.340000 12.970000  24.540000 ;
        RECT 12.770000  24.770000 12.970000  24.970000 ;
        RECT 12.770000  25.200000 12.970000  25.400000 ;
        RECT 12.770000  25.630000 12.970000  25.830000 ;
        RECT 12.770000  26.060000 12.970000  26.260000 ;
        RECT 12.770000  26.490000 12.970000  26.690000 ;
        RECT 12.770000  26.920000 12.970000  27.120000 ;
        RECT 12.770000  27.350000 12.970000  27.550000 ;
        RECT 12.770000  27.780000 12.970000  27.980000 ;
        RECT 12.770000  28.210000 12.970000  28.410000 ;
        RECT 13.175000  23.910000 13.375000  24.110000 ;
        RECT 13.175000  24.340000 13.375000  24.540000 ;
        RECT 13.175000  24.770000 13.375000  24.970000 ;
        RECT 13.175000  25.200000 13.375000  25.400000 ;
        RECT 13.175000  25.630000 13.375000  25.830000 ;
        RECT 13.175000  26.060000 13.375000  26.260000 ;
        RECT 13.175000  26.490000 13.375000  26.690000 ;
        RECT 13.175000  26.920000 13.375000  27.120000 ;
        RECT 13.175000  27.350000 13.375000  27.550000 ;
        RECT 13.175000  27.780000 13.375000  27.980000 ;
        RECT 13.175000  28.210000 13.375000  28.410000 ;
        RECT 13.580000  23.910000 13.780000  24.110000 ;
        RECT 13.580000  24.340000 13.780000  24.540000 ;
        RECT 13.580000  24.770000 13.780000  24.970000 ;
        RECT 13.580000  25.200000 13.780000  25.400000 ;
        RECT 13.580000  25.630000 13.780000  25.830000 ;
        RECT 13.580000  26.060000 13.780000  26.260000 ;
        RECT 13.580000  26.490000 13.780000  26.690000 ;
        RECT 13.580000  26.920000 13.780000  27.120000 ;
        RECT 13.580000  27.350000 13.780000  27.550000 ;
        RECT 13.580000  27.780000 13.780000  27.980000 ;
        RECT 13.580000  28.210000 13.780000  28.410000 ;
        RECT 13.985000  23.910000 14.185000  24.110000 ;
        RECT 13.985000  24.340000 14.185000  24.540000 ;
        RECT 13.985000  24.770000 14.185000  24.970000 ;
        RECT 13.985000  25.200000 14.185000  25.400000 ;
        RECT 13.985000  25.630000 14.185000  25.830000 ;
        RECT 13.985000  26.060000 14.185000  26.260000 ;
        RECT 13.985000  26.490000 14.185000  26.690000 ;
        RECT 13.985000  26.920000 14.185000  27.120000 ;
        RECT 13.985000  27.350000 14.185000  27.550000 ;
        RECT 13.985000  27.780000 14.185000  27.980000 ;
        RECT 13.985000  28.210000 14.185000  28.410000 ;
        RECT 14.390000  23.910000 14.590000  24.110000 ;
        RECT 14.390000  24.340000 14.590000  24.540000 ;
        RECT 14.390000  24.770000 14.590000  24.970000 ;
        RECT 14.390000  25.200000 14.590000  25.400000 ;
        RECT 14.390000  25.630000 14.590000  25.830000 ;
        RECT 14.390000  26.060000 14.590000  26.260000 ;
        RECT 14.390000  26.490000 14.590000  26.690000 ;
        RECT 14.390000  26.920000 14.590000  27.120000 ;
        RECT 14.390000  27.350000 14.590000  27.550000 ;
        RECT 14.390000  27.780000 14.590000  27.980000 ;
        RECT 14.390000  28.210000 14.590000  28.410000 ;
        RECT 14.795000  23.910000 14.995000  24.110000 ;
        RECT 14.795000  24.340000 14.995000  24.540000 ;
        RECT 14.795000  24.770000 14.995000  24.970000 ;
        RECT 14.795000  25.200000 14.995000  25.400000 ;
        RECT 14.795000  25.630000 14.995000  25.830000 ;
        RECT 14.795000  26.060000 14.995000  26.260000 ;
        RECT 14.795000  26.490000 14.995000  26.690000 ;
        RECT 14.795000  26.920000 14.995000  27.120000 ;
        RECT 14.795000  27.350000 14.995000  27.550000 ;
        RECT 14.795000  27.780000 14.995000  27.980000 ;
        RECT 14.795000  28.210000 14.995000  28.410000 ;
        RECT 15.200000  23.910000 15.400000  24.110000 ;
        RECT 15.200000  24.340000 15.400000  24.540000 ;
        RECT 15.200000  24.770000 15.400000  24.970000 ;
        RECT 15.200000  25.200000 15.400000  25.400000 ;
        RECT 15.200000  25.630000 15.400000  25.830000 ;
        RECT 15.200000  26.060000 15.400000  26.260000 ;
        RECT 15.200000  26.490000 15.400000  26.690000 ;
        RECT 15.200000  26.920000 15.400000  27.120000 ;
        RECT 15.200000  27.350000 15.400000  27.550000 ;
        RECT 15.200000  27.780000 15.400000  27.980000 ;
        RECT 15.200000  28.210000 15.400000  28.410000 ;
        RECT 15.605000  23.910000 15.805000  24.110000 ;
        RECT 15.605000  24.340000 15.805000  24.540000 ;
        RECT 15.605000  24.770000 15.805000  24.970000 ;
        RECT 15.605000  25.200000 15.805000  25.400000 ;
        RECT 15.605000  25.630000 15.805000  25.830000 ;
        RECT 15.605000  26.060000 15.805000  26.260000 ;
        RECT 15.605000  26.490000 15.805000  26.690000 ;
        RECT 15.605000  26.920000 15.805000  27.120000 ;
        RECT 15.605000  27.350000 15.805000  27.550000 ;
        RECT 15.605000  27.780000 15.805000  27.980000 ;
        RECT 15.605000  28.210000 15.805000  28.410000 ;
        RECT 16.010000  23.910000 16.210000  24.110000 ;
        RECT 16.010000  24.340000 16.210000  24.540000 ;
        RECT 16.010000  24.770000 16.210000  24.970000 ;
        RECT 16.010000  25.200000 16.210000  25.400000 ;
        RECT 16.010000  25.630000 16.210000  25.830000 ;
        RECT 16.010000  26.060000 16.210000  26.260000 ;
        RECT 16.010000  26.490000 16.210000  26.690000 ;
        RECT 16.010000  26.920000 16.210000  27.120000 ;
        RECT 16.010000  27.350000 16.210000  27.550000 ;
        RECT 16.010000  27.780000 16.210000  27.980000 ;
        RECT 16.010000  28.210000 16.210000  28.410000 ;
        RECT 16.415000  23.910000 16.615000  24.110000 ;
        RECT 16.415000  24.340000 16.615000  24.540000 ;
        RECT 16.415000  24.770000 16.615000  24.970000 ;
        RECT 16.415000  25.200000 16.615000  25.400000 ;
        RECT 16.415000  25.630000 16.615000  25.830000 ;
        RECT 16.415000  26.060000 16.615000  26.260000 ;
        RECT 16.415000  26.490000 16.615000  26.690000 ;
        RECT 16.415000  26.920000 16.615000  27.120000 ;
        RECT 16.415000  27.350000 16.615000  27.550000 ;
        RECT 16.415000  27.780000 16.615000  27.980000 ;
        RECT 16.415000  28.210000 16.615000  28.410000 ;
        RECT 16.820000  23.910000 17.020000  24.110000 ;
        RECT 16.820000  24.340000 17.020000  24.540000 ;
        RECT 16.820000  24.770000 17.020000  24.970000 ;
        RECT 16.820000  25.200000 17.020000  25.400000 ;
        RECT 16.820000  25.630000 17.020000  25.830000 ;
        RECT 16.820000  26.060000 17.020000  26.260000 ;
        RECT 16.820000  26.490000 17.020000  26.690000 ;
        RECT 16.820000  26.920000 17.020000  27.120000 ;
        RECT 16.820000  27.350000 17.020000  27.550000 ;
        RECT 16.820000  27.780000 17.020000  27.980000 ;
        RECT 16.820000  28.210000 17.020000  28.410000 ;
        RECT 17.225000  23.910000 17.425000  24.110000 ;
        RECT 17.225000  24.340000 17.425000  24.540000 ;
        RECT 17.225000  24.770000 17.425000  24.970000 ;
        RECT 17.225000  25.200000 17.425000  25.400000 ;
        RECT 17.225000  25.630000 17.425000  25.830000 ;
        RECT 17.225000  26.060000 17.425000  26.260000 ;
        RECT 17.225000  26.490000 17.425000  26.690000 ;
        RECT 17.225000  26.920000 17.425000  27.120000 ;
        RECT 17.225000  27.350000 17.425000  27.550000 ;
        RECT 17.225000  27.780000 17.425000  27.980000 ;
        RECT 17.225000  28.210000 17.425000  28.410000 ;
        RECT 17.630000  23.910000 17.830000  24.110000 ;
        RECT 17.630000  24.340000 17.830000  24.540000 ;
        RECT 17.630000  24.770000 17.830000  24.970000 ;
        RECT 17.630000  25.200000 17.830000  25.400000 ;
        RECT 17.630000  25.630000 17.830000  25.830000 ;
        RECT 17.630000  26.060000 17.830000  26.260000 ;
        RECT 17.630000  26.490000 17.830000  26.690000 ;
        RECT 17.630000  26.920000 17.830000  27.120000 ;
        RECT 17.630000  27.350000 17.830000  27.550000 ;
        RECT 17.630000  27.780000 17.830000  27.980000 ;
        RECT 17.630000  28.210000 17.830000  28.410000 ;
        RECT 18.035000  23.910000 18.235000  24.110000 ;
        RECT 18.035000  24.340000 18.235000  24.540000 ;
        RECT 18.035000  24.770000 18.235000  24.970000 ;
        RECT 18.035000  25.200000 18.235000  25.400000 ;
        RECT 18.035000  25.630000 18.235000  25.830000 ;
        RECT 18.035000  26.060000 18.235000  26.260000 ;
        RECT 18.035000  26.490000 18.235000  26.690000 ;
        RECT 18.035000  26.920000 18.235000  27.120000 ;
        RECT 18.035000  27.350000 18.235000  27.550000 ;
        RECT 18.035000  27.780000 18.235000  27.980000 ;
        RECT 18.035000  28.210000 18.235000  28.410000 ;
        RECT 18.440000  23.910000 18.640000  24.110000 ;
        RECT 18.440000  24.340000 18.640000  24.540000 ;
        RECT 18.440000  24.770000 18.640000  24.970000 ;
        RECT 18.440000  25.200000 18.640000  25.400000 ;
        RECT 18.440000  25.630000 18.640000  25.830000 ;
        RECT 18.440000  26.060000 18.640000  26.260000 ;
        RECT 18.440000  26.490000 18.640000  26.690000 ;
        RECT 18.440000  26.920000 18.640000  27.120000 ;
        RECT 18.440000  27.350000 18.640000  27.550000 ;
        RECT 18.440000  27.780000 18.640000  27.980000 ;
        RECT 18.440000  28.210000 18.640000  28.410000 ;
        RECT 18.845000  23.910000 19.045000  24.110000 ;
        RECT 18.845000  24.340000 19.045000  24.540000 ;
        RECT 18.845000  24.770000 19.045000  24.970000 ;
        RECT 18.845000  25.200000 19.045000  25.400000 ;
        RECT 18.845000  25.630000 19.045000  25.830000 ;
        RECT 18.845000  26.060000 19.045000  26.260000 ;
        RECT 18.845000  26.490000 19.045000  26.690000 ;
        RECT 18.845000  26.920000 19.045000  27.120000 ;
        RECT 18.845000  27.350000 19.045000  27.550000 ;
        RECT 18.845000  27.780000 19.045000  27.980000 ;
        RECT 18.845000  28.210000 19.045000  28.410000 ;
        RECT 19.250000  23.910000 19.450000  24.110000 ;
        RECT 19.250000  24.340000 19.450000  24.540000 ;
        RECT 19.250000  24.770000 19.450000  24.970000 ;
        RECT 19.250000  25.200000 19.450000  25.400000 ;
        RECT 19.250000  25.630000 19.450000  25.830000 ;
        RECT 19.250000  26.060000 19.450000  26.260000 ;
        RECT 19.250000  26.490000 19.450000  26.690000 ;
        RECT 19.250000  26.920000 19.450000  27.120000 ;
        RECT 19.250000  27.350000 19.450000  27.550000 ;
        RECT 19.250000  27.780000 19.450000  27.980000 ;
        RECT 19.250000  28.210000 19.450000  28.410000 ;
        RECT 19.655000  23.910000 19.855000  24.110000 ;
        RECT 19.655000  24.340000 19.855000  24.540000 ;
        RECT 19.655000  24.770000 19.855000  24.970000 ;
        RECT 19.655000  25.200000 19.855000  25.400000 ;
        RECT 19.655000  25.630000 19.855000  25.830000 ;
        RECT 19.655000  26.060000 19.855000  26.260000 ;
        RECT 19.655000  26.490000 19.855000  26.690000 ;
        RECT 19.655000  26.920000 19.855000  27.120000 ;
        RECT 19.655000  27.350000 19.855000  27.550000 ;
        RECT 19.655000  27.780000 19.855000  27.980000 ;
        RECT 19.655000  28.210000 19.855000  28.410000 ;
        RECT 20.060000  23.910000 20.260000  24.110000 ;
        RECT 20.060000  24.340000 20.260000  24.540000 ;
        RECT 20.060000  24.770000 20.260000  24.970000 ;
        RECT 20.060000  25.200000 20.260000  25.400000 ;
        RECT 20.060000  25.630000 20.260000  25.830000 ;
        RECT 20.060000  26.060000 20.260000  26.260000 ;
        RECT 20.060000  26.490000 20.260000  26.690000 ;
        RECT 20.060000  26.920000 20.260000  27.120000 ;
        RECT 20.060000  27.350000 20.260000  27.550000 ;
        RECT 20.060000  27.780000 20.260000  27.980000 ;
        RECT 20.060000  28.210000 20.260000  28.410000 ;
        RECT 20.465000  23.910000 20.665000  24.110000 ;
        RECT 20.465000  24.340000 20.665000  24.540000 ;
        RECT 20.465000  24.770000 20.665000  24.970000 ;
        RECT 20.465000  25.200000 20.665000  25.400000 ;
        RECT 20.465000  25.630000 20.665000  25.830000 ;
        RECT 20.465000  26.060000 20.665000  26.260000 ;
        RECT 20.465000  26.490000 20.665000  26.690000 ;
        RECT 20.465000  26.920000 20.665000  27.120000 ;
        RECT 20.465000  27.350000 20.665000  27.550000 ;
        RECT 20.465000  27.780000 20.665000  27.980000 ;
        RECT 20.465000  28.210000 20.665000  28.410000 ;
        RECT 20.870000  23.910000 21.070000  24.110000 ;
        RECT 20.870000  24.340000 21.070000  24.540000 ;
        RECT 20.870000  24.770000 21.070000  24.970000 ;
        RECT 20.870000  25.200000 21.070000  25.400000 ;
        RECT 20.870000  25.630000 21.070000  25.830000 ;
        RECT 20.870000  26.060000 21.070000  26.260000 ;
        RECT 20.870000  26.490000 21.070000  26.690000 ;
        RECT 20.870000  26.920000 21.070000  27.120000 ;
        RECT 20.870000  27.350000 21.070000  27.550000 ;
        RECT 20.870000  27.780000 21.070000  27.980000 ;
        RECT 20.870000  28.210000 21.070000  28.410000 ;
        RECT 21.275000  23.910000 21.475000  24.110000 ;
        RECT 21.275000  24.340000 21.475000  24.540000 ;
        RECT 21.275000  24.770000 21.475000  24.970000 ;
        RECT 21.275000  25.200000 21.475000  25.400000 ;
        RECT 21.275000  25.630000 21.475000  25.830000 ;
        RECT 21.275000  26.060000 21.475000  26.260000 ;
        RECT 21.275000  26.490000 21.475000  26.690000 ;
        RECT 21.275000  26.920000 21.475000  27.120000 ;
        RECT 21.275000  27.350000 21.475000  27.550000 ;
        RECT 21.275000  27.780000 21.475000  27.980000 ;
        RECT 21.275000  28.210000 21.475000  28.410000 ;
        RECT 21.680000  23.910000 21.880000  24.110000 ;
        RECT 21.680000  24.340000 21.880000  24.540000 ;
        RECT 21.680000  24.770000 21.880000  24.970000 ;
        RECT 21.680000  25.200000 21.880000  25.400000 ;
        RECT 21.680000  25.630000 21.880000  25.830000 ;
        RECT 21.680000  26.060000 21.880000  26.260000 ;
        RECT 21.680000  26.490000 21.880000  26.690000 ;
        RECT 21.680000  26.920000 21.880000  27.120000 ;
        RECT 21.680000  27.350000 21.880000  27.550000 ;
        RECT 21.680000  27.780000 21.880000  27.980000 ;
        RECT 21.680000  28.210000 21.880000  28.410000 ;
        RECT 22.085000  23.910000 22.285000  24.110000 ;
        RECT 22.085000  24.340000 22.285000  24.540000 ;
        RECT 22.085000  24.770000 22.285000  24.970000 ;
        RECT 22.085000  25.200000 22.285000  25.400000 ;
        RECT 22.085000  25.630000 22.285000  25.830000 ;
        RECT 22.085000  26.060000 22.285000  26.260000 ;
        RECT 22.085000  26.490000 22.285000  26.690000 ;
        RECT 22.085000  26.920000 22.285000  27.120000 ;
        RECT 22.085000  27.350000 22.285000  27.550000 ;
        RECT 22.085000  27.780000 22.285000  27.980000 ;
        RECT 22.085000  28.210000 22.285000  28.410000 ;
        RECT 22.490000  23.910000 22.690000  24.110000 ;
        RECT 22.490000  24.340000 22.690000  24.540000 ;
        RECT 22.490000  24.770000 22.690000  24.970000 ;
        RECT 22.490000  25.200000 22.690000  25.400000 ;
        RECT 22.490000  25.630000 22.690000  25.830000 ;
        RECT 22.490000  26.060000 22.690000  26.260000 ;
        RECT 22.490000  26.490000 22.690000  26.690000 ;
        RECT 22.490000  26.920000 22.690000  27.120000 ;
        RECT 22.490000  27.350000 22.690000  27.550000 ;
        RECT 22.490000  27.780000 22.690000  27.980000 ;
        RECT 22.490000  28.210000 22.690000  28.410000 ;
        RECT 22.895000  23.910000 23.095000  24.110000 ;
        RECT 22.895000  24.340000 23.095000  24.540000 ;
        RECT 22.895000  24.770000 23.095000  24.970000 ;
        RECT 22.895000  25.200000 23.095000  25.400000 ;
        RECT 22.895000  25.630000 23.095000  25.830000 ;
        RECT 22.895000  26.060000 23.095000  26.260000 ;
        RECT 22.895000  26.490000 23.095000  26.690000 ;
        RECT 22.895000  26.920000 23.095000  27.120000 ;
        RECT 22.895000  27.350000 23.095000  27.550000 ;
        RECT 22.895000  27.780000 23.095000  27.980000 ;
        RECT 22.895000  28.210000 23.095000  28.410000 ;
        RECT 23.300000  23.910000 23.500000  24.110000 ;
        RECT 23.300000  24.340000 23.500000  24.540000 ;
        RECT 23.300000  24.770000 23.500000  24.970000 ;
        RECT 23.300000  25.200000 23.500000  25.400000 ;
        RECT 23.300000  25.630000 23.500000  25.830000 ;
        RECT 23.300000  26.060000 23.500000  26.260000 ;
        RECT 23.300000  26.490000 23.500000  26.690000 ;
        RECT 23.300000  26.920000 23.500000  27.120000 ;
        RECT 23.300000  27.350000 23.500000  27.550000 ;
        RECT 23.300000  27.780000 23.500000  27.980000 ;
        RECT 23.300000  28.210000 23.500000  28.410000 ;
        RECT 23.705000  23.910000 23.905000  24.110000 ;
        RECT 23.705000  24.340000 23.905000  24.540000 ;
        RECT 23.705000  24.770000 23.905000  24.970000 ;
        RECT 23.705000  25.200000 23.905000  25.400000 ;
        RECT 23.705000  25.630000 23.905000  25.830000 ;
        RECT 23.705000  26.060000 23.905000  26.260000 ;
        RECT 23.705000  26.490000 23.905000  26.690000 ;
        RECT 23.705000  26.920000 23.905000  27.120000 ;
        RECT 23.705000  27.350000 23.905000  27.550000 ;
        RECT 23.705000  27.780000 23.905000  27.980000 ;
        RECT 23.705000  28.210000 23.905000  28.410000 ;
        RECT 24.110000  23.910000 24.310000  24.110000 ;
        RECT 24.110000  24.340000 24.310000  24.540000 ;
        RECT 24.110000  24.770000 24.310000  24.970000 ;
        RECT 24.110000  25.200000 24.310000  25.400000 ;
        RECT 24.110000  25.630000 24.310000  25.830000 ;
        RECT 24.110000  26.060000 24.310000  26.260000 ;
        RECT 24.110000  26.490000 24.310000  26.690000 ;
        RECT 24.110000  26.920000 24.310000  27.120000 ;
        RECT 24.110000  27.350000 24.310000  27.550000 ;
        RECT 24.110000  27.780000 24.310000  27.980000 ;
        RECT 24.110000  28.210000 24.310000  28.410000 ;
        RECT 50.845000  23.910000 51.045000  24.110000 ;
        RECT 50.845000  24.340000 51.045000  24.540000 ;
        RECT 50.845000  24.770000 51.045000  24.970000 ;
        RECT 50.845000  25.200000 51.045000  25.400000 ;
        RECT 50.845000  25.630000 51.045000  25.830000 ;
        RECT 50.845000  26.060000 51.045000  26.260000 ;
        RECT 50.845000  26.490000 51.045000  26.690000 ;
        RECT 50.845000  26.920000 51.045000  27.120000 ;
        RECT 50.845000  27.350000 51.045000  27.550000 ;
        RECT 50.845000  27.780000 51.045000  27.980000 ;
        RECT 50.845000  28.210000 51.045000  28.410000 ;
        RECT 51.255000  23.910000 51.455000  24.110000 ;
        RECT 51.255000  24.340000 51.455000  24.540000 ;
        RECT 51.255000  24.770000 51.455000  24.970000 ;
        RECT 51.255000  25.200000 51.455000  25.400000 ;
        RECT 51.255000  25.630000 51.455000  25.830000 ;
        RECT 51.255000  26.060000 51.455000  26.260000 ;
        RECT 51.255000  26.490000 51.455000  26.690000 ;
        RECT 51.255000  26.920000 51.455000  27.120000 ;
        RECT 51.255000  27.350000 51.455000  27.550000 ;
        RECT 51.255000  27.780000 51.455000  27.980000 ;
        RECT 51.255000  28.210000 51.455000  28.410000 ;
        RECT 51.665000  23.910000 51.865000  24.110000 ;
        RECT 51.665000  24.340000 51.865000  24.540000 ;
        RECT 51.665000  24.770000 51.865000  24.970000 ;
        RECT 51.665000  25.200000 51.865000  25.400000 ;
        RECT 51.665000  25.630000 51.865000  25.830000 ;
        RECT 51.665000  26.060000 51.865000  26.260000 ;
        RECT 51.665000  26.490000 51.865000  26.690000 ;
        RECT 51.665000  26.920000 51.865000  27.120000 ;
        RECT 51.665000  27.350000 51.865000  27.550000 ;
        RECT 51.665000  27.780000 51.865000  27.980000 ;
        RECT 51.665000  28.210000 51.865000  28.410000 ;
        RECT 52.075000  23.910000 52.275000  24.110000 ;
        RECT 52.075000  24.340000 52.275000  24.540000 ;
        RECT 52.075000  24.770000 52.275000  24.970000 ;
        RECT 52.075000  25.200000 52.275000  25.400000 ;
        RECT 52.075000  25.630000 52.275000  25.830000 ;
        RECT 52.075000  26.060000 52.275000  26.260000 ;
        RECT 52.075000  26.490000 52.275000  26.690000 ;
        RECT 52.075000  26.920000 52.275000  27.120000 ;
        RECT 52.075000  27.350000 52.275000  27.550000 ;
        RECT 52.075000  27.780000 52.275000  27.980000 ;
        RECT 52.075000  28.210000 52.275000  28.410000 ;
        RECT 52.485000  23.910000 52.685000  24.110000 ;
        RECT 52.485000  24.340000 52.685000  24.540000 ;
        RECT 52.485000  24.770000 52.685000  24.970000 ;
        RECT 52.485000  25.200000 52.685000  25.400000 ;
        RECT 52.485000  25.630000 52.685000  25.830000 ;
        RECT 52.485000  26.060000 52.685000  26.260000 ;
        RECT 52.485000  26.490000 52.685000  26.690000 ;
        RECT 52.485000  26.920000 52.685000  27.120000 ;
        RECT 52.485000  27.350000 52.685000  27.550000 ;
        RECT 52.485000  27.780000 52.685000  27.980000 ;
        RECT 52.485000  28.210000 52.685000  28.410000 ;
        RECT 52.895000  23.910000 53.095000  24.110000 ;
        RECT 52.895000  24.340000 53.095000  24.540000 ;
        RECT 52.895000  24.770000 53.095000  24.970000 ;
        RECT 52.895000  25.200000 53.095000  25.400000 ;
        RECT 52.895000  25.630000 53.095000  25.830000 ;
        RECT 52.895000  26.060000 53.095000  26.260000 ;
        RECT 52.895000  26.490000 53.095000  26.690000 ;
        RECT 52.895000  26.920000 53.095000  27.120000 ;
        RECT 52.895000  27.350000 53.095000  27.550000 ;
        RECT 52.895000  27.780000 53.095000  27.980000 ;
        RECT 52.895000  28.210000 53.095000  28.410000 ;
        RECT 53.305000  23.910000 53.505000  24.110000 ;
        RECT 53.305000  24.340000 53.505000  24.540000 ;
        RECT 53.305000  24.770000 53.505000  24.970000 ;
        RECT 53.305000  25.200000 53.505000  25.400000 ;
        RECT 53.305000  25.630000 53.505000  25.830000 ;
        RECT 53.305000  26.060000 53.505000  26.260000 ;
        RECT 53.305000  26.490000 53.505000  26.690000 ;
        RECT 53.305000  26.920000 53.505000  27.120000 ;
        RECT 53.305000  27.350000 53.505000  27.550000 ;
        RECT 53.305000  27.780000 53.505000  27.980000 ;
        RECT 53.305000  28.210000 53.505000  28.410000 ;
        RECT 53.715000  23.910000 53.915000  24.110000 ;
        RECT 53.715000  24.340000 53.915000  24.540000 ;
        RECT 53.715000  24.770000 53.915000  24.970000 ;
        RECT 53.715000  25.200000 53.915000  25.400000 ;
        RECT 53.715000  25.630000 53.915000  25.830000 ;
        RECT 53.715000  26.060000 53.915000  26.260000 ;
        RECT 53.715000  26.490000 53.915000  26.690000 ;
        RECT 53.715000  26.920000 53.915000  27.120000 ;
        RECT 53.715000  27.350000 53.915000  27.550000 ;
        RECT 53.715000  27.780000 53.915000  27.980000 ;
        RECT 53.715000  28.210000 53.915000  28.410000 ;
        RECT 54.125000  23.910000 54.325000  24.110000 ;
        RECT 54.125000  24.340000 54.325000  24.540000 ;
        RECT 54.125000  24.770000 54.325000  24.970000 ;
        RECT 54.125000  25.200000 54.325000  25.400000 ;
        RECT 54.125000  25.630000 54.325000  25.830000 ;
        RECT 54.125000  26.060000 54.325000  26.260000 ;
        RECT 54.125000  26.490000 54.325000  26.690000 ;
        RECT 54.125000  26.920000 54.325000  27.120000 ;
        RECT 54.125000  27.350000 54.325000  27.550000 ;
        RECT 54.125000  27.780000 54.325000  27.980000 ;
        RECT 54.125000  28.210000 54.325000  28.410000 ;
        RECT 54.535000  23.910000 54.735000  24.110000 ;
        RECT 54.535000  24.340000 54.735000  24.540000 ;
        RECT 54.535000  24.770000 54.735000  24.970000 ;
        RECT 54.535000  25.200000 54.735000  25.400000 ;
        RECT 54.535000  25.630000 54.735000  25.830000 ;
        RECT 54.535000  26.060000 54.735000  26.260000 ;
        RECT 54.535000  26.490000 54.735000  26.690000 ;
        RECT 54.535000  26.920000 54.735000  27.120000 ;
        RECT 54.535000  27.350000 54.735000  27.550000 ;
        RECT 54.535000  27.780000 54.735000  27.980000 ;
        RECT 54.535000  28.210000 54.735000  28.410000 ;
        RECT 54.945000  23.910000 55.145000  24.110000 ;
        RECT 54.945000  24.340000 55.145000  24.540000 ;
        RECT 54.945000  24.770000 55.145000  24.970000 ;
        RECT 54.945000  25.200000 55.145000  25.400000 ;
        RECT 54.945000  25.630000 55.145000  25.830000 ;
        RECT 54.945000  26.060000 55.145000  26.260000 ;
        RECT 54.945000  26.490000 55.145000  26.690000 ;
        RECT 54.945000  26.920000 55.145000  27.120000 ;
        RECT 54.945000  27.350000 55.145000  27.550000 ;
        RECT 54.945000  27.780000 55.145000  27.980000 ;
        RECT 54.945000  28.210000 55.145000  28.410000 ;
        RECT 55.355000  23.910000 55.555000  24.110000 ;
        RECT 55.355000  24.340000 55.555000  24.540000 ;
        RECT 55.355000  24.770000 55.555000  24.970000 ;
        RECT 55.355000  25.200000 55.555000  25.400000 ;
        RECT 55.355000  25.630000 55.555000  25.830000 ;
        RECT 55.355000  26.060000 55.555000  26.260000 ;
        RECT 55.355000  26.490000 55.555000  26.690000 ;
        RECT 55.355000  26.920000 55.555000  27.120000 ;
        RECT 55.355000  27.350000 55.555000  27.550000 ;
        RECT 55.355000  27.780000 55.555000  27.980000 ;
        RECT 55.355000  28.210000 55.555000  28.410000 ;
        RECT 55.765000  23.910000 55.965000  24.110000 ;
        RECT 55.765000  24.340000 55.965000  24.540000 ;
        RECT 55.765000  24.770000 55.965000  24.970000 ;
        RECT 55.765000  25.200000 55.965000  25.400000 ;
        RECT 55.765000  25.630000 55.965000  25.830000 ;
        RECT 55.765000  26.060000 55.965000  26.260000 ;
        RECT 55.765000  26.490000 55.965000  26.690000 ;
        RECT 55.765000  26.920000 55.965000  27.120000 ;
        RECT 55.765000  27.350000 55.965000  27.550000 ;
        RECT 55.765000  27.780000 55.965000  27.980000 ;
        RECT 55.765000  28.210000 55.965000  28.410000 ;
        RECT 56.175000  23.910000 56.375000  24.110000 ;
        RECT 56.175000  24.340000 56.375000  24.540000 ;
        RECT 56.175000  24.770000 56.375000  24.970000 ;
        RECT 56.175000  25.200000 56.375000  25.400000 ;
        RECT 56.175000  25.630000 56.375000  25.830000 ;
        RECT 56.175000  26.060000 56.375000  26.260000 ;
        RECT 56.175000  26.490000 56.375000  26.690000 ;
        RECT 56.175000  26.920000 56.375000  27.120000 ;
        RECT 56.175000  27.350000 56.375000  27.550000 ;
        RECT 56.175000  27.780000 56.375000  27.980000 ;
        RECT 56.175000  28.210000 56.375000  28.410000 ;
        RECT 56.585000  23.910000 56.785000  24.110000 ;
        RECT 56.585000  24.340000 56.785000  24.540000 ;
        RECT 56.585000  24.770000 56.785000  24.970000 ;
        RECT 56.585000  25.200000 56.785000  25.400000 ;
        RECT 56.585000  25.630000 56.785000  25.830000 ;
        RECT 56.585000  26.060000 56.785000  26.260000 ;
        RECT 56.585000  26.490000 56.785000  26.690000 ;
        RECT 56.585000  26.920000 56.785000  27.120000 ;
        RECT 56.585000  27.350000 56.785000  27.550000 ;
        RECT 56.585000  27.780000 56.785000  27.980000 ;
        RECT 56.585000  28.210000 56.785000  28.410000 ;
        RECT 56.990000  23.910000 57.190000  24.110000 ;
        RECT 56.990000  24.340000 57.190000  24.540000 ;
        RECT 56.990000  24.770000 57.190000  24.970000 ;
        RECT 56.990000  25.200000 57.190000  25.400000 ;
        RECT 56.990000  25.630000 57.190000  25.830000 ;
        RECT 56.990000  26.060000 57.190000  26.260000 ;
        RECT 56.990000  26.490000 57.190000  26.690000 ;
        RECT 56.990000  26.920000 57.190000  27.120000 ;
        RECT 56.990000  27.350000 57.190000  27.550000 ;
        RECT 56.990000  27.780000 57.190000  27.980000 ;
        RECT 56.990000  28.210000 57.190000  28.410000 ;
        RECT 57.395000  23.910000 57.595000  24.110000 ;
        RECT 57.395000  24.340000 57.595000  24.540000 ;
        RECT 57.395000  24.770000 57.595000  24.970000 ;
        RECT 57.395000  25.200000 57.595000  25.400000 ;
        RECT 57.395000  25.630000 57.595000  25.830000 ;
        RECT 57.395000  26.060000 57.595000  26.260000 ;
        RECT 57.395000  26.490000 57.595000  26.690000 ;
        RECT 57.395000  26.920000 57.595000  27.120000 ;
        RECT 57.395000  27.350000 57.595000  27.550000 ;
        RECT 57.395000  27.780000 57.595000  27.980000 ;
        RECT 57.395000  28.210000 57.595000  28.410000 ;
        RECT 57.800000  23.910000 58.000000  24.110000 ;
        RECT 57.800000  24.340000 58.000000  24.540000 ;
        RECT 57.800000  24.770000 58.000000  24.970000 ;
        RECT 57.800000  25.200000 58.000000  25.400000 ;
        RECT 57.800000  25.630000 58.000000  25.830000 ;
        RECT 57.800000  26.060000 58.000000  26.260000 ;
        RECT 57.800000  26.490000 58.000000  26.690000 ;
        RECT 57.800000  26.920000 58.000000  27.120000 ;
        RECT 57.800000  27.350000 58.000000  27.550000 ;
        RECT 57.800000  27.780000 58.000000  27.980000 ;
        RECT 57.800000  28.210000 58.000000  28.410000 ;
        RECT 58.205000  23.910000 58.405000  24.110000 ;
        RECT 58.205000  24.340000 58.405000  24.540000 ;
        RECT 58.205000  24.770000 58.405000  24.970000 ;
        RECT 58.205000  25.200000 58.405000  25.400000 ;
        RECT 58.205000  25.630000 58.405000  25.830000 ;
        RECT 58.205000  26.060000 58.405000  26.260000 ;
        RECT 58.205000  26.490000 58.405000  26.690000 ;
        RECT 58.205000  26.920000 58.405000  27.120000 ;
        RECT 58.205000  27.350000 58.405000  27.550000 ;
        RECT 58.205000  27.780000 58.405000  27.980000 ;
        RECT 58.205000  28.210000 58.405000  28.410000 ;
        RECT 58.610000  23.910000 58.810000  24.110000 ;
        RECT 58.610000  24.340000 58.810000  24.540000 ;
        RECT 58.610000  24.770000 58.810000  24.970000 ;
        RECT 58.610000  25.200000 58.810000  25.400000 ;
        RECT 58.610000  25.630000 58.810000  25.830000 ;
        RECT 58.610000  26.060000 58.810000  26.260000 ;
        RECT 58.610000  26.490000 58.810000  26.690000 ;
        RECT 58.610000  26.920000 58.810000  27.120000 ;
        RECT 58.610000  27.350000 58.810000  27.550000 ;
        RECT 58.610000  27.780000 58.810000  27.980000 ;
        RECT 58.610000  28.210000 58.810000  28.410000 ;
        RECT 59.015000  23.910000 59.215000  24.110000 ;
        RECT 59.015000  24.340000 59.215000  24.540000 ;
        RECT 59.015000  24.770000 59.215000  24.970000 ;
        RECT 59.015000  25.200000 59.215000  25.400000 ;
        RECT 59.015000  25.630000 59.215000  25.830000 ;
        RECT 59.015000  26.060000 59.215000  26.260000 ;
        RECT 59.015000  26.490000 59.215000  26.690000 ;
        RECT 59.015000  26.920000 59.215000  27.120000 ;
        RECT 59.015000  27.350000 59.215000  27.550000 ;
        RECT 59.015000  27.780000 59.215000  27.980000 ;
        RECT 59.015000  28.210000 59.215000  28.410000 ;
        RECT 59.420000  23.910000 59.620000  24.110000 ;
        RECT 59.420000  24.340000 59.620000  24.540000 ;
        RECT 59.420000  24.770000 59.620000  24.970000 ;
        RECT 59.420000  25.200000 59.620000  25.400000 ;
        RECT 59.420000  25.630000 59.620000  25.830000 ;
        RECT 59.420000  26.060000 59.620000  26.260000 ;
        RECT 59.420000  26.490000 59.620000  26.690000 ;
        RECT 59.420000  26.920000 59.620000  27.120000 ;
        RECT 59.420000  27.350000 59.620000  27.550000 ;
        RECT 59.420000  27.780000 59.620000  27.980000 ;
        RECT 59.420000  28.210000 59.620000  28.410000 ;
        RECT 59.825000  23.910000 60.025000  24.110000 ;
        RECT 59.825000  24.340000 60.025000  24.540000 ;
        RECT 59.825000  24.770000 60.025000  24.970000 ;
        RECT 59.825000  25.200000 60.025000  25.400000 ;
        RECT 59.825000  25.630000 60.025000  25.830000 ;
        RECT 59.825000  26.060000 60.025000  26.260000 ;
        RECT 59.825000  26.490000 60.025000  26.690000 ;
        RECT 59.825000  26.920000 60.025000  27.120000 ;
        RECT 59.825000  27.350000 60.025000  27.550000 ;
        RECT 59.825000  27.780000 60.025000  27.980000 ;
        RECT 59.825000  28.210000 60.025000  28.410000 ;
        RECT 60.230000  23.910000 60.430000  24.110000 ;
        RECT 60.230000  24.340000 60.430000  24.540000 ;
        RECT 60.230000  24.770000 60.430000  24.970000 ;
        RECT 60.230000  25.200000 60.430000  25.400000 ;
        RECT 60.230000  25.630000 60.430000  25.830000 ;
        RECT 60.230000  26.060000 60.430000  26.260000 ;
        RECT 60.230000  26.490000 60.430000  26.690000 ;
        RECT 60.230000  26.920000 60.430000  27.120000 ;
        RECT 60.230000  27.350000 60.430000  27.550000 ;
        RECT 60.230000  27.780000 60.430000  27.980000 ;
        RECT 60.230000  28.210000 60.430000  28.410000 ;
        RECT 60.635000  23.910000 60.835000  24.110000 ;
        RECT 60.635000  24.340000 60.835000  24.540000 ;
        RECT 60.635000  24.770000 60.835000  24.970000 ;
        RECT 60.635000  25.200000 60.835000  25.400000 ;
        RECT 60.635000  25.630000 60.835000  25.830000 ;
        RECT 60.635000  26.060000 60.835000  26.260000 ;
        RECT 60.635000  26.490000 60.835000  26.690000 ;
        RECT 60.635000  26.920000 60.835000  27.120000 ;
        RECT 60.635000  27.350000 60.835000  27.550000 ;
        RECT 60.635000  27.780000 60.835000  27.980000 ;
        RECT 60.635000  28.210000 60.835000  28.410000 ;
        RECT 61.040000  23.910000 61.240000  24.110000 ;
        RECT 61.040000  24.340000 61.240000  24.540000 ;
        RECT 61.040000  24.770000 61.240000  24.970000 ;
        RECT 61.040000  25.200000 61.240000  25.400000 ;
        RECT 61.040000  25.630000 61.240000  25.830000 ;
        RECT 61.040000  26.060000 61.240000  26.260000 ;
        RECT 61.040000  26.490000 61.240000  26.690000 ;
        RECT 61.040000  26.920000 61.240000  27.120000 ;
        RECT 61.040000  27.350000 61.240000  27.550000 ;
        RECT 61.040000  27.780000 61.240000  27.980000 ;
        RECT 61.040000  28.210000 61.240000  28.410000 ;
        RECT 61.445000  23.910000 61.645000  24.110000 ;
        RECT 61.445000  24.340000 61.645000  24.540000 ;
        RECT 61.445000  24.770000 61.645000  24.970000 ;
        RECT 61.445000  25.200000 61.645000  25.400000 ;
        RECT 61.445000  25.630000 61.645000  25.830000 ;
        RECT 61.445000  26.060000 61.645000  26.260000 ;
        RECT 61.445000  26.490000 61.645000  26.690000 ;
        RECT 61.445000  26.920000 61.645000  27.120000 ;
        RECT 61.445000  27.350000 61.645000  27.550000 ;
        RECT 61.445000  27.780000 61.645000  27.980000 ;
        RECT 61.445000  28.210000 61.645000  28.410000 ;
        RECT 61.850000  23.910000 62.050000  24.110000 ;
        RECT 61.850000  24.340000 62.050000  24.540000 ;
        RECT 61.850000  24.770000 62.050000  24.970000 ;
        RECT 61.850000  25.200000 62.050000  25.400000 ;
        RECT 61.850000  25.630000 62.050000  25.830000 ;
        RECT 61.850000  26.060000 62.050000  26.260000 ;
        RECT 61.850000  26.490000 62.050000  26.690000 ;
        RECT 61.850000  26.920000 62.050000  27.120000 ;
        RECT 61.850000  27.350000 62.050000  27.550000 ;
        RECT 61.850000  27.780000 62.050000  27.980000 ;
        RECT 61.850000  28.210000 62.050000  28.410000 ;
        RECT 62.140000 173.900000 62.340000 174.100000 ;
        RECT 62.140000 174.300000 62.340000 174.500000 ;
        RECT 62.140000 174.700000 62.340000 174.900000 ;
        RECT 62.140000 175.100000 62.340000 175.300000 ;
        RECT 62.140000 175.500000 62.340000 175.700000 ;
        RECT 62.140000 175.900000 62.340000 176.100000 ;
        RECT 62.140000 176.300000 62.340000 176.500000 ;
        RECT 62.140000 176.700000 62.340000 176.900000 ;
        RECT 62.140000 177.100000 62.340000 177.300000 ;
        RECT 62.140000 177.500000 62.340000 177.700000 ;
        RECT 62.140000 177.900000 62.340000 178.100000 ;
        RECT 62.140000 178.300000 62.340000 178.500000 ;
        RECT 62.140000 178.700000 62.340000 178.900000 ;
        RECT 62.140000 179.100000 62.340000 179.300000 ;
        RECT 62.140000 179.500000 62.340000 179.700000 ;
        RECT 62.140000 179.900000 62.340000 180.100000 ;
        RECT 62.140000 180.300000 62.340000 180.500000 ;
        RECT 62.140000 180.700000 62.340000 180.900000 ;
        RECT 62.140000 181.100000 62.340000 181.300000 ;
        RECT 62.140000 181.505000 62.340000 181.705000 ;
        RECT 62.140000 181.910000 62.340000 182.110000 ;
        RECT 62.140000 182.315000 62.340000 182.515000 ;
        RECT 62.140000 182.720000 62.340000 182.920000 ;
        RECT 62.140000 183.125000 62.340000 183.325000 ;
        RECT 62.140000 183.530000 62.340000 183.730000 ;
        RECT 62.140000 183.935000 62.340000 184.135000 ;
        RECT 62.140000 184.340000 62.340000 184.540000 ;
        RECT 62.140000 184.745000 62.340000 184.945000 ;
        RECT 62.140000 185.150000 62.340000 185.350000 ;
        RECT 62.140000 185.555000 62.340000 185.755000 ;
        RECT 62.140000 185.960000 62.340000 186.160000 ;
        RECT 62.140000 186.365000 62.340000 186.565000 ;
        RECT 62.140000 186.770000 62.340000 186.970000 ;
        RECT 62.140000 187.175000 62.340000 187.375000 ;
        RECT 62.140000 187.580000 62.340000 187.780000 ;
        RECT 62.140000 187.985000 62.340000 188.185000 ;
        RECT 62.140000 188.390000 62.340000 188.590000 ;
        RECT 62.140000 188.795000 62.340000 188.995000 ;
        RECT 62.140000 189.200000 62.340000 189.400000 ;
        RECT 62.140000 189.605000 62.340000 189.805000 ;
        RECT 62.140000 190.010000 62.340000 190.210000 ;
        RECT 62.140000 190.415000 62.340000 190.615000 ;
        RECT 62.140000 190.820000 62.340000 191.020000 ;
        RECT 62.140000 191.225000 62.340000 191.425000 ;
        RECT 62.140000 191.630000 62.340000 191.830000 ;
        RECT 62.140000 192.035000 62.340000 192.235000 ;
        RECT 62.140000 192.440000 62.340000 192.640000 ;
        RECT 62.140000 192.845000 62.340000 193.045000 ;
        RECT 62.140000 193.250000 62.340000 193.450000 ;
        RECT 62.140000 193.655000 62.340000 193.855000 ;
        RECT 62.140000 194.060000 62.340000 194.260000 ;
        RECT 62.140000 194.465000 62.340000 194.665000 ;
        RECT 62.140000 194.870000 62.340000 195.070000 ;
        RECT 62.140000 195.275000 62.340000 195.475000 ;
        RECT 62.140000 195.680000 62.340000 195.880000 ;
        RECT 62.140000 196.085000 62.340000 196.285000 ;
        RECT 62.140000 196.490000 62.340000 196.690000 ;
        RECT 62.140000 196.895000 62.340000 197.095000 ;
        RECT 62.140000 197.300000 62.340000 197.500000 ;
        RECT 62.140000 197.705000 62.340000 197.905000 ;
        RECT 62.255000  23.910000 62.455000  24.110000 ;
        RECT 62.255000  24.340000 62.455000  24.540000 ;
        RECT 62.255000  24.770000 62.455000  24.970000 ;
        RECT 62.255000  25.200000 62.455000  25.400000 ;
        RECT 62.255000  25.630000 62.455000  25.830000 ;
        RECT 62.255000  26.060000 62.455000  26.260000 ;
        RECT 62.255000  26.490000 62.455000  26.690000 ;
        RECT 62.255000  26.920000 62.455000  27.120000 ;
        RECT 62.255000  27.350000 62.455000  27.550000 ;
        RECT 62.255000  27.780000 62.455000  27.980000 ;
        RECT 62.255000  28.210000 62.455000  28.410000 ;
        RECT 62.550000 173.900000 62.750000 174.100000 ;
        RECT 62.550000 174.300000 62.750000 174.500000 ;
        RECT 62.550000 174.700000 62.750000 174.900000 ;
        RECT 62.550000 175.100000 62.750000 175.300000 ;
        RECT 62.550000 175.500000 62.750000 175.700000 ;
        RECT 62.550000 175.900000 62.750000 176.100000 ;
        RECT 62.550000 176.300000 62.750000 176.500000 ;
        RECT 62.550000 176.700000 62.750000 176.900000 ;
        RECT 62.550000 177.100000 62.750000 177.300000 ;
        RECT 62.550000 177.500000 62.750000 177.700000 ;
        RECT 62.550000 177.900000 62.750000 178.100000 ;
        RECT 62.550000 178.300000 62.750000 178.500000 ;
        RECT 62.550000 178.700000 62.750000 178.900000 ;
        RECT 62.550000 179.100000 62.750000 179.300000 ;
        RECT 62.550000 179.500000 62.750000 179.700000 ;
        RECT 62.550000 179.900000 62.750000 180.100000 ;
        RECT 62.550000 180.300000 62.750000 180.500000 ;
        RECT 62.550000 180.700000 62.750000 180.900000 ;
        RECT 62.550000 181.100000 62.750000 181.300000 ;
        RECT 62.550000 181.505000 62.750000 181.705000 ;
        RECT 62.550000 181.910000 62.750000 182.110000 ;
        RECT 62.550000 182.315000 62.750000 182.515000 ;
        RECT 62.550000 182.720000 62.750000 182.920000 ;
        RECT 62.550000 183.125000 62.750000 183.325000 ;
        RECT 62.550000 183.530000 62.750000 183.730000 ;
        RECT 62.550000 183.935000 62.750000 184.135000 ;
        RECT 62.550000 184.340000 62.750000 184.540000 ;
        RECT 62.550000 184.745000 62.750000 184.945000 ;
        RECT 62.550000 185.150000 62.750000 185.350000 ;
        RECT 62.550000 185.555000 62.750000 185.755000 ;
        RECT 62.550000 185.960000 62.750000 186.160000 ;
        RECT 62.550000 186.365000 62.750000 186.565000 ;
        RECT 62.550000 186.770000 62.750000 186.970000 ;
        RECT 62.550000 187.175000 62.750000 187.375000 ;
        RECT 62.550000 187.580000 62.750000 187.780000 ;
        RECT 62.550000 187.985000 62.750000 188.185000 ;
        RECT 62.550000 188.390000 62.750000 188.590000 ;
        RECT 62.550000 188.795000 62.750000 188.995000 ;
        RECT 62.550000 189.200000 62.750000 189.400000 ;
        RECT 62.550000 189.605000 62.750000 189.805000 ;
        RECT 62.550000 190.010000 62.750000 190.210000 ;
        RECT 62.550000 190.415000 62.750000 190.615000 ;
        RECT 62.550000 190.820000 62.750000 191.020000 ;
        RECT 62.550000 191.225000 62.750000 191.425000 ;
        RECT 62.550000 191.630000 62.750000 191.830000 ;
        RECT 62.550000 192.035000 62.750000 192.235000 ;
        RECT 62.550000 192.440000 62.750000 192.640000 ;
        RECT 62.550000 192.845000 62.750000 193.045000 ;
        RECT 62.550000 193.250000 62.750000 193.450000 ;
        RECT 62.550000 193.655000 62.750000 193.855000 ;
        RECT 62.550000 194.060000 62.750000 194.260000 ;
        RECT 62.550000 194.465000 62.750000 194.665000 ;
        RECT 62.550000 194.870000 62.750000 195.070000 ;
        RECT 62.550000 195.275000 62.750000 195.475000 ;
        RECT 62.550000 195.680000 62.750000 195.880000 ;
        RECT 62.550000 196.085000 62.750000 196.285000 ;
        RECT 62.550000 196.490000 62.750000 196.690000 ;
        RECT 62.550000 196.895000 62.750000 197.095000 ;
        RECT 62.550000 197.300000 62.750000 197.500000 ;
        RECT 62.550000 197.705000 62.750000 197.905000 ;
        RECT 62.660000  23.910000 62.860000  24.110000 ;
        RECT 62.660000  24.340000 62.860000  24.540000 ;
        RECT 62.660000  24.770000 62.860000  24.970000 ;
        RECT 62.660000  25.200000 62.860000  25.400000 ;
        RECT 62.660000  25.630000 62.860000  25.830000 ;
        RECT 62.660000  26.060000 62.860000  26.260000 ;
        RECT 62.660000  26.490000 62.860000  26.690000 ;
        RECT 62.660000  26.920000 62.860000  27.120000 ;
        RECT 62.660000  27.350000 62.860000  27.550000 ;
        RECT 62.660000  27.780000 62.860000  27.980000 ;
        RECT 62.660000  28.210000 62.860000  28.410000 ;
        RECT 62.960000 173.900000 63.160000 174.100000 ;
        RECT 62.960000 174.300000 63.160000 174.500000 ;
        RECT 62.960000 174.700000 63.160000 174.900000 ;
        RECT 62.960000 175.100000 63.160000 175.300000 ;
        RECT 62.960000 175.500000 63.160000 175.700000 ;
        RECT 62.960000 175.900000 63.160000 176.100000 ;
        RECT 62.960000 176.300000 63.160000 176.500000 ;
        RECT 62.960000 176.700000 63.160000 176.900000 ;
        RECT 62.960000 177.100000 63.160000 177.300000 ;
        RECT 62.960000 177.500000 63.160000 177.700000 ;
        RECT 62.960000 177.900000 63.160000 178.100000 ;
        RECT 62.960000 178.300000 63.160000 178.500000 ;
        RECT 62.960000 178.700000 63.160000 178.900000 ;
        RECT 62.960000 179.100000 63.160000 179.300000 ;
        RECT 62.960000 179.500000 63.160000 179.700000 ;
        RECT 62.960000 179.900000 63.160000 180.100000 ;
        RECT 62.960000 180.300000 63.160000 180.500000 ;
        RECT 62.960000 180.700000 63.160000 180.900000 ;
        RECT 62.960000 181.100000 63.160000 181.300000 ;
        RECT 62.960000 181.505000 63.160000 181.705000 ;
        RECT 62.960000 181.910000 63.160000 182.110000 ;
        RECT 62.960000 182.315000 63.160000 182.515000 ;
        RECT 62.960000 182.720000 63.160000 182.920000 ;
        RECT 62.960000 183.125000 63.160000 183.325000 ;
        RECT 62.960000 183.530000 63.160000 183.730000 ;
        RECT 62.960000 183.935000 63.160000 184.135000 ;
        RECT 62.960000 184.340000 63.160000 184.540000 ;
        RECT 62.960000 184.745000 63.160000 184.945000 ;
        RECT 62.960000 185.150000 63.160000 185.350000 ;
        RECT 62.960000 185.555000 63.160000 185.755000 ;
        RECT 62.960000 185.960000 63.160000 186.160000 ;
        RECT 62.960000 186.365000 63.160000 186.565000 ;
        RECT 62.960000 186.770000 63.160000 186.970000 ;
        RECT 62.960000 187.175000 63.160000 187.375000 ;
        RECT 62.960000 187.580000 63.160000 187.780000 ;
        RECT 62.960000 187.985000 63.160000 188.185000 ;
        RECT 62.960000 188.390000 63.160000 188.590000 ;
        RECT 62.960000 188.795000 63.160000 188.995000 ;
        RECT 62.960000 189.200000 63.160000 189.400000 ;
        RECT 62.960000 189.605000 63.160000 189.805000 ;
        RECT 62.960000 190.010000 63.160000 190.210000 ;
        RECT 62.960000 190.415000 63.160000 190.615000 ;
        RECT 62.960000 190.820000 63.160000 191.020000 ;
        RECT 62.960000 191.225000 63.160000 191.425000 ;
        RECT 62.960000 191.630000 63.160000 191.830000 ;
        RECT 62.960000 192.035000 63.160000 192.235000 ;
        RECT 62.960000 192.440000 63.160000 192.640000 ;
        RECT 62.960000 192.845000 63.160000 193.045000 ;
        RECT 62.960000 193.250000 63.160000 193.450000 ;
        RECT 62.960000 193.655000 63.160000 193.855000 ;
        RECT 62.960000 194.060000 63.160000 194.260000 ;
        RECT 62.960000 194.465000 63.160000 194.665000 ;
        RECT 62.960000 194.870000 63.160000 195.070000 ;
        RECT 62.960000 195.275000 63.160000 195.475000 ;
        RECT 62.960000 195.680000 63.160000 195.880000 ;
        RECT 62.960000 196.085000 63.160000 196.285000 ;
        RECT 62.960000 196.490000 63.160000 196.690000 ;
        RECT 62.960000 196.895000 63.160000 197.095000 ;
        RECT 62.960000 197.300000 63.160000 197.500000 ;
        RECT 62.960000 197.705000 63.160000 197.905000 ;
        RECT 63.065000  23.910000 63.265000  24.110000 ;
        RECT 63.065000  24.340000 63.265000  24.540000 ;
        RECT 63.065000  24.770000 63.265000  24.970000 ;
        RECT 63.065000  25.200000 63.265000  25.400000 ;
        RECT 63.065000  25.630000 63.265000  25.830000 ;
        RECT 63.065000  26.060000 63.265000  26.260000 ;
        RECT 63.065000  26.490000 63.265000  26.690000 ;
        RECT 63.065000  26.920000 63.265000  27.120000 ;
        RECT 63.065000  27.350000 63.265000  27.550000 ;
        RECT 63.065000  27.780000 63.265000  27.980000 ;
        RECT 63.065000  28.210000 63.265000  28.410000 ;
        RECT 63.370000 173.900000 63.570000 174.100000 ;
        RECT 63.370000 174.300000 63.570000 174.500000 ;
        RECT 63.370000 174.700000 63.570000 174.900000 ;
        RECT 63.370000 175.100000 63.570000 175.300000 ;
        RECT 63.370000 175.500000 63.570000 175.700000 ;
        RECT 63.370000 175.900000 63.570000 176.100000 ;
        RECT 63.370000 176.300000 63.570000 176.500000 ;
        RECT 63.370000 176.700000 63.570000 176.900000 ;
        RECT 63.370000 177.100000 63.570000 177.300000 ;
        RECT 63.370000 177.500000 63.570000 177.700000 ;
        RECT 63.370000 177.900000 63.570000 178.100000 ;
        RECT 63.370000 178.300000 63.570000 178.500000 ;
        RECT 63.370000 178.700000 63.570000 178.900000 ;
        RECT 63.370000 179.100000 63.570000 179.300000 ;
        RECT 63.370000 179.500000 63.570000 179.700000 ;
        RECT 63.370000 179.900000 63.570000 180.100000 ;
        RECT 63.370000 180.300000 63.570000 180.500000 ;
        RECT 63.370000 180.700000 63.570000 180.900000 ;
        RECT 63.370000 181.100000 63.570000 181.300000 ;
        RECT 63.370000 181.505000 63.570000 181.705000 ;
        RECT 63.370000 181.910000 63.570000 182.110000 ;
        RECT 63.370000 182.315000 63.570000 182.515000 ;
        RECT 63.370000 182.720000 63.570000 182.920000 ;
        RECT 63.370000 183.125000 63.570000 183.325000 ;
        RECT 63.370000 183.530000 63.570000 183.730000 ;
        RECT 63.370000 183.935000 63.570000 184.135000 ;
        RECT 63.370000 184.340000 63.570000 184.540000 ;
        RECT 63.370000 184.745000 63.570000 184.945000 ;
        RECT 63.370000 185.150000 63.570000 185.350000 ;
        RECT 63.370000 185.555000 63.570000 185.755000 ;
        RECT 63.370000 185.960000 63.570000 186.160000 ;
        RECT 63.370000 186.365000 63.570000 186.565000 ;
        RECT 63.370000 186.770000 63.570000 186.970000 ;
        RECT 63.370000 187.175000 63.570000 187.375000 ;
        RECT 63.370000 187.580000 63.570000 187.780000 ;
        RECT 63.370000 187.985000 63.570000 188.185000 ;
        RECT 63.370000 188.390000 63.570000 188.590000 ;
        RECT 63.370000 188.795000 63.570000 188.995000 ;
        RECT 63.370000 189.200000 63.570000 189.400000 ;
        RECT 63.370000 189.605000 63.570000 189.805000 ;
        RECT 63.370000 190.010000 63.570000 190.210000 ;
        RECT 63.370000 190.415000 63.570000 190.615000 ;
        RECT 63.370000 190.820000 63.570000 191.020000 ;
        RECT 63.370000 191.225000 63.570000 191.425000 ;
        RECT 63.370000 191.630000 63.570000 191.830000 ;
        RECT 63.370000 192.035000 63.570000 192.235000 ;
        RECT 63.370000 192.440000 63.570000 192.640000 ;
        RECT 63.370000 192.845000 63.570000 193.045000 ;
        RECT 63.370000 193.250000 63.570000 193.450000 ;
        RECT 63.370000 193.655000 63.570000 193.855000 ;
        RECT 63.370000 194.060000 63.570000 194.260000 ;
        RECT 63.370000 194.465000 63.570000 194.665000 ;
        RECT 63.370000 194.870000 63.570000 195.070000 ;
        RECT 63.370000 195.275000 63.570000 195.475000 ;
        RECT 63.370000 195.680000 63.570000 195.880000 ;
        RECT 63.370000 196.085000 63.570000 196.285000 ;
        RECT 63.370000 196.490000 63.570000 196.690000 ;
        RECT 63.370000 196.895000 63.570000 197.095000 ;
        RECT 63.370000 197.300000 63.570000 197.500000 ;
        RECT 63.370000 197.705000 63.570000 197.905000 ;
        RECT 63.470000  23.910000 63.670000  24.110000 ;
        RECT 63.470000  24.340000 63.670000  24.540000 ;
        RECT 63.470000  24.770000 63.670000  24.970000 ;
        RECT 63.470000  25.200000 63.670000  25.400000 ;
        RECT 63.470000  25.630000 63.670000  25.830000 ;
        RECT 63.470000  26.060000 63.670000  26.260000 ;
        RECT 63.470000  26.490000 63.670000  26.690000 ;
        RECT 63.470000  26.920000 63.670000  27.120000 ;
        RECT 63.470000  27.350000 63.670000  27.550000 ;
        RECT 63.470000  27.780000 63.670000  27.980000 ;
        RECT 63.470000  28.210000 63.670000  28.410000 ;
        RECT 63.780000 173.900000 63.980000 174.100000 ;
        RECT 63.780000 174.300000 63.980000 174.500000 ;
        RECT 63.780000 174.700000 63.980000 174.900000 ;
        RECT 63.780000 175.100000 63.980000 175.300000 ;
        RECT 63.780000 175.500000 63.980000 175.700000 ;
        RECT 63.780000 175.900000 63.980000 176.100000 ;
        RECT 63.780000 176.300000 63.980000 176.500000 ;
        RECT 63.780000 176.700000 63.980000 176.900000 ;
        RECT 63.780000 177.100000 63.980000 177.300000 ;
        RECT 63.780000 177.500000 63.980000 177.700000 ;
        RECT 63.780000 177.900000 63.980000 178.100000 ;
        RECT 63.780000 178.300000 63.980000 178.500000 ;
        RECT 63.780000 178.700000 63.980000 178.900000 ;
        RECT 63.780000 179.100000 63.980000 179.300000 ;
        RECT 63.780000 179.500000 63.980000 179.700000 ;
        RECT 63.780000 179.900000 63.980000 180.100000 ;
        RECT 63.780000 180.300000 63.980000 180.500000 ;
        RECT 63.780000 180.700000 63.980000 180.900000 ;
        RECT 63.780000 181.100000 63.980000 181.300000 ;
        RECT 63.780000 181.505000 63.980000 181.705000 ;
        RECT 63.780000 181.910000 63.980000 182.110000 ;
        RECT 63.780000 182.315000 63.980000 182.515000 ;
        RECT 63.780000 182.720000 63.980000 182.920000 ;
        RECT 63.780000 183.125000 63.980000 183.325000 ;
        RECT 63.780000 183.530000 63.980000 183.730000 ;
        RECT 63.780000 183.935000 63.980000 184.135000 ;
        RECT 63.780000 184.340000 63.980000 184.540000 ;
        RECT 63.780000 184.745000 63.980000 184.945000 ;
        RECT 63.780000 185.150000 63.980000 185.350000 ;
        RECT 63.780000 185.555000 63.980000 185.755000 ;
        RECT 63.780000 185.960000 63.980000 186.160000 ;
        RECT 63.780000 186.365000 63.980000 186.565000 ;
        RECT 63.780000 186.770000 63.980000 186.970000 ;
        RECT 63.780000 187.175000 63.980000 187.375000 ;
        RECT 63.780000 187.580000 63.980000 187.780000 ;
        RECT 63.780000 187.985000 63.980000 188.185000 ;
        RECT 63.780000 188.390000 63.980000 188.590000 ;
        RECT 63.780000 188.795000 63.980000 188.995000 ;
        RECT 63.780000 189.200000 63.980000 189.400000 ;
        RECT 63.780000 189.605000 63.980000 189.805000 ;
        RECT 63.780000 190.010000 63.980000 190.210000 ;
        RECT 63.780000 190.415000 63.980000 190.615000 ;
        RECT 63.780000 190.820000 63.980000 191.020000 ;
        RECT 63.780000 191.225000 63.980000 191.425000 ;
        RECT 63.780000 191.630000 63.980000 191.830000 ;
        RECT 63.780000 192.035000 63.980000 192.235000 ;
        RECT 63.780000 192.440000 63.980000 192.640000 ;
        RECT 63.780000 192.845000 63.980000 193.045000 ;
        RECT 63.780000 193.250000 63.980000 193.450000 ;
        RECT 63.780000 193.655000 63.980000 193.855000 ;
        RECT 63.780000 194.060000 63.980000 194.260000 ;
        RECT 63.780000 194.465000 63.980000 194.665000 ;
        RECT 63.780000 194.870000 63.980000 195.070000 ;
        RECT 63.780000 195.275000 63.980000 195.475000 ;
        RECT 63.780000 195.680000 63.980000 195.880000 ;
        RECT 63.780000 196.085000 63.980000 196.285000 ;
        RECT 63.780000 196.490000 63.980000 196.690000 ;
        RECT 63.780000 196.895000 63.980000 197.095000 ;
        RECT 63.780000 197.300000 63.980000 197.500000 ;
        RECT 63.780000 197.705000 63.980000 197.905000 ;
        RECT 63.875000  23.910000 64.075000  24.110000 ;
        RECT 63.875000  24.340000 64.075000  24.540000 ;
        RECT 63.875000  24.770000 64.075000  24.970000 ;
        RECT 63.875000  25.200000 64.075000  25.400000 ;
        RECT 63.875000  25.630000 64.075000  25.830000 ;
        RECT 63.875000  26.060000 64.075000  26.260000 ;
        RECT 63.875000  26.490000 64.075000  26.690000 ;
        RECT 63.875000  26.920000 64.075000  27.120000 ;
        RECT 63.875000  27.350000 64.075000  27.550000 ;
        RECT 63.875000  27.780000 64.075000  27.980000 ;
        RECT 63.875000  28.210000 64.075000  28.410000 ;
        RECT 64.190000 173.900000 64.390000 174.100000 ;
        RECT 64.190000 174.300000 64.390000 174.500000 ;
        RECT 64.190000 174.700000 64.390000 174.900000 ;
        RECT 64.190000 175.100000 64.390000 175.300000 ;
        RECT 64.190000 175.500000 64.390000 175.700000 ;
        RECT 64.190000 175.900000 64.390000 176.100000 ;
        RECT 64.190000 176.300000 64.390000 176.500000 ;
        RECT 64.190000 176.700000 64.390000 176.900000 ;
        RECT 64.190000 177.100000 64.390000 177.300000 ;
        RECT 64.190000 177.500000 64.390000 177.700000 ;
        RECT 64.190000 177.900000 64.390000 178.100000 ;
        RECT 64.190000 178.300000 64.390000 178.500000 ;
        RECT 64.190000 178.700000 64.390000 178.900000 ;
        RECT 64.190000 179.100000 64.390000 179.300000 ;
        RECT 64.190000 179.500000 64.390000 179.700000 ;
        RECT 64.190000 179.900000 64.390000 180.100000 ;
        RECT 64.190000 180.300000 64.390000 180.500000 ;
        RECT 64.190000 180.700000 64.390000 180.900000 ;
        RECT 64.190000 181.100000 64.390000 181.300000 ;
        RECT 64.190000 181.505000 64.390000 181.705000 ;
        RECT 64.190000 181.910000 64.390000 182.110000 ;
        RECT 64.190000 182.315000 64.390000 182.515000 ;
        RECT 64.190000 182.720000 64.390000 182.920000 ;
        RECT 64.190000 183.125000 64.390000 183.325000 ;
        RECT 64.190000 183.530000 64.390000 183.730000 ;
        RECT 64.190000 183.935000 64.390000 184.135000 ;
        RECT 64.190000 184.340000 64.390000 184.540000 ;
        RECT 64.190000 184.745000 64.390000 184.945000 ;
        RECT 64.190000 185.150000 64.390000 185.350000 ;
        RECT 64.190000 185.555000 64.390000 185.755000 ;
        RECT 64.190000 185.960000 64.390000 186.160000 ;
        RECT 64.190000 186.365000 64.390000 186.565000 ;
        RECT 64.190000 186.770000 64.390000 186.970000 ;
        RECT 64.190000 187.175000 64.390000 187.375000 ;
        RECT 64.190000 187.580000 64.390000 187.780000 ;
        RECT 64.190000 187.985000 64.390000 188.185000 ;
        RECT 64.190000 188.390000 64.390000 188.590000 ;
        RECT 64.190000 188.795000 64.390000 188.995000 ;
        RECT 64.190000 189.200000 64.390000 189.400000 ;
        RECT 64.190000 189.605000 64.390000 189.805000 ;
        RECT 64.190000 190.010000 64.390000 190.210000 ;
        RECT 64.190000 190.415000 64.390000 190.615000 ;
        RECT 64.190000 190.820000 64.390000 191.020000 ;
        RECT 64.190000 191.225000 64.390000 191.425000 ;
        RECT 64.190000 191.630000 64.390000 191.830000 ;
        RECT 64.190000 192.035000 64.390000 192.235000 ;
        RECT 64.190000 192.440000 64.390000 192.640000 ;
        RECT 64.190000 192.845000 64.390000 193.045000 ;
        RECT 64.190000 193.250000 64.390000 193.450000 ;
        RECT 64.190000 193.655000 64.390000 193.855000 ;
        RECT 64.190000 194.060000 64.390000 194.260000 ;
        RECT 64.190000 194.465000 64.390000 194.665000 ;
        RECT 64.190000 194.870000 64.390000 195.070000 ;
        RECT 64.190000 195.275000 64.390000 195.475000 ;
        RECT 64.190000 195.680000 64.390000 195.880000 ;
        RECT 64.190000 196.085000 64.390000 196.285000 ;
        RECT 64.190000 196.490000 64.390000 196.690000 ;
        RECT 64.190000 196.895000 64.390000 197.095000 ;
        RECT 64.190000 197.300000 64.390000 197.500000 ;
        RECT 64.190000 197.705000 64.390000 197.905000 ;
        RECT 64.280000  23.910000 64.480000  24.110000 ;
        RECT 64.280000  24.340000 64.480000  24.540000 ;
        RECT 64.280000  24.770000 64.480000  24.970000 ;
        RECT 64.280000  25.200000 64.480000  25.400000 ;
        RECT 64.280000  25.630000 64.480000  25.830000 ;
        RECT 64.280000  26.060000 64.480000  26.260000 ;
        RECT 64.280000  26.490000 64.480000  26.690000 ;
        RECT 64.280000  26.920000 64.480000  27.120000 ;
        RECT 64.280000  27.350000 64.480000  27.550000 ;
        RECT 64.280000  27.780000 64.480000  27.980000 ;
        RECT 64.280000  28.210000 64.480000  28.410000 ;
        RECT 64.600000 173.900000 64.800000 174.100000 ;
        RECT 64.600000 174.300000 64.800000 174.500000 ;
        RECT 64.600000 174.700000 64.800000 174.900000 ;
        RECT 64.600000 175.100000 64.800000 175.300000 ;
        RECT 64.600000 175.500000 64.800000 175.700000 ;
        RECT 64.600000 175.900000 64.800000 176.100000 ;
        RECT 64.600000 176.300000 64.800000 176.500000 ;
        RECT 64.600000 176.700000 64.800000 176.900000 ;
        RECT 64.600000 177.100000 64.800000 177.300000 ;
        RECT 64.600000 177.500000 64.800000 177.700000 ;
        RECT 64.600000 177.900000 64.800000 178.100000 ;
        RECT 64.600000 178.300000 64.800000 178.500000 ;
        RECT 64.600000 178.700000 64.800000 178.900000 ;
        RECT 64.600000 179.100000 64.800000 179.300000 ;
        RECT 64.600000 179.500000 64.800000 179.700000 ;
        RECT 64.600000 179.900000 64.800000 180.100000 ;
        RECT 64.600000 180.300000 64.800000 180.500000 ;
        RECT 64.600000 180.700000 64.800000 180.900000 ;
        RECT 64.600000 181.100000 64.800000 181.300000 ;
        RECT 64.600000 181.505000 64.800000 181.705000 ;
        RECT 64.600000 181.910000 64.800000 182.110000 ;
        RECT 64.600000 182.315000 64.800000 182.515000 ;
        RECT 64.600000 182.720000 64.800000 182.920000 ;
        RECT 64.600000 183.125000 64.800000 183.325000 ;
        RECT 64.600000 183.530000 64.800000 183.730000 ;
        RECT 64.600000 183.935000 64.800000 184.135000 ;
        RECT 64.600000 184.340000 64.800000 184.540000 ;
        RECT 64.600000 184.745000 64.800000 184.945000 ;
        RECT 64.600000 185.150000 64.800000 185.350000 ;
        RECT 64.600000 185.555000 64.800000 185.755000 ;
        RECT 64.600000 185.960000 64.800000 186.160000 ;
        RECT 64.600000 186.365000 64.800000 186.565000 ;
        RECT 64.600000 186.770000 64.800000 186.970000 ;
        RECT 64.600000 187.175000 64.800000 187.375000 ;
        RECT 64.600000 187.580000 64.800000 187.780000 ;
        RECT 64.600000 187.985000 64.800000 188.185000 ;
        RECT 64.600000 188.390000 64.800000 188.590000 ;
        RECT 64.600000 188.795000 64.800000 188.995000 ;
        RECT 64.600000 189.200000 64.800000 189.400000 ;
        RECT 64.600000 189.605000 64.800000 189.805000 ;
        RECT 64.600000 190.010000 64.800000 190.210000 ;
        RECT 64.600000 190.415000 64.800000 190.615000 ;
        RECT 64.600000 190.820000 64.800000 191.020000 ;
        RECT 64.600000 191.225000 64.800000 191.425000 ;
        RECT 64.600000 191.630000 64.800000 191.830000 ;
        RECT 64.600000 192.035000 64.800000 192.235000 ;
        RECT 64.600000 192.440000 64.800000 192.640000 ;
        RECT 64.600000 192.845000 64.800000 193.045000 ;
        RECT 64.600000 193.250000 64.800000 193.450000 ;
        RECT 64.600000 193.655000 64.800000 193.855000 ;
        RECT 64.600000 194.060000 64.800000 194.260000 ;
        RECT 64.600000 194.465000 64.800000 194.665000 ;
        RECT 64.600000 194.870000 64.800000 195.070000 ;
        RECT 64.600000 195.275000 64.800000 195.475000 ;
        RECT 64.600000 195.680000 64.800000 195.880000 ;
        RECT 64.600000 196.085000 64.800000 196.285000 ;
        RECT 64.600000 196.490000 64.800000 196.690000 ;
        RECT 64.600000 196.895000 64.800000 197.095000 ;
        RECT 64.600000 197.300000 64.800000 197.500000 ;
        RECT 64.600000 197.705000 64.800000 197.905000 ;
        RECT 64.685000  23.910000 64.885000  24.110000 ;
        RECT 64.685000  24.340000 64.885000  24.540000 ;
        RECT 64.685000  24.770000 64.885000  24.970000 ;
        RECT 64.685000  25.200000 64.885000  25.400000 ;
        RECT 64.685000  25.630000 64.885000  25.830000 ;
        RECT 64.685000  26.060000 64.885000  26.260000 ;
        RECT 64.685000  26.490000 64.885000  26.690000 ;
        RECT 64.685000  26.920000 64.885000  27.120000 ;
        RECT 64.685000  27.350000 64.885000  27.550000 ;
        RECT 64.685000  27.780000 64.885000  27.980000 ;
        RECT 64.685000  28.210000 64.885000  28.410000 ;
        RECT 65.010000 173.900000 65.210000 174.100000 ;
        RECT 65.010000 174.300000 65.210000 174.500000 ;
        RECT 65.010000 174.700000 65.210000 174.900000 ;
        RECT 65.010000 175.100000 65.210000 175.300000 ;
        RECT 65.010000 175.500000 65.210000 175.700000 ;
        RECT 65.010000 175.900000 65.210000 176.100000 ;
        RECT 65.010000 176.300000 65.210000 176.500000 ;
        RECT 65.010000 176.700000 65.210000 176.900000 ;
        RECT 65.010000 177.100000 65.210000 177.300000 ;
        RECT 65.010000 177.500000 65.210000 177.700000 ;
        RECT 65.010000 177.900000 65.210000 178.100000 ;
        RECT 65.010000 178.300000 65.210000 178.500000 ;
        RECT 65.010000 178.700000 65.210000 178.900000 ;
        RECT 65.010000 179.100000 65.210000 179.300000 ;
        RECT 65.010000 179.500000 65.210000 179.700000 ;
        RECT 65.010000 179.900000 65.210000 180.100000 ;
        RECT 65.010000 180.300000 65.210000 180.500000 ;
        RECT 65.010000 180.700000 65.210000 180.900000 ;
        RECT 65.010000 181.100000 65.210000 181.300000 ;
        RECT 65.010000 181.505000 65.210000 181.705000 ;
        RECT 65.010000 181.910000 65.210000 182.110000 ;
        RECT 65.010000 182.315000 65.210000 182.515000 ;
        RECT 65.010000 182.720000 65.210000 182.920000 ;
        RECT 65.010000 183.125000 65.210000 183.325000 ;
        RECT 65.010000 183.530000 65.210000 183.730000 ;
        RECT 65.010000 183.935000 65.210000 184.135000 ;
        RECT 65.010000 184.340000 65.210000 184.540000 ;
        RECT 65.010000 184.745000 65.210000 184.945000 ;
        RECT 65.010000 185.150000 65.210000 185.350000 ;
        RECT 65.010000 185.555000 65.210000 185.755000 ;
        RECT 65.010000 185.960000 65.210000 186.160000 ;
        RECT 65.010000 186.365000 65.210000 186.565000 ;
        RECT 65.010000 186.770000 65.210000 186.970000 ;
        RECT 65.010000 187.175000 65.210000 187.375000 ;
        RECT 65.010000 187.580000 65.210000 187.780000 ;
        RECT 65.010000 187.985000 65.210000 188.185000 ;
        RECT 65.010000 188.390000 65.210000 188.590000 ;
        RECT 65.010000 188.795000 65.210000 188.995000 ;
        RECT 65.010000 189.200000 65.210000 189.400000 ;
        RECT 65.010000 189.605000 65.210000 189.805000 ;
        RECT 65.010000 190.010000 65.210000 190.210000 ;
        RECT 65.010000 190.415000 65.210000 190.615000 ;
        RECT 65.010000 190.820000 65.210000 191.020000 ;
        RECT 65.010000 191.225000 65.210000 191.425000 ;
        RECT 65.010000 191.630000 65.210000 191.830000 ;
        RECT 65.010000 192.035000 65.210000 192.235000 ;
        RECT 65.010000 192.440000 65.210000 192.640000 ;
        RECT 65.010000 192.845000 65.210000 193.045000 ;
        RECT 65.010000 193.250000 65.210000 193.450000 ;
        RECT 65.010000 193.655000 65.210000 193.855000 ;
        RECT 65.010000 194.060000 65.210000 194.260000 ;
        RECT 65.010000 194.465000 65.210000 194.665000 ;
        RECT 65.010000 194.870000 65.210000 195.070000 ;
        RECT 65.010000 195.275000 65.210000 195.475000 ;
        RECT 65.010000 195.680000 65.210000 195.880000 ;
        RECT 65.010000 196.085000 65.210000 196.285000 ;
        RECT 65.010000 196.490000 65.210000 196.690000 ;
        RECT 65.010000 196.895000 65.210000 197.095000 ;
        RECT 65.010000 197.300000 65.210000 197.500000 ;
        RECT 65.010000 197.705000 65.210000 197.905000 ;
        RECT 65.090000  23.910000 65.290000  24.110000 ;
        RECT 65.090000  24.340000 65.290000  24.540000 ;
        RECT 65.090000  24.770000 65.290000  24.970000 ;
        RECT 65.090000  25.200000 65.290000  25.400000 ;
        RECT 65.090000  25.630000 65.290000  25.830000 ;
        RECT 65.090000  26.060000 65.290000  26.260000 ;
        RECT 65.090000  26.490000 65.290000  26.690000 ;
        RECT 65.090000  26.920000 65.290000  27.120000 ;
        RECT 65.090000  27.350000 65.290000  27.550000 ;
        RECT 65.090000  27.780000 65.290000  27.980000 ;
        RECT 65.090000  28.210000 65.290000  28.410000 ;
        RECT 65.420000 173.900000 65.620000 174.100000 ;
        RECT 65.420000 174.300000 65.620000 174.500000 ;
        RECT 65.420000 174.700000 65.620000 174.900000 ;
        RECT 65.420000 175.100000 65.620000 175.300000 ;
        RECT 65.420000 175.500000 65.620000 175.700000 ;
        RECT 65.420000 175.900000 65.620000 176.100000 ;
        RECT 65.420000 176.300000 65.620000 176.500000 ;
        RECT 65.420000 176.700000 65.620000 176.900000 ;
        RECT 65.420000 177.100000 65.620000 177.300000 ;
        RECT 65.420000 177.500000 65.620000 177.700000 ;
        RECT 65.420000 177.900000 65.620000 178.100000 ;
        RECT 65.420000 178.300000 65.620000 178.500000 ;
        RECT 65.420000 178.700000 65.620000 178.900000 ;
        RECT 65.420000 179.100000 65.620000 179.300000 ;
        RECT 65.420000 179.500000 65.620000 179.700000 ;
        RECT 65.420000 179.900000 65.620000 180.100000 ;
        RECT 65.420000 180.300000 65.620000 180.500000 ;
        RECT 65.420000 180.700000 65.620000 180.900000 ;
        RECT 65.420000 181.100000 65.620000 181.300000 ;
        RECT 65.420000 181.505000 65.620000 181.705000 ;
        RECT 65.420000 181.910000 65.620000 182.110000 ;
        RECT 65.420000 182.315000 65.620000 182.515000 ;
        RECT 65.420000 182.720000 65.620000 182.920000 ;
        RECT 65.420000 183.125000 65.620000 183.325000 ;
        RECT 65.420000 183.530000 65.620000 183.730000 ;
        RECT 65.420000 183.935000 65.620000 184.135000 ;
        RECT 65.420000 184.340000 65.620000 184.540000 ;
        RECT 65.420000 184.745000 65.620000 184.945000 ;
        RECT 65.420000 185.150000 65.620000 185.350000 ;
        RECT 65.420000 185.555000 65.620000 185.755000 ;
        RECT 65.420000 185.960000 65.620000 186.160000 ;
        RECT 65.420000 186.365000 65.620000 186.565000 ;
        RECT 65.420000 186.770000 65.620000 186.970000 ;
        RECT 65.420000 187.175000 65.620000 187.375000 ;
        RECT 65.420000 187.580000 65.620000 187.780000 ;
        RECT 65.420000 187.985000 65.620000 188.185000 ;
        RECT 65.420000 188.390000 65.620000 188.590000 ;
        RECT 65.420000 188.795000 65.620000 188.995000 ;
        RECT 65.420000 189.200000 65.620000 189.400000 ;
        RECT 65.420000 189.605000 65.620000 189.805000 ;
        RECT 65.420000 190.010000 65.620000 190.210000 ;
        RECT 65.420000 190.415000 65.620000 190.615000 ;
        RECT 65.420000 190.820000 65.620000 191.020000 ;
        RECT 65.420000 191.225000 65.620000 191.425000 ;
        RECT 65.420000 191.630000 65.620000 191.830000 ;
        RECT 65.420000 192.035000 65.620000 192.235000 ;
        RECT 65.420000 192.440000 65.620000 192.640000 ;
        RECT 65.420000 192.845000 65.620000 193.045000 ;
        RECT 65.420000 193.250000 65.620000 193.450000 ;
        RECT 65.420000 193.655000 65.620000 193.855000 ;
        RECT 65.420000 194.060000 65.620000 194.260000 ;
        RECT 65.420000 194.465000 65.620000 194.665000 ;
        RECT 65.420000 194.870000 65.620000 195.070000 ;
        RECT 65.420000 195.275000 65.620000 195.475000 ;
        RECT 65.420000 195.680000 65.620000 195.880000 ;
        RECT 65.420000 196.085000 65.620000 196.285000 ;
        RECT 65.420000 196.490000 65.620000 196.690000 ;
        RECT 65.420000 196.895000 65.620000 197.095000 ;
        RECT 65.420000 197.300000 65.620000 197.500000 ;
        RECT 65.420000 197.705000 65.620000 197.905000 ;
        RECT 65.495000  23.910000 65.695000  24.110000 ;
        RECT 65.495000  24.340000 65.695000  24.540000 ;
        RECT 65.495000  24.770000 65.695000  24.970000 ;
        RECT 65.495000  25.200000 65.695000  25.400000 ;
        RECT 65.495000  25.630000 65.695000  25.830000 ;
        RECT 65.495000  26.060000 65.695000  26.260000 ;
        RECT 65.495000  26.490000 65.695000  26.690000 ;
        RECT 65.495000  26.920000 65.695000  27.120000 ;
        RECT 65.495000  27.350000 65.695000  27.550000 ;
        RECT 65.495000  27.780000 65.695000  27.980000 ;
        RECT 65.495000  28.210000 65.695000  28.410000 ;
        RECT 65.830000 173.900000 66.030000 174.100000 ;
        RECT 65.830000 174.300000 66.030000 174.500000 ;
        RECT 65.830000 174.700000 66.030000 174.900000 ;
        RECT 65.830000 175.100000 66.030000 175.300000 ;
        RECT 65.830000 175.500000 66.030000 175.700000 ;
        RECT 65.830000 175.900000 66.030000 176.100000 ;
        RECT 65.830000 176.300000 66.030000 176.500000 ;
        RECT 65.830000 176.700000 66.030000 176.900000 ;
        RECT 65.830000 177.100000 66.030000 177.300000 ;
        RECT 65.830000 177.500000 66.030000 177.700000 ;
        RECT 65.830000 177.900000 66.030000 178.100000 ;
        RECT 65.830000 178.300000 66.030000 178.500000 ;
        RECT 65.830000 178.700000 66.030000 178.900000 ;
        RECT 65.830000 179.100000 66.030000 179.300000 ;
        RECT 65.830000 179.500000 66.030000 179.700000 ;
        RECT 65.830000 179.900000 66.030000 180.100000 ;
        RECT 65.830000 180.300000 66.030000 180.500000 ;
        RECT 65.830000 180.700000 66.030000 180.900000 ;
        RECT 65.830000 181.100000 66.030000 181.300000 ;
        RECT 65.830000 181.505000 66.030000 181.705000 ;
        RECT 65.830000 181.910000 66.030000 182.110000 ;
        RECT 65.830000 182.315000 66.030000 182.515000 ;
        RECT 65.830000 182.720000 66.030000 182.920000 ;
        RECT 65.830000 183.125000 66.030000 183.325000 ;
        RECT 65.830000 183.530000 66.030000 183.730000 ;
        RECT 65.830000 183.935000 66.030000 184.135000 ;
        RECT 65.830000 184.340000 66.030000 184.540000 ;
        RECT 65.830000 184.745000 66.030000 184.945000 ;
        RECT 65.830000 185.150000 66.030000 185.350000 ;
        RECT 65.830000 185.555000 66.030000 185.755000 ;
        RECT 65.830000 185.960000 66.030000 186.160000 ;
        RECT 65.830000 186.365000 66.030000 186.565000 ;
        RECT 65.830000 186.770000 66.030000 186.970000 ;
        RECT 65.830000 187.175000 66.030000 187.375000 ;
        RECT 65.830000 187.580000 66.030000 187.780000 ;
        RECT 65.830000 187.985000 66.030000 188.185000 ;
        RECT 65.830000 188.390000 66.030000 188.590000 ;
        RECT 65.830000 188.795000 66.030000 188.995000 ;
        RECT 65.830000 189.200000 66.030000 189.400000 ;
        RECT 65.830000 189.605000 66.030000 189.805000 ;
        RECT 65.830000 190.010000 66.030000 190.210000 ;
        RECT 65.830000 190.415000 66.030000 190.615000 ;
        RECT 65.830000 190.820000 66.030000 191.020000 ;
        RECT 65.830000 191.225000 66.030000 191.425000 ;
        RECT 65.830000 191.630000 66.030000 191.830000 ;
        RECT 65.830000 192.035000 66.030000 192.235000 ;
        RECT 65.830000 192.440000 66.030000 192.640000 ;
        RECT 65.830000 192.845000 66.030000 193.045000 ;
        RECT 65.830000 193.250000 66.030000 193.450000 ;
        RECT 65.830000 193.655000 66.030000 193.855000 ;
        RECT 65.830000 194.060000 66.030000 194.260000 ;
        RECT 65.830000 194.465000 66.030000 194.665000 ;
        RECT 65.830000 194.870000 66.030000 195.070000 ;
        RECT 65.830000 195.275000 66.030000 195.475000 ;
        RECT 65.830000 195.680000 66.030000 195.880000 ;
        RECT 65.830000 196.085000 66.030000 196.285000 ;
        RECT 65.830000 196.490000 66.030000 196.690000 ;
        RECT 65.830000 196.895000 66.030000 197.095000 ;
        RECT 65.830000 197.300000 66.030000 197.500000 ;
        RECT 65.830000 197.705000 66.030000 197.905000 ;
        RECT 65.900000  23.910000 66.100000  24.110000 ;
        RECT 65.900000  24.340000 66.100000  24.540000 ;
        RECT 65.900000  24.770000 66.100000  24.970000 ;
        RECT 65.900000  25.200000 66.100000  25.400000 ;
        RECT 65.900000  25.630000 66.100000  25.830000 ;
        RECT 65.900000  26.060000 66.100000  26.260000 ;
        RECT 65.900000  26.490000 66.100000  26.690000 ;
        RECT 65.900000  26.920000 66.100000  27.120000 ;
        RECT 65.900000  27.350000 66.100000  27.550000 ;
        RECT 65.900000  27.780000 66.100000  27.980000 ;
        RECT 65.900000  28.210000 66.100000  28.410000 ;
        RECT 66.240000 173.900000 66.440000 174.100000 ;
        RECT 66.240000 174.300000 66.440000 174.500000 ;
        RECT 66.240000 174.700000 66.440000 174.900000 ;
        RECT 66.240000 175.100000 66.440000 175.300000 ;
        RECT 66.240000 175.500000 66.440000 175.700000 ;
        RECT 66.240000 175.900000 66.440000 176.100000 ;
        RECT 66.240000 176.300000 66.440000 176.500000 ;
        RECT 66.240000 176.700000 66.440000 176.900000 ;
        RECT 66.240000 177.100000 66.440000 177.300000 ;
        RECT 66.240000 177.500000 66.440000 177.700000 ;
        RECT 66.240000 177.900000 66.440000 178.100000 ;
        RECT 66.240000 178.300000 66.440000 178.500000 ;
        RECT 66.240000 178.700000 66.440000 178.900000 ;
        RECT 66.240000 179.100000 66.440000 179.300000 ;
        RECT 66.240000 179.500000 66.440000 179.700000 ;
        RECT 66.240000 179.900000 66.440000 180.100000 ;
        RECT 66.240000 180.300000 66.440000 180.500000 ;
        RECT 66.240000 180.700000 66.440000 180.900000 ;
        RECT 66.240000 181.100000 66.440000 181.300000 ;
        RECT 66.240000 181.505000 66.440000 181.705000 ;
        RECT 66.240000 181.910000 66.440000 182.110000 ;
        RECT 66.240000 182.315000 66.440000 182.515000 ;
        RECT 66.240000 182.720000 66.440000 182.920000 ;
        RECT 66.240000 183.125000 66.440000 183.325000 ;
        RECT 66.240000 183.530000 66.440000 183.730000 ;
        RECT 66.240000 183.935000 66.440000 184.135000 ;
        RECT 66.240000 184.340000 66.440000 184.540000 ;
        RECT 66.240000 184.745000 66.440000 184.945000 ;
        RECT 66.240000 185.150000 66.440000 185.350000 ;
        RECT 66.240000 185.555000 66.440000 185.755000 ;
        RECT 66.240000 185.960000 66.440000 186.160000 ;
        RECT 66.240000 186.365000 66.440000 186.565000 ;
        RECT 66.240000 186.770000 66.440000 186.970000 ;
        RECT 66.240000 187.175000 66.440000 187.375000 ;
        RECT 66.240000 187.580000 66.440000 187.780000 ;
        RECT 66.240000 187.985000 66.440000 188.185000 ;
        RECT 66.240000 188.390000 66.440000 188.590000 ;
        RECT 66.240000 188.795000 66.440000 188.995000 ;
        RECT 66.240000 189.200000 66.440000 189.400000 ;
        RECT 66.240000 189.605000 66.440000 189.805000 ;
        RECT 66.240000 190.010000 66.440000 190.210000 ;
        RECT 66.240000 190.415000 66.440000 190.615000 ;
        RECT 66.240000 190.820000 66.440000 191.020000 ;
        RECT 66.240000 191.225000 66.440000 191.425000 ;
        RECT 66.240000 191.630000 66.440000 191.830000 ;
        RECT 66.240000 192.035000 66.440000 192.235000 ;
        RECT 66.240000 192.440000 66.440000 192.640000 ;
        RECT 66.240000 192.845000 66.440000 193.045000 ;
        RECT 66.240000 193.250000 66.440000 193.450000 ;
        RECT 66.240000 193.655000 66.440000 193.855000 ;
        RECT 66.240000 194.060000 66.440000 194.260000 ;
        RECT 66.240000 194.465000 66.440000 194.665000 ;
        RECT 66.240000 194.870000 66.440000 195.070000 ;
        RECT 66.240000 195.275000 66.440000 195.475000 ;
        RECT 66.240000 195.680000 66.440000 195.880000 ;
        RECT 66.240000 196.085000 66.440000 196.285000 ;
        RECT 66.240000 196.490000 66.440000 196.690000 ;
        RECT 66.240000 196.895000 66.440000 197.095000 ;
        RECT 66.240000 197.300000 66.440000 197.500000 ;
        RECT 66.240000 197.705000 66.440000 197.905000 ;
        RECT 66.305000  23.910000 66.505000  24.110000 ;
        RECT 66.305000  24.340000 66.505000  24.540000 ;
        RECT 66.305000  24.770000 66.505000  24.970000 ;
        RECT 66.305000  25.200000 66.505000  25.400000 ;
        RECT 66.305000  25.630000 66.505000  25.830000 ;
        RECT 66.305000  26.060000 66.505000  26.260000 ;
        RECT 66.305000  26.490000 66.505000  26.690000 ;
        RECT 66.305000  26.920000 66.505000  27.120000 ;
        RECT 66.305000  27.350000 66.505000  27.550000 ;
        RECT 66.305000  27.780000 66.505000  27.980000 ;
        RECT 66.305000  28.210000 66.505000  28.410000 ;
        RECT 66.650000 173.900000 66.850000 174.100000 ;
        RECT 66.650000 174.300000 66.850000 174.500000 ;
        RECT 66.650000 174.700000 66.850000 174.900000 ;
        RECT 66.650000 175.100000 66.850000 175.300000 ;
        RECT 66.650000 175.500000 66.850000 175.700000 ;
        RECT 66.650000 175.900000 66.850000 176.100000 ;
        RECT 66.650000 176.300000 66.850000 176.500000 ;
        RECT 66.650000 176.700000 66.850000 176.900000 ;
        RECT 66.650000 177.100000 66.850000 177.300000 ;
        RECT 66.650000 177.500000 66.850000 177.700000 ;
        RECT 66.650000 177.900000 66.850000 178.100000 ;
        RECT 66.650000 178.300000 66.850000 178.500000 ;
        RECT 66.650000 178.700000 66.850000 178.900000 ;
        RECT 66.650000 179.100000 66.850000 179.300000 ;
        RECT 66.650000 179.500000 66.850000 179.700000 ;
        RECT 66.650000 179.900000 66.850000 180.100000 ;
        RECT 66.650000 180.300000 66.850000 180.500000 ;
        RECT 66.650000 180.700000 66.850000 180.900000 ;
        RECT 66.650000 181.100000 66.850000 181.300000 ;
        RECT 66.650000 181.505000 66.850000 181.705000 ;
        RECT 66.650000 181.910000 66.850000 182.110000 ;
        RECT 66.650000 182.315000 66.850000 182.515000 ;
        RECT 66.650000 182.720000 66.850000 182.920000 ;
        RECT 66.650000 183.125000 66.850000 183.325000 ;
        RECT 66.650000 183.530000 66.850000 183.730000 ;
        RECT 66.650000 183.935000 66.850000 184.135000 ;
        RECT 66.650000 184.340000 66.850000 184.540000 ;
        RECT 66.650000 184.745000 66.850000 184.945000 ;
        RECT 66.650000 185.150000 66.850000 185.350000 ;
        RECT 66.650000 185.555000 66.850000 185.755000 ;
        RECT 66.650000 185.960000 66.850000 186.160000 ;
        RECT 66.650000 186.365000 66.850000 186.565000 ;
        RECT 66.650000 186.770000 66.850000 186.970000 ;
        RECT 66.650000 187.175000 66.850000 187.375000 ;
        RECT 66.650000 187.580000 66.850000 187.780000 ;
        RECT 66.650000 187.985000 66.850000 188.185000 ;
        RECT 66.650000 188.390000 66.850000 188.590000 ;
        RECT 66.650000 188.795000 66.850000 188.995000 ;
        RECT 66.650000 189.200000 66.850000 189.400000 ;
        RECT 66.650000 189.605000 66.850000 189.805000 ;
        RECT 66.650000 190.010000 66.850000 190.210000 ;
        RECT 66.650000 190.415000 66.850000 190.615000 ;
        RECT 66.650000 190.820000 66.850000 191.020000 ;
        RECT 66.650000 191.225000 66.850000 191.425000 ;
        RECT 66.650000 191.630000 66.850000 191.830000 ;
        RECT 66.650000 192.035000 66.850000 192.235000 ;
        RECT 66.650000 192.440000 66.850000 192.640000 ;
        RECT 66.650000 192.845000 66.850000 193.045000 ;
        RECT 66.650000 193.250000 66.850000 193.450000 ;
        RECT 66.650000 193.655000 66.850000 193.855000 ;
        RECT 66.650000 194.060000 66.850000 194.260000 ;
        RECT 66.650000 194.465000 66.850000 194.665000 ;
        RECT 66.650000 194.870000 66.850000 195.070000 ;
        RECT 66.650000 195.275000 66.850000 195.475000 ;
        RECT 66.650000 195.680000 66.850000 195.880000 ;
        RECT 66.650000 196.085000 66.850000 196.285000 ;
        RECT 66.650000 196.490000 66.850000 196.690000 ;
        RECT 66.650000 196.895000 66.850000 197.095000 ;
        RECT 66.650000 197.300000 66.850000 197.500000 ;
        RECT 66.650000 197.705000 66.850000 197.905000 ;
        RECT 66.710000  23.910000 66.910000  24.110000 ;
        RECT 66.710000  24.340000 66.910000  24.540000 ;
        RECT 66.710000  24.770000 66.910000  24.970000 ;
        RECT 66.710000  25.200000 66.910000  25.400000 ;
        RECT 66.710000  25.630000 66.910000  25.830000 ;
        RECT 66.710000  26.060000 66.910000  26.260000 ;
        RECT 66.710000  26.490000 66.910000  26.690000 ;
        RECT 66.710000  26.920000 66.910000  27.120000 ;
        RECT 66.710000  27.350000 66.910000  27.550000 ;
        RECT 66.710000  27.780000 66.910000  27.980000 ;
        RECT 66.710000  28.210000 66.910000  28.410000 ;
        RECT 67.060000 173.900000 67.260000 174.100000 ;
        RECT 67.060000 174.300000 67.260000 174.500000 ;
        RECT 67.060000 174.700000 67.260000 174.900000 ;
        RECT 67.060000 175.100000 67.260000 175.300000 ;
        RECT 67.060000 175.500000 67.260000 175.700000 ;
        RECT 67.060000 175.900000 67.260000 176.100000 ;
        RECT 67.060000 176.300000 67.260000 176.500000 ;
        RECT 67.060000 176.700000 67.260000 176.900000 ;
        RECT 67.060000 177.100000 67.260000 177.300000 ;
        RECT 67.060000 177.500000 67.260000 177.700000 ;
        RECT 67.060000 177.900000 67.260000 178.100000 ;
        RECT 67.060000 178.300000 67.260000 178.500000 ;
        RECT 67.060000 178.700000 67.260000 178.900000 ;
        RECT 67.060000 179.100000 67.260000 179.300000 ;
        RECT 67.060000 179.500000 67.260000 179.700000 ;
        RECT 67.060000 179.900000 67.260000 180.100000 ;
        RECT 67.060000 180.300000 67.260000 180.500000 ;
        RECT 67.060000 180.700000 67.260000 180.900000 ;
        RECT 67.060000 181.100000 67.260000 181.300000 ;
        RECT 67.060000 181.505000 67.260000 181.705000 ;
        RECT 67.060000 181.910000 67.260000 182.110000 ;
        RECT 67.060000 182.315000 67.260000 182.515000 ;
        RECT 67.060000 182.720000 67.260000 182.920000 ;
        RECT 67.060000 183.125000 67.260000 183.325000 ;
        RECT 67.060000 183.530000 67.260000 183.730000 ;
        RECT 67.060000 183.935000 67.260000 184.135000 ;
        RECT 67.060000 184.340000 67.260000 184.540000 ;
        RECT 67.060000 184.745000 67.260000 184.945000 ;
        RECT 67.060000 185.150000 67.260000 185.350000 ;
        RECT 67.060000 185.555000 67.260000 185.755000 ;
        RECT 67.060000 185.960000 67.260000 186.160000 ;
        RECT 67.060000 186.365000 67.260000 186.565000 ;
        RECT 67.060000 186.770000 67.260000 186.970000 ;
        RECT 67.060000 187.175000 67.260000 187.375000 ;
        RECT 67.060000 187.580000 67.260000 187.780000 ;
        RECT 67.060000 187.985000 67.260000 188.185000 ;
        RECT 67.060000 188.390000 67.260000 188.590000 ;
        RECT 67.060000 188.795000 67.260000 188.995000 ;
        RECT 67.060000 189.200000 67.260000 189.400000 ;
        RECT 67.060000 189.605000 67.260000 189.805000 ;
        RECT 67.060000 190.010000 67.260000 190.210000 ;
        RECT 67.060000 190.415000 67.260000 190.615000 ;
        RECT 67.060000 190.820000 67.260000 191.020000 ;
        RECT 67.060000 191.225000 67.260000 191.425000 ;
        RECT 67.060000 191.630000 67.260000 191.830000 ;
        RECT 67.060000 192.035000 67.260000 192.235000 ;
        RECT 67.060000 192.440000 67.260000 192.640000 ;
        RECT 67.060000 192.845000 67.260000 193.045000 ;
        RECT 67.060000 193.250000 67.260000 193.450000 ;
        RECT 67.060000 193.655000 67.260000 193.855000 ;
        RECT 67.060000 194.060000 67.260000 194.260000 ;
        RECT 67.060000 194.465000 67.260000 194.665000 ;
        RECT 67.060000 194.870000 67.260000 195.070000 ;
        RECT 67.060000 195.275000 67.260000 195.475000 ;
        RECT 67.060000 195.680000 67.260000 195.880000 ;
        RECT 67.060000 196.085000 67.260000 196.285000 ;
        RECT 67.060000 196.490000 67.260000 196.690000 ;
        RECT 67.060000 196.895000 67.260000 197.095000 ;
        RECT 67.060000 197.300000 67.260000 197.500000 ;
        RECT 67.060000 197.705000 67.260000 197.905000 ;
        RECT 67.115000  23.910000 67.315000  24.110000 ;
        RECT 67.115000  24.340000 67.315000  24.540000 ;
        RECT 67.115000  24.770000 67.315000  24.970000 ;
        RECT 67.115000  25.200000 67.315000  25.400000 ;
        RECT 67.115000  25.630000 67.315000  25.830000 ;
        RECT 67.115000  26.060000 67.315000  26.260000 ;
        RECT 67.115000  26.490000 67.315000  26.690000 ;
        RECT 67.115000  26.920000 67.315000  27.120000 ;
        RECT 67.115000  27.350000 67.315000  27.550000 ;
        RECT 67.115000  27.780000 67.315000  27.980000 ;
        RECT 67.115000  28.210000 67.315000  28.410000 ;
        RECT 67.470000 173.900000 67.670000 174.100000 ;
        RECT 67.470000 174.300000 67.670000 174.500000 ;
        RECT 67.470000 174.700000 67.670000 174.900000 ;
        RECT 67.470000 175.100000 67.670000 175.300000 ;
        RECT 67.470000 175.500000 67.670000 175.700000 ;
        RECT 67.470000 175.900000 67.670000 176.100000 ;
        RECT 67.470000 176.300000 67.670000 176.500000 ;
        RECT 67.470000 176.700000 67.670000 176.900000 ;
        RECT 67.470000 177.100000 67.670000 177.300000 ;
        RECT 67.470000 177.500000 67.670000 177.700000 ;
        RECT 67.470000 177.900000 67.670000 178.100000 ;
        RECT 67.470000 178.300000 67.670000 178.500000 ;
        RECT 67.470000 178.700000 67.670000 178.900000 ;
        RECT 67.470000 179.100000 67.670000 179.300000 ;
        RECT 67.470000 179.500000 67.670000 179.700000 ;
        RECT 67.470000 179.900000 67.670000 180.100000 ;
        RECT 67.470000 180.300000 67.670000 180.500000 ;
        RECT 67.470000 180.700000 67.670000 180.900000 ;
        RECT 67.470000 181.100000 67.670000 181.300000 ;
        RECT 67.470000 181.505000 67.670000 181.705000 ;
        RECT 67.470000 181.910000 67.670000 182.110000 ;
        RECT 67.470000 182.315000 67.670000 182.515000 ;
        RECT 67.470000 182.720000 67.670000 182.920000 ;
        RECT 67.470000 183.125000 67.670000 183.325000 ;
        RECT 67.470000 183.530000 67.670000 183.730000 ;
        RECT 67.470000 183.935000 67.670000 184.135000 ;
        RECT 67.470000 184.340000 67.670000 184.540000 ;
        RECT 67.470000 184.745000 67.670000 184.945000 ;
        RECT 67.470000 185.150000 67.670000 185.350000 ;
        RECT 67.470000 185.555000 67.670000 185.755000 ;
        RECT 67.470000 185.960000 67.670000 186.160000 ;
        RECT 67.470000 186.365000 67.670000 186.565000 ;
        RECT 67.470000 186.770000 67.670000 186.970000 ;
        RECT 67.470000 187.175000 67.670000 187.375000 ;
        RECT 67.470000 187.580000 67.670000 187.780000 ;
        RECT 67.470000 187.985000 67.670000 188.185000 ;
        RECT 67.470000 188.390000 67.670000 188.590000 ;
        RECT 67.470000 188.795000 67.670000 188.995000 ;
        RECT 67.470000 189.200000 67.670000 189.400000 ;
        RECT 67.470000 189.605000 67.670000 189.805000 ;
        RECT 67.470000 190.010000 67.670000 190.210000 ;
        RECT 67.470000 190.415000 67.670000 190.615000 ;
        RECT 67.470000 190.820000 67.670000 191.020000 ;
        RECT 67.470000 191.225000 67.670000 191.425000 ;
        RECT 67.470000 191.630000 67.670000 191.830000 ;
        RECT 67.470000 192.035000 67.670000 192.235000 ;
        RECT 67.470000 192.440000 67.670000 192.640000 ;
        RECT 67.470000 192.845000 67.670000 193.045000 ;
        RECT 67.470000 193.250000 67.670000 193.450000 ;
        RECT 67.470000 193.655000 67.670000 193.855000 ;
        RECT 67.470000 194.060000 67.670000 194.260000 ;
        RECT 67.470000 194.465000 67.670000 194.665000 ;
        RECT 67.470000 194.870000 67.670000 195.070000 ;
        RECT 67.470000 195.275000 67.670000 195.475000 ;
        RECT 67.470000 195.680000 67.670000 195.880000 ;
        RECT 67.470000 196.085000 67.670000 196.285000 ;
        RECT 67.470000 196.490000 67.670000 196.690000 ;
        RECT 67.470000 196.895000 67.670000 197.095000 ;
        RECT 67.470000 197.300000 67.670000 197.500000 ;
        RECT 67.470000 197.705000 67.670000 197.905000 ;
        RECT 67.520000  23.910000 67.720000  24.110000 ;
        RECT 67.520000  24.340000 67.720000  24.540000 ;
        RECT 67.520000  24.770000 67.720000  24.970000 ;
        RECT 67.520000  25.200000 67.720000  25.400000 ;
        RECT 67.520000  25.630000 67.720000  25.830000 ;
        RECT 67.520000  26.060000 67.720000  26.260000 ;
        RECT 67.520000  26.490000 67.720000  26.690000 ;
        RECT 67.520000  26.920000 67.720000  27.120000 ;
        RECT 67.520000  27.350000 67.720000  27.550000 ;
        RECT 67.520000  27.780000 67.720000  27.980000 ;
        RECT 67.520000  28.210000 67.720000  28.410000 ;
        RECT 67.880000 173.900000 68.080000 174.100000 ;
        RECT 67.880000 174.300000 68.080000 174.500000 ;
        RECT 67.880000 174.700000 68.080000 174.900000 ;
        RECT 67.880000 175.100000 68.080000 175.300000 ;
        RECT 67.880000 175.500000 68.080000 175.700000 ;
        RECT 67.880000 175.900000 68.080000 176.100000 ;
        RECT 67.880000 176.300000 68.080000 176.500000 ;
        RECT 67.880000 176.700000 68.080000 176.900000 ;
        RECT 67.880000 177.100000 68.080000 177.300000 ;
        RECT 67.880000 177.500000 68.080000 177.700000 ;
        RECT 67.880000 177.900000 68.080000 178.100000 ;
        RECT 67.880000 178.300000 68.080000 178.500000 ;
        RECT 67.880000 178.700000 68.080000 178.900000 ;
        RECT 67.880000 179.100000 68.080000 179.300000 ;
        RECT 67.880000 179.500000 68.080000 179.700000 ;
        RECT 67.880000 179.900000 68.080000 180.100000 ;
        RECT 67.880000 180.300000 68.080000 180.500000 ;
        RECT 67.880000 180.700000 68.080000 180.900000 ;
        RECT 67.880000 181.100000 68.080000 181.300000 ;
        RECT 67.880000 181.505000 68.080000 181.705000 ;
        RECT 67.880000 181.910000 68.080000 182.110000 ;
        RECT 67.880000 182.315000 68.080000 182.515000 ;
        RECT 67.880000 182.720000 68.080000 182.920000 ;
        RECT 67.880000 183.125000 68.080000 183.325000 ;
        RECT 67.880000 183.530000 68.080000 183.730000 ;
        RECT 67.880000 183.935000 68.080000 184.135000 ;
        RECT 67.880000 184.340000 68.080000 184.540000 ;
        RECT 67.880000 184.745000 68.080000 184.945000 ;
        RECT 67.880000 185.150000 68.080000 185.350000 ;
        RECT 67.880000 185.555000 68.080000 185.755000 ;
        RECT 67.880000 185.960000 68.080000 186.160000 ;
        RECT 67.880000 186.365000 68.080000 186.565000 ;
        RECT 67.880000 186.770000 68.080000 186.970000 ;
        RECT 67.880000 187.175000 68.080000 187.375000 ;
        RECT 67.880000 187.580000 68.080000 187.780000 ;
        RECT 67.880000 187.985000 68.080000 188.185000 ;
        RECT 67.880000 188.390000 68.080000 188.590000 ;
        RECT 67.880000 188.795000 68.080000 188.995000 ;
        RECT 67.880000 189.200000 68.080000 189.400000 ;
        RECT 67.880000 189.605000 68.080000 189.805000 ;
        RECT 67.880000 190.010000 68.080000 190.210000 ;
        RECT 67.880000 190.415000 68.080000 190.615000 ;
        RECT 67.880000 190.820000 68.080000 191.020000 ;
        RECT 67.880000 191.225000 68.080000 191.425000 ;
        RECT 67.880000 191.630000 68.080000 191.830000 ;
        RECT 67.880000 192.035000 68.080000 192.235000 ;
        RECT 67.880000 192.440000 68.080000 192.640000 ;
        RECT 67.880000 192.845000 68.080000 193.045000 ;
        RECT 67.880000 193.250000 68.080000 193.450000 ;
        RECT 67.880000 193.655000 68.080000 193.855000 ;
        RECT 67.880000 194.060000 68.080000 194.260000 ;
        RECT 67.880000 194.465000 68.080000 194.665000 ;
        RECT 67.880000 194.870000 68.080000 195.070000 ;
        RECT 67.880000 195.275000 68.080000 195.475000 ;
        RECT 67.880000 195.680000 68.080000 195.880000 ;
        RECT 67.880000 196.085000 68.080000 196.285000 ;
        RECT 67.880000 196.490000 68.080000 196.690000 ;
        RECT 67.880000 196.895000 68.080000 197.095000 ;
        RECT 67.880000 197.300000 68.080000 197.500000 ;
        RECT 67.880000 197.705000 68.080000 197.905000 ;
        RECT 67.925000  23.910000 68.125000  24.110000 ;
        RECT 67.925000  24.340000 68.125000  24.540000 ;
        RECT 67.925000  24.770000 68.125000  24.970000 ;
        RECT 67.925000  25.200000 68.125000  25.400000 ;
        RECT 67.925000  25.630000 68.125000  25.830000 ;
        RECT 67.925000  26.060000 68.125000  26.260000 ;
        RECT 67.925000  26.490000 68.125000  26.690000 ;
        RECT 67.925000  26.920000 68.125000  27.120000 ;
        RECT 67.925000  27.350000 68.125000  27.550000 ;
        RECT 67.925000  27.780000 68.125000  27.980000 ;
        RECT 67.925000  28.210000 68.125000  28.410000 ;
        RECT 68.290000 173.900000 68.490000 174.100000 ;
        RECT 68.290000 174.300000 68.490000 174.500000 ;
        RECT 68.290000 174.700000 68.490000 174.900000 ;
        RECT 68.290000 175.100000 68.490000 175.300000 ;
        RECT 68.290000 175.500000 68.490000 175.700000 ;
        RECT 68.290000 175.900000 68.490000 176.100000 ;
        RECT 68.290000 176.300000 68.490000 176.500000 ;
        RECT 68.290000 176.700000 68.490000 176.900000 ;
        RECT 68.290000 177.100000 68.490000 177.300000 ;
        RECT 68.290000 177.500000 68.490000 177.700000 ;
        RECT 68.290000 177.900000 68.490000 178.100000 ;
        RECT 68.290000 178.300000 68.490000 178.500000 ;
        RECT 68.290000 178.700000 68.490000 178.900000 ;
        RECT 68.290000 179.100000 68.490000 179.300000 ;
        RECT 68.290000 179.500000 68.490000 179.700000 ;
        RECT 68.290000 179.900000 68.490000 180.100000 ;
        RECT 68.290000 180.300000 68.490000 180.500000 ;
        RECT 68.290000 180.700000 68.490000 180.900000 ;
        RECT 68.290000 181.100000 68.490000 181.300000 ;
        RECT 68.290000 181.505000 68.490000 181.705000 ;
        RECT 68.290000 181.910000 68.490000 182.110000 ;
        RECT 68.290000 182.315000 68.490000 182.515000 ;
        RECT 68.290000 182.720000 68.490000 182.920000 ;
        RECT 68.290000 183.125000 68.490000 183.325000 ;
        RECT 68.290000 183.530000 68.490000 183.730000 ;
        RECT 68.290000 183.935000 68.490000 184.135000 ;
        RECT 68.290000 184.340000 68.490000 184.540000 ;
        RECT 68.290000 184.745000 68.490000 184.945000 ;
        RECT 68.290000 185.150000 68.490000 185.350000 ;
        RECT 68.290000 185.555000 68.490000 185.755000 ;
        RECT 68.290000 185.960000 68.490000 186.160000 ;
        RECT 68.290000 186.365000 68.490000 186.565000 ;
        RECT 68.290000 186.770000 68.490000 186.970000 ;
        RECT 68.290000 187.175000 68.490000 187.375000 ;
        RECT 68.290000 187.580000 68.490000 187.780000 ;
        RECT 68.290000 187.985000 68.490000 188.185000 ;
        RECT 68.290000 188.390000 68.490000 188.590000 ;
        RECT 68.290000 188.795000 68.490000 188.995000 ;
        RECT 68.290000 189.200000 68.490000 189.400000 ;
        RECT 68.290000 189.605000 68.490000 189.805000 ;
        RECT 68.290000 190.010000 68.490000 190.210000 ;
        RECT 68.290000 190.415000 68.490000 190.615000 ;
        RECT 68.290000 190.820000 68.490000 191.020000 ;
        RECT 68.290000 191.225000 68.490000 191.425000 ;
        RECT 68.290000 191.630000 68.490000 191.830000 ;
        RECT 68.290000 192.035000 68.490000 192.235000 ;
        RECT 68.290000 192.440000 68.490000 192.640000 ;
        RECT 68.290000 192.845000 68.490000 193.045000 ;
        RECT 68.290000 193.250000 68.490000 193.450000 ;
        RECT 68.290000 193.655000 68.490000 193.855000 ;
        RECT 68.290000 194.060000 68.490000 194.260000 ;
        RECT 68.290000 194.465000 68.490000 194.665000 ;
        RECT 68.290000 194.870000 68.490000 195.070000 ;
        RECT 68.290000 195.275000 68.490000 195.475000 ;
        RECT 68.290000 195.680000 68.490000 195.880000 ;
        RECT 68.290000 196.085000 68.490000 196.285000 ;
        RECT 68.290000 196.490000 68.490000 196.690000 ;
        RECT 68.290000 196.895000 68.490000 197.095000 ;
        RECT 68.290000 197.300000 68.490000 197.500000 ;
        RECT 68.290000 197.705000 68.490000 197.905000 ;
        RECT 68.330000  23.910000 68.530000  24.110000 ;
        RECT 68.330000  24.340000 68.530000  24.540000 ;
        RECT 68.330000  24.770000 68.530000  24.970000 ;
        RECT 68.330000  25.200000 68.530000  25.400000 ;
        RECT 68.330000  25.630000 68.530000  25.830000 ;
        RECT 68.330000  26.060000 68.530000  26.260000 ;
        RECT 68.330000  26.490000 68.530000  26.690000 ;
        RECT 68.330000  26.920000 68.530000  27.120000 ;
        RECT 68.330000  27.350000 68.530000  27.550000 ;
        RECT 68.330000  27.780000 68.530000  27.980000 ;
        RECT 68.330000  28.210000 68.530000  28.410000 ;
        RECT 68.700000 173.900000 68.900000 174.100000 ;
        RECT 68.700000 174.300000 68.900000 174.500000 ;
        RECT 68.700000 174.700000 68.900000 174.900000 ;
        RECT 68.700000 175.100000 68.900000 175.300000 ;
        RECT 68.700000 175.500000 68.900000 175.700000 ;
        RECT 68.700000 175.900000 68.900000 176.100000 ;
        RECT 68.700000 176.300000 68.900000 176.500000 ;
        RECT 68.700000 176.700000 68.900000 176.900000 ;
        RECT 68.700000 177.100000 68.900000 177.300000 ;
        RECT 68.700000 177.500000 68.900000 177.700000 ;
        RECT 68.700000 177.900000 68.900000 178.100000 ;
        RECT 68.700000 178.300000 68.900000 178.500000 ;
        RECT 68.700000 178.700000 68.900000 178.900000 ;
        RECT 68.700000 179.100000 68.900000 179.300000 ;
        RECT 68.700000 179.500000 68.900000 179.700000 ;
        RECT 68.700000 179.900000 68.900000 180.100000 ;
        RECT 68.700000 180.300000 68.900000 180.500000 ;
        RECT 68.700000 180.700000 68.900000 180.900000 ;
        RECT 68.700000 181.100000 68.900000 181.300000 ;
        RECT 68.700000 181.505000 68.900000 181.705000 ;
        RECT 68.700000 181.910000 68.900000 182.110000 ;
        RECT 68.700000 182.315000 68.900000 182.515000 ;
        RECT 68.700000 182.720000 68.900000 182.920000 ;
        RECT 68.700000 183.125000 68.900000 183.325000 ;
        RECT 68.700000 183.530000 68.900000 183.730000 ;
        RECT 68.700000 183.935000 68.900000 184.135000 ;
        RECT 68.700000 184.340000 68.900000 184.540000 ;
        RECT 68.700000 184.745000 68.900000 184.945000 ;
        RECT 68.700000 185.150000 68.900000 185.350000 ;
        RECT 68.700000 185.555000 68.900000 185.755000 ;
        RECT 68.700000 185.960000 68.900000 186.160000 ;
        RECT 68.700000 186.365000 68.900000 186.565000 ;
        RECT 68.700000 186.770000 68.900000 186.970000 ;
        RECT 68.700000 187.175000 68.900000 187.375000 ;
        RECT 68.700000 187.580000 68.900000 187.780000 ;
        RECT 68.700000 187.985000 68.900000 188.185000 ;
        RECT 68.700000 188.390000 68.900000 188.590000 ;
        RECT 68.700000 188.795000 68.900000 188.995000 ;
        RECT 68.700000 189.200000 68.900000 189.400000 ;
        RECT 68.700000 189.605000 68.900000 189.805000 ;
        RECT 68.700000 190.010000 68.900000 190.210000 ;
        RECT 68.700000 190.415000 68.900000 190.615000 ;
        RECT 68.700000 190.820000 68.900000 191.020000 ;
        RECT 68.700000 191.225000 68.900000 191.425000 ;
        RECT 68.700000 191.630000 68.900000 191.830000 ;
        RECT 68.700000 192.035000 68.900000 192.235000 ;
        RECT 68.700000 192.440000 68.900000 192.640000 ;
        RECT 68.700000 192.845000 68.900000 193.045000 ;
        RECT 68.700000 193.250000 68.900000 193.450000 ;
        RECT 68.700000 193.655000 68.900000 193.855000 ;
        RECT 68.700000 194.060000 68.900000 194.260000 ;
        RECT 68.700000 194.465000 68.900000 194.665000 ;
        RECT 68.700000 194.870000 68.900000 195.070000 ;
        RECT 68.700000 195.275000 68.900000 195.475000 ;
        RECT 68.700000 195.680000 68.900000 195.880000 ;
        RECT 68.700000 196.085000 68.900000 196.285000 ;
        RECT 68.700000 196.490000 68.900000 196.690000 ;
        RECT 68.700000 196.895000 68.900000 197.095000 ;
        RECT 68.700000 197.300000 68.900000 197.500000 ;
        RECT 68.700000 197.705000 68.900000 197.905000 ;
        RECT 68.735000  23.910000 68.935000  24.110000 ;
        RECT 68.735000  24.340000 68.935000  24.540000 ;
        RECT 68.735000  24.770000 68.935000  24.970000 ;
        RECT 68.735000  25.200000 68.935000  25.400000 ;
        RECT 68.735000  25.630000 68.935000  25.830000 ;
        RECT 68.735000  26.060000 68.935000  26.260000 ;
        RECT 68.735000  26.490000 68.935000  26.690000 ;
        RECT 68.735000  26.920000 68.935000  27.120000 ;
        RECT 68.735000  27.350000 68.935000  27.550000 ;
        RECT 68.735000  27.780000 68.935000  27.980000 ;
        RECT 68.735000  28.210000 68.935000  28.410000 ;
        RECT 69.110000 173.900000 69.310000 174.100000 ;
        RECT 69.110000 174.300000 69.310000 174.500000 ;
        RECT 69.110000 174.700000 69.310000 174.900000 ;
        RECT 69.110000 175.100000 69.310000 175.300000 ;
        RECT 69.110000 175.500000 69.310000 175.700000 ;
        RECT 69.110000 175.900000 69.310000 176.100000 ;
        RECT 69.110000 176.300000 69.310000 176.500000 ;
        RECT 69.110000 176.700000 69.310000 176.900000 ;
        RECT 69.110000 177.100000 69.310000 177.300000 ;
        RECT 69.110000 177.500000 69.310000 177.700000 ;
        RECT 69.110000 177.900000 69.310000 178.100000 ;
        RECT 69.110000 178.300000 69.310000 178.500000 ;
        RECT 69.110000 178.700000 69.310000 178.900000 ;
        RECT 69.110000 179.100000 69.310000 179.300000 ;
        RECT 69.110000 179.500000 69.310000 179.700000 ;
        RECT 69.110000 179.900000 69.310000 180.100000 ;
        RECT 69.110000 180.300000 69.310000 180.500000 ;
        RECT 69.110000 180.700000 69.310000 180.900000 ;
        RECT 69.110000 181.100000 69.310000 181.300000 ;
        RECT 69.110000 181.505000 69.310000 181.705000 ;
        RECT 69.110000 181.910000 69.310000 182.110000 ;
        RECT 69.110000 182.315000 69.310000 182.515000 ;
        RECT 69.110000 182.720000 69.310000 182.920000 ;
        RECT 69.110000 183.125000 69.310000 183.325000 ;
        RECT 69.110000 183.530000 69.310000 183.730000 ;
        RECT 69.110000 183.935000 69.310000 184.135000 ;
        RECT 69.110000 184.340000 69.310000 184.540000 ;
        RECT 69.110000 184.745000 69.310000 184.945000 ;
        RECT 69.110000 185.150000 69.310000 185.350000 ;
        RECT 69.110000 185.555000 69.310000 185.755000 ;
        RECT 69.110000 185.960000 69.310000 186.160000 ;
        RECT 69.110000 186.365000 69.310000 186.565000 ;
        RECT 69.110000 186.770000 69.310000 186.970000 ;
        RECT 69.110000 187.175000 69.310000 187.375000 ;
        RECT 69.110000 187.580000 69.310000 187.780000 ;
        RECT 69.110000 187.985000 69.310000 188.185000 ;
        RECT 69.110000 188.390000 69.310000 188.590000 ;
        RECT 69.110000 188.795000 69.310000 188.995000 ;
        RECT 69.110000 189.200000 69.310000 189.400000 ;
        RECT 69.110000 189.605000 69.310000 189.805000 ;
        RECT 69.110000 190.010000 69.310000 190.210000 ;
        RECT 69.110000 190.415000 69.310000 190.615000 ;
        RECT 69.110000 190.820000 69.310000 191.020000 ;
        RECT 69.110000 191.225000 69.310000 191.425000 ;
        RECT 69.110000 191.630000 69.310000 191.830000 ;
        RECT 69.110000 192.035000 69.310000 192.235000 ;
        RECT 69.110000 192.440000 69.310000 192.640000 ;
        RECT 69.110000 192.845000 69.310000 193.045000 ;
        RECT 69.110000 193.250000 69.310000 193.450000 ;
        RECT 69.110000 193.655000 69.310000 193.855000 ;
        RECT 69.110000 194.060000 69.310000 194.260000 ;
        RECT 69.110000 194.465000 69.310000 194.665000 ;
        RECT 69.110000 194.870000 69.310000 195.070000 ;
        RECT 69.110000 195.275000 69.310000 195.475000 ;
        RECT 69.110000 195.680000 69.310000 195.880000 ;
        RECT 69.110000 196.085000 69.310000 196.285000 ;
        RECT 69.110000 196.490000 69.310000 196.690000 ;
        RECT 69.110000 196.895000 69.310000 197.095000 ;
        RECT 69.110000 197.300000 69.310000 197.500000 ;
        RECT 69.110000 197.705000 69.310000 197.905000 ;
        RECT 69.140000  23.910000 69.340000  24.110000 ;
        RECT 69.140000  24.340000 69.340000  24.540000 ;
        RECT 69.140000  24.770000 69.340000  24.970000 ;
        RECT 69.140000  25.200000 69.340000  25.400000 ;
        RECT 69.140000  25.630000 69.340000  25.830000 ;
        RECT 69.140000  26.060000 69.340000  26.260000 ;
        RECT 69.140000  26.490000 69.340000  26.690000 ;
        RECT 69.140000  26.920000 69.340000  27.120000 ;
        RECT 69.140000  27.350000 69.340000  27.550000 ;
        RECT 69.140000  27.780000 69.340000  27.980000 ;
        RECT 69.140000  28.210000 69.340000  28.410000 ;
        RECT 69.520000 173.900000 69.720000 174.100000 ;
        RECT 69.520000 174.300000 69.720000 174.500000 ;
        RECT 69.520000 174.700000 69.720000 174.900000 ;
        RECT 69.520000 175.100000 69.720000 175.300000 ;
        RECT 69.520000 175.500000 69.720000 175.700000 ;
        RECT 69.520000 175.900000 69.720000 176.100000 ;
        RECT 69.520000 176.300000 69.720000 176.500000 ;
        RECT 69.520000 176.700000 69.720000 176.900000 ;
        RECT 69.520000 177.100000 69.720000 177.300000 ;
        RECT 69.520000 177.500000 69.720000 177.700000 ;
        RECT 69.520000 177.900000 69.720000 178.100000 ;
        RECT 69.520000 178.300000 69.720000 178.500000 ;
        RECT 69.520000 178.700000 69.720000 178.900000 ;
        RECT 69.520000 179.100000 69.720000 179.300000 ;
        RECT 69.520000 179.500000 69.720000 179.700000 ;
        RECT 69.520000 179.900000 69.720000 180.100000 ;
        RECT 69.520000 180.300000 69.720000 180.500000 ;
        RECT 69.520000 180.700000 69.720000 180.900000 ;
        RECT 69.520000 181.100000 69.720000 181.300000 ;
        RECT 69.520000 181.505000 69.720000 181.705000 ;
        RECT 69.520000 181.910000 69.720000 182.110000 ;
        RECT 69.520000 182.315000 69.720000 182.515000 ;
        RECT 69.520000 182.720000 69.720000 182.920000 ;
        RECT 69.520000 183.125000 69.720000 183.325000 ;
        RECT 69.520000 183.530000 69.720000 183.730000 ;
        RECT 69.520000 183.935000 69.720000 184.135000 ;
        RECT 69.520000 184.340000 69.720000 184.540000 ;
        RECT 69.520000 184.745000 69.720000 184.945000 ;
        RECT 69.520000 185.150000 69.720000 185.350000 ;
        RECT 69.520000 185.555000 69.720000 185.755000 ;
        RECT 69.520000 185.960000 69.720000 186.160000 ;
        RECT 69.520000 186.365000 69.720000 186.565000 ;
        RECT 69.520000 186.770000 69.720000 186.970000 ;
        RECT 69.520000 187.175000 69.720000 187.375000 ;
        RECT 69.520000 187.580000 69.720000 187.780000 ;
        RECT 69.520000 187.985000 69.720000 188.185000 ;
        RECT 69.520000 188.390000 69.720000 188.590000 ;
        RECT 69.520000 188.795000 69.720000 188.995000 ;
        RECT 69.520000 189.200000 69.720000 189.400000 ;
        RECT 69.520000 189.605000 69.720000 189.805000 ;
        RECT 69.520000 190.010000 69.720000 190.210000 ;
        RECT 69.520000 190.415000 69.720000 190.615000 ;
        RECT 69.520000 190.820000 69.720000 191.020000 ;
        RECT 69.520000 191.225000 69.720000 191.425000 ;
        RECT 69.520000 191.630000 69.720000 191.830000 ;
        RECT 69.520000 192.035000 69.720000 192.235000 ;
        RECT 69.520000 192.440000 69.720000 192.640000 ;
        RECT 69.520000 192.845000 69.720000 193.045000 ;
        RECT 69.520000 193.250000 69.720000 193.450000 ;
        RECT 69.520000 193.655000 69.720000 193.855000 ;
        RECT 69.520000 194.060000 69.720000 194.260000 ;
        RECT 69.520000 194.465000 69.720000 194.665000 ;
        RECT 69.520000 194.870000 69.720000 195.070000 ;
        RECT 69.520000 195.275000 69.720000 195.475000 ;
        RECT 69.520000 195.680000 69.720000 195.880000 ;
        RECT 69.520000 196.085000 69.720000 196.285000 ;
        RECT 69.520000 196.490000 69.720000 196.690000 ;
        RECT 69.520000 196.895000 69.720000 197.095000 ;
        RECT 69.520000 197.300000 69.720000 197.500000 ;
        RECT 69.520000 197.705000 69.720000 197.905000 ;
        RECT 69.545000  23.910000 69.745000  24.110000 ;
        RECT 69.545000  24.340000 69.745000  24.540000 ;
        RECT 69.545000  24.770000 69.745000  24.970000 ;
        RECT 69.545000  25.200000 69.745000  25.400000 ;
        RECT 69.545000  25.630000 69.745000  25.830000 ;
        RECT 69.545000  26.060000 69.745000  26.260000 ;
        RECT 69.545000  26.490000 69.745000  26.690000 ;
        RECT 69.545000  26.920000 69.745000  27.120000 ;
        RECT 69.545000  27.350000 69.745000  27.550000 ;
        RECT 69.545000  27.780000 69.745000  27.980000 ;
        RECT 69.545000  28.210000 69.745000  28.410000 ;
        RECT 69.930000 173.900000 70.130000 174.100000 ;
        RECT 69.930000 174.300000 70.130000 174.500000 ;
        RECT 69.930000 174.700000 70.130000 174.900000 ;
        RECT 69.930000 175.100000 70.130000 175.300000 ;
        RECT 69.930000 175.500000 70.130000 175.700000 ;
        RECT 69.930000 175.900000 70.130000 176.100000 ;
        RECT 69.930000 176.300000 70.130000 176.500000 ;
        RECT 69.930000 176.700000 70.130000 176.900000 ;
        RECT 69.930000 177.100000 70.130000 177.300000 ;
        RECT 69.930000 177.500000 70.130000 177.700000 ;
        RECT 69.930000 177.900000 70.130000 178.100000 ;
        RECT 69.930000 178.300000 70.130000 178.500000 ;
        RECT 69.930000 178.700000 70.130000 178.900000 ;
        RECT 69.930000 179.100000 70.130000 179.300000 ;
        RECT 69.930000 179.500000 70.130000 179.700000 ;
        RECT 69.930000 179.900000 70.130000 180.100000 ;
        RECT 69.930000 180.300000 70.130000 180.500000 ;
        RECT 69.930000 180.700000 70.130000 180.900000 ;
        RECT 69.930000 181.100000 70.130000 181.300000 ;
        RECT 69.930000 181.505000 70.130000 181.705000 ;
        RECT 69.930000 181.910000 70.130000 182.110000 ;
        RECT 69.930000 182.315000 70.130000 182.515000 ;
        RECT 69.930000 182.720000 70.130000 182.920000 ;
        RECT 69.930000 183.125000 70.130000 183.325000 ;
        RECT 69.930000 183.530000 70.130000 183.730000 ;
        RECT 69.930000 183.935000 70.130000 184.135000 ;
        RECT 69.930000 184.340000 70.130000 184.540000 ;
        RECT 69.930000 184.745000 70.130000 184.945000 ;
        RECT 69.930000 185.150000 70.130000 185.350000 ;
        RECT 69.930000 185.555000 70.130000 185.755000 ;
        RECT 69.930000 185.960000 70.130000 186.160000 ;
        RECT 69.930000 186.365000 70.130000 186.565000 ;
        RECT 69.930000 186.770000 70.130000 186.970000 ;
        RECT 69.930000 187.175000 70.130000 187.375000 ;
        RECT 69.930000 187.580000 70.130000 187.780000 ;
        RECT 69.930000 187.985000 70.130000 188.185000 ;
        RECT 69.930000 188.390000 70.130000 188.590000 ;
        RECT 69.930000 188.795000 70.130000 188.995000 ;
        RECT 69.930000 189.200000 70.130000 189.400000 ;
        RECT 69.930000 189.605000 70.130000 189.805000 ;
        RECT 69.930000 190.010000 70.130000 190.210000 ;
        RECT 69.930000 190.415000 70.130000 190.615000 ;
        RECT 69.930000 190.820000 70.130000 191.020000 ;
        RECT 69.930000 191.225000 70.130000 191.425000 ;
        RECT 69.930000 191.630000 70.130000 191.830000 ;
        RECT 69.930000 192.035000 70.130000 192.235000 ;
        RECT 69.930000 192.440000 70.130000 192.640000 ;
        RECT 69.930000 192.845000 70.130000 193.045000 ;
        RECT 69.930000 193.250000 70.130000 193.450000 ;
        RECT 69.930000 193.655000 70.130000 193.855000 ;
        RECT 69.930000 194.060000 70.130000 194.260000 ;
        RECT 69.930000 194.465000 70.130000 194.665000 ;
        RECT 69.930000 194.870000 70.130000 195.070000 ;
        RECT 69.930000 195.275000 70.130000 195.475000 ;
        RECT 69.930000 195.680000 70.130000 195.880000 ;
        RECT 69.930000 196.085000 70.130000 196.285000 ;
        RECT 69.930000 196.490000 70.130000 196.690000 ;
        RECT 69.930000 196.895000 70.130000 197.095000 ;
        RECT 69.930000 197.300000 70.130000 197.500000 ;
        RECT 69.930000 197.705000 70.130000 197.905000 ;
        RECT 69.950000  23.910000 70.150000  24.110000 ;
        RECT 69.950000  24.340000 70.150000  24.540000 ;
        RECT 69.950000  24.770000 70.150000  24.970000 ;
        RECT 69.950000  25.200000 70.150000  25.400000 ;
        RECT 69.950000  25.630000 70.150000  25.830000 ;
        RECT 69.950000  26.060000 70.150000  26.260000 ;
        RECT 69.950000  26.490000 70.150000  26.690000 ;
        RECT 69.950000  26.920000 70.150000  27.120000 ;
        RECT 69.950000  27.350000 70.150000  27.550000 ;
        RECT 69.950000  27.780000 70.150000  27.980000 ;
        RECT 69.950000  28.210000 70.150000  28.410000 ;
        RECT 70.340000 173.900000 70.540000 174.100000 ;
        RECT 70.340000 174.300000 70.540000 174.500000 ;
        RECT 70.340000 174.700000 70.540000 174.900000 ;
        RECT 70.340000 175.100000 70.540000 175.300000 ;
        RECT 70.340000 175.500000 70.540000 175.700000 ;
        RECT 70.340000 175.900000 70.540000 176.100000 ;
        RECT 70.340000 176.300000 70.540000 176.500000 ;
        RECT 70.340000 176.700000 70.540000 176.900000 ;
        RECT 70.340000 177.100000 70.540000 177.300000 ;
        RECT 70.340000 177.500000 70.540000 177.700000 ;
        RECT 70.340000 177.900000 70.540000 178.100000 ;
        RECT 70.340000 178.300000 70.540000 178.500000 ;
        RECT 70.340000 178.700000 70.540000 178.900000 ;
        RECT 70.340000 179.100000 70.540000 179.300000 ;
        RECT 70.340000 179.500000 70.540000 179.700000 ;
        RECT 70.340000 179.900000 70.540000 180.100000 ;
        RECT 70.340000 180.300000 70.540000 180.500000 ;
        RECT 70.340000 180.700000 70.540000 180.900000 ;
        RECT 70.340000 181.100000 70.540000 181.300000 ;
        RECT 70.340000 181.505000 70.540000 181.705000 ;
        RECT 70.340000 181.910000 70.540000 182.110000 ;
        RECT 70.340000 182.315000 70.540000 182.515000 ;
        RECT 70.340000 182.720000 70.540000 182.920000 ;
        RECT 70.340000 183.125000 70.540000 183.325000 ;
        RECT 70.340000 183.530000 70.540000 183.730000 ;
        RECT 70.340000 183.935000 70.540000 184.135000 ;
        RECT 70.340000 184.340000 70.540000 184.540000 ;
        RECT 70.340000 184.745000 70.540000 184.945000 ;
        RECT 70.340000 185.150000 70.540000 185.350000 ;
        RECT 70.340000 185.555000 70.540000 185.755000 ;
        RECT 70.340000 185.960000 70.540000 186.160000 ;
        RECT 70.340000 186.365000 70.540000 186.565000 ;
        RECT 70.340000 186.770000 70.540000 186.970000 ;
        RECT 70.340000 187.175000 70.540000 187.375000 ;
        RECT 70.340000 187.580000 70.540000 187.780000 ;
        RECT 70.340000 187.985000 70.540000 188.185000 ;
        RECT 70.340000 188.390000 70.540000 188.590000 ;
        RECT 70.340000 188.795000 70.540000 188.995000 ;
        RECT 70.340000 189.200000 70.540000 189.400000 ;
        RECT 70.340000 189.605000 70.540000 189.805000 ;
        RECT 70.340000 190.010000 70.540000 190.210000 ;
        RECT 70.340000 190.415000 70.540000 190.615000 ;
        RECT 70.340000 190.820000 70.540000 191.020000 ;
        RECT 70.340000 191.225000 70.540000 191.425000 ;
        RECT 70.340000 191.630000 70.540000 191.830000 ;
        RECT 70.340000 192.035000 70.540000 192.235000 ;
        RECT 70.340000 192.440000 70.540000 192.640000 ;
        RECT 70.340000 192.845000 70.540000 193.045000 ;
        RECT 70.340000 193.250000 70.540000 193.450000 ;
        RECT 70.340000 193.655000 70.540000 193.855000 ;
        RECT 70.340000 194.060000 70.540000 194.260000 ;
        RECT 70.340000 194.465000 70.540000 194.665000 ;
        RECT 70.340000 194.870000 70.540000 195.070000 ;
        RECT 70.340000 195.275000 70.540000 195.475000 ;
        RECT 70.340000 195.680000 70.540000 195.880000 ;
        RECT 70.340000 196.085000 70.540000 196.285000 ;
        RECT 70.340000 196.490000 70.540000 196.690000 ;
        RECT 70.340000 196.895000 70.540000 197.095000 ;
        RECT 70.340000 197.300000 70.540000 197.500000 ;
        RECT 70.340000 197.705000 70.540000 197.905000 ;
        RECT 70.355000  23.910000 70.555000  24.110000 ;
        RECT 70.355000  24.340000 70.555000  24.540000 ;
        RECT 70.355000  24.770000 70.555000  24.970000 ;
        RECT 70.355000  25.200000 70.555000  25.400000 ;
        RECT 70.355000  25.630000 70.555000  25.830000 ;
        RECT 70.355000  26.060000 70.555000  26.260000 ;
        RECT 70.355000  26.490000 70.555000  26.690000 ;
        RECT 70.355000  26.920000 70.555000  27.120000 ;
        RECT 70.355000  27.350000 70.555000  27.550000 ;
        RECT 70.355000  27.780000 70.555000  27.980000 ;
        RECT 70.355000  28.210000 70.555000  28.410000 ;
        RECT 70.750000 173.900000 70.950000 174.100000 ;
        RECT 70.750000 174.300000 70.950000 174.500000 ;
        RECT 70.750000 174.700000 70.950000 174.900000 ;
        RECT 70.750000 175.100000 70.950000 175.300000 ;
        RECT 70.750000 175.500000 70.950000 175.700000 ;
        RECT 70.750000 175.900000 70.950000 176.100000 ;
        RECT 70.750000 176.300000 70.950000 176.500000 ;
        RECT 70.750000 176.700000 70.950000 176.900000 ;
        RECT 70.750000 177.100000 70.950000 177.300000 ;
        RECT 70.750000 177.500000 70.950000 177.700000 ;
        RECT 70.750000 177.900000 70.950000 178.100000 ;
        RECT 70.750000 178.300000 70.950000 178.500000 ;
        RECT 70.750000 178.700000 70.950000 178.900000 ;
        RECT 70.750000 179.100000 70.950000 179.300000 ;
        RECT 70.750000 179.500000 70.950000 179.700000 ;
        RECT 70.750000 179.900000 70.950000 180.100000 ;
        RECT 70.750000 180.300000 70.950000 180.500000 ;
        RECT 70.750000 180.700000 70.950000 180.900000 ;
        RECT 70.750000 181.100000 70.950000 181.300000 ;
        RECT 70.750000 181.505000 70.950000 181.705000 ;
        RECT 70.750000 181.910000 70.950000 182.110000 ;
        RECT 70.750000 182.315000 70.950000 182.515000 ;
        RECT 70.750000 182.720000 70.950000 182.920000 ;
        RECT 70.750000 183.125000 70.950000 183.325000 ;
        RECT 70.750000 183.530000 70.950000 183.730000 ;
        RECT 70.750000 183.935000 70.950000 184.135000 ;
        RECT 70.750000 184.340000 70.950000 184.540000 ;
        RECT 70.750000 184.745000 70.950000 184.945000 ;
        RECT 70.750000 185.150000 70.950000 185.350000 ;
        RECT 70.750000 185.555000 70.950000 185.755000 ;
        RECT 70.750000 185.960000 70.950000 186.160000 ;
        RECT 70.750000 186.365000 70.950000 186.565000 ;
        RECT 70.750000 186.770000 70.950000 186.970000 ;
        RECT 70.750000 187.175000 70.950000 187.375000 ;
        RECT 70.750000 187.580000 70.950000 187.780000 ;
        RECT 70.750000 187.985000 70.950000 188.185000 ;
        RECT 70.750000 188.390000 70.950000 188.590000 ;
        RECT 70.750000 188.795000 70.950000 188.995000 ;
        RECT 70.750000 189.200000 70.950000 189.400000 ;
        RECT 70.750000 189.605000 70.950000 189.805000 ;
        RECT 70.750000 190.010000 70.950000 190.210000 ;
        RECT 70.750000 190.415000 70.950000 190.615000 ;
        RECT 70.750000 190.820000 70.950000 191.020000 ;
        RECT 70.750000 191.225000 70.950000 191.425000 ;
        RECT 70.750000 191.630000 70.950000 191.830000 ;
        RECT 70.750000 192.035000 70.950000 192.235000 ;
        RECT 70.750000 192.440000 70.950000 192.640000 ;
        RECT 70.750000 192.845000 70.950000 193.045000 ;
        RECT 70.750000 193.250000 70.950000 193.450000 ;
        RECT 70.750000 193.655000 70.950000 193.855000 ;
        RECT 70.750000 194.060000 70.950000 194.260000 ;
        RECT 70.750000 194.465000 70.950000 194.665000 ;
        RECT 70.750000 194.870000 70.950000 195.070000 ;
        RECT 70.750000 195.275000 70.950000 195.475000 ;
        RECT 70.750000 195.680000 70.950000 195.880000 ;
        RECT 70.750000 196.085000 70.950000 196.285000 ;
        RECT 70.750000 196.490000 70.950000 196.690000 ;
        RECT 70.750000 196.895000 70.950000 197.095000 ;
        RECT 70.750000 197.300000 70.950000 197.500000 ;
        RECT 70.750000 197.705000 70.950000 197.905000 ;
        RECT 70.760000  23.910000 70.960000  24.110000 ;
        RECT 70.760000  24.340000 70.960000  24.540000 ;
        RECT 70.760000  24.770000 70.960000  24.970000 ;
        RECT 70.760000  25.200000 70.960000  25.400000 ;
        RECT 70.760000  25.630000 70.960000  25.830000 ;
        RECT 70.760000  26.060000 70.960000  26.260000 ;
        RECT 70.760000  26.490000 70.960000  26.690000 ;
        RECT 70.760000  26.920000 70.960000  27.120000 ;
        RECT 70.760000  27.350000 70.960000  27.550000 ;
        RECT 70.760000  27.780000 70.960000  27.980000 ;
        RECT 70.760000  28.210000 70.960000  28.410000 ;
        RECT 71.160000 173.900000 71.360000 174.100000 ;
        RECT 71.160000 174.300000 71.360000 174.500000 ;
        RECT 71.160000 174.700000 71.360000 174.900000 ;
        RECT 71.160000 175.100000 71.360000 175.300000 ;
        RECT 71.160000 175.500000 71.360000 175.700000 ;
        RECT 71.160000 175.900000 71.360000 176.100000 ;
        RECT 71.160000 176.300000 71.360000 176.500000 ;
        RECT 71.160000 176.700000 71.360000 176.900000 ;
        RECT 71.160000 177.100000 71.360000 177.300000 ;
        RECT 71.160000 177.500000 71.360000 177.700000 ;
        RECT 71.160000 177.900000 71.360000 178.100000 ;
        RECT 71.160000 178.300000 71.360000 178.500000 ;
        RECT 71.160000 178.700000 71.360000 178.900000 ;
        RECT 71.160000 179.100000 71.360000 179.300000 ;
        RECT 71.160000 179.500000 71.360000 179.700000 ;
        RECT 71.160000 179.900000 71.360000 180.100000 ;
        RECT 71.160000 180.300000 71.360000 180.500000 ;
        RECT 71.160000 180.700000 71.360000 180.900000 ;
        RECT 71.160000 181.100000 71.360000 181.300000 ;
        RECT 71.160000 181.505000 71.360000 181.705000 ;
        RECT 71.160000 181.910000 71.360000 182.110000 ;
        RECT 71.160000 182.315000 71.360000 182.515000 ;
        RECT 71.160000 182.720000 71.360000 182.920000 ;
        RECT 71.160000 183.125000 71.360000 183.325000 ;
        RECT 71.160000 183.530000 71.360000 183.730000 ;
        RECT 71.160000 183.935000 71.360000 184.135000 ;
        RECT 71.160000 184.340000 71.360000 184.540000 ;
        RECT 71.160000 184.745000 71.360000 184.945000 ;
        RECT 71.160000 185.150000 71.360000 185.350000 ;
        RECT 71.160000 185.555000 71.360000 185.755000 ;
        RECT 71.160000 185.960000 71.360000 186.160000 ;
        RECT 71.160000 186.365000 71.360000 186.565000 ;
        RECT 71.160000 186.770000 71.360000 186.970000 ;
        RECT 71.160000 187.175000 71.360000 187.375000 ;
        RECT 71.160000 187.580000 71.360000 187.780000 ;
        RECT 71.160000 187.985000 71.360000 188.185000 ;
        RECT 71.160000 188.390000 71.360000 188.590000 ;
        RECT 71.160000 188.795000 71.360000 188.995000 ;
        RECT 71.160000 189.200000 71.360000 189.400000 ;
        RECT 71.160000 189.605000 71.360000 189.805000 ;
        RECT 71.160000 190.010000 71.360000 190.210000 ;
        RECT 71.160000 190.415000 71.360000 190.615000 ;
        RECT 71.160000 190.820000 71.360000 191.020000 ;
        RECT 71.160000 191.225000 71.360000 191.425000 ;
        RECT 71.160000 191.630000 71.360000 191.830000 ;
        RECT 71.160000 192.035000 71.360000 192.235000 ;
        RECT 71.160000 192.440000 71.360000 192.640000 ;
        RECT 71.160000 192.845000 71.360000 193.045000 ;
        RECT 71.160000 193.250000 71.360000 193.450000 ;
        RECT 71.160000 193.655000 71.360000 193.855000 ;
        RECT 71.160000 194.060000 71.360000 194.260000 ;
        RECT 71.160000 194.465000 71.360000 194.665000 ;
        RECT 71.160000 194.870000 71.360000 195.070000 ;
        RECT 71.160000 195.275000 71.360000 195.475000 ;
        RECT 71.160000 195.680000 71.360000 195.880000 ;
        RECT 71.160000 196.085000 71.360000 196.285000 ;
        RECT 71.160000 196.490000 71.360000 196.690000 ;
        RECT 71.160000 196.895000 71.360000 197.095000 ;
        RECT 71.160000 197.300000 71.360000 197.500000 ;
        RECT 71.160000 197.705000 71.360000 197.905000 ;
        RECT 71.165000  23.910000 71.365000  24.110000 ;
        RECT 71.165000  24.340000 71.365000  24.540000 ;
        RECT 71.165000  24.770000 71.365000  24.970000 ;
        RECT 71.165000  25.200000 71.365000  25.400000 ;
        RECT 71.165000  25.630000 71.365000  25.830000 ;
        RECT 71.165000  26.060000 71.365000  26.260000 ;
        RECT 71.165000  26.490000 71.365000  26.690000 ;
        RECT 71.165000  26.920000 71.365000  27.120000 ;
        RECT 71.165000  27.350000 71.365000  27.550000 ;
        RECT 71.165000  27.780000 71.365000  27.980000 ;
        RECT 71.165000  28.210000 71.365000  28.410000 ;
        RECT 71.570000  23.910000 71.770000  24.110000 ;
        RECT 71.570000  24.340000 71.770000  24.540000 ;
        RECT 71.570000  24.770000 71.770000  24.970000 ;
        RECT 71.570000  25.200000 71.770000  25.400000 ;
        RECT 71.570000  25.630000 71.770000  25.830000 ;
        RECT 71.570000  26.060000 71.770000  26.260000 ;
        RECT 71.570000  26.490000 71.770000  26.690000 ;
        RECT 71.570000  26.920000 71.770000  27.120000 ;
        RECT 71.570000  27.350000 71.770000  27.550000 ;
        RECT 71.570000  27.780000 71.770000  27.980000 ;
        RECT 71.570000  28.210000 71.770000  28.410000 ;
        RECT 71.570000 173.900000 71.770000 174.100000 ;
        RECT 71.570000 174.300000 71.770000 174.500000 ;
        RECT 71.570000 174.700000 71.770000 174.900000 ;
        RECT 71.570000 175.100000 71.770000 175.300000 ;
        RECT 71.570000 175.500000 71.770000 175.700000 ;
        RECT 71.570000 175.900000 71.770000 176.100000 ;
        RECT 71.570000 176.300000 71.770000 176.500000 ;
        RECT 71.570000 176.700000 71.770000 176.900000 ;
        RECT 71.570000 177.100000 71.770000 177.300000 ;
        RECT 71.570000 177.500000 71.770000 177.700000 ;
        RECT 71.570000 177.900000 71.770000 178.100000 ;
        RECT 71.570000 178.300000 71.770000 178.500000 ;
        RECT 71.570000 178.700000 71.770000 178.900000 ;
        RECT 71.570000 179.100000 71.770000 179.300000 ;
        RECT 71.570000 179.500000 71.770000 179.700000 ;
        RECT 71.570000 179.900000 71.770000 180.100000 ;
        RECT 71.570000 180.300000 71.770000 180.500000 ;
        RECT 71.570000 180.700000 71.770000 180.900000 ;
        RECT 71.570000 181.100000 71.770000 181.300000 ;
        RECT 71.570000 181.505000 71.770000 181.705000 ;
        RECT 71.570000 181.910000 71.770000 182.110000 ;
        RECT 71.570000 182.315000 71.770000 182.515000 ;
        RECT 71.570000 182.720000 71.770000 182.920000 ;
        RECT 71.570000 183.125000 71.770000 183.325000 ;
        RECT 71.570000 183.530000 71.770000 183.730000 ;
        RECT 71.570000 183.935000 71.770000 184.135000 ;
        RECT 71.570000 184.340000 71.770000 184.540000 ;
        RECT 71.570000 184.745000 71.770000 184.945000 ;
        RECT 71.570000 185.150000 71.770000 185.350000 ;
        RECT 71.570000 185.555000 71.770000 185.755000 ;
        RECT 71.570000 185.960000 71.770000 186.160000 ;
        RECT 71.570000 186.365000 71.770000 186.565000 ;
        RECT 71.570000 186.770000 71.770000 186.970000 ;
        RECT 71.570000 187.175000 71.770000 187.375000 ;
        RECT 71.570000 187.580000 71.770000 187.780000 ;
        RECT 71.570000 187.985000 71.770000 188.185000 ;
        RECT 71.570000 188.390000 71.770000 188.590000 ;
        RECT 71.570000 188.795000 71.770000 188.995000 ;
        RECT 71.570000 189.200000 71.770000 189.400000 ;
        RECT 71.570000 189.605000 71.770000 189.805000 ;
        RECT 71.570000 190.010000 71.770000 190.210000 ;
        RECT 71.570000 190.415000 71.770000 190.615000 ;
        RECT 71.570000 190.820000 71.770000 191.020000 ;
        RECT 71.570000 191.225000 71.770000 191.425000 ;
        RECT 71.570000 191.630000 71.770000 191.830000 ;
        RECT 71.570000 192.035000 71.770000 192.235000 ;
        RECT 71.570000 192.440000 71.770000 192.640000 ;
        RECT 71.570000 192.845000 71.770000 193.045000 ;
        RECT 71.570000 193.250000 71.770000 193.450000 ;
        RECT 71.570000 193.655000 71.770000 193.855000 ;
        RECT 71.570000 194.060000 71.770000 194.260000 ;
        RECT 71.570000 194.465000 71.770000 194.665000 ;
        RECT 71.570000 194.870000 71.770000 195.070000 ;
        RECT 71.570000 195.275000 71.770000 195.475000 ;
        RECT 71.570000 195.680000 71.770000 195.880000 ;
        RECT 71.570000 196.085000 71.770000 196.285000 ;
        RECT 71.570000 196.490000 71.770000 196.690000 ;
        RECT 71.570000 196.895000 71.770000 197.095000 ;
        RECT 71.570000 197.300000 71.770000 197.500000 ;
        RECT 71.570000 197.705000 71.770000 197.905000 ;
        RECT 71.975000  23.910000 72.175000  24.110000 ;
        RECT 71.975000  24.340000 72.175000  24.540000 ;
        RECT 71.975000  24.770000 72.175000  24.970000 ;
        RECT 71.975000  25.200000 72.175000  25.400000 ;
        RECT 71.975000  25.630000 72.175000  25.830000 ;
        RECT 71.975000  26.060000 72.175000  26.260000 ;
        RECT 71.975000  26.490000 72.175000  26.690000 ;
        RECT 71.975000  26.920000 72.175000  27.120000 ;
        RECT 71.975000  27.350000 72.175000  27.550000 ;
        RECT 71.975000  27.780000 72.175000  27.980000 ;
        RECT 71.975000  28.210000 72.175000  28.410000 ;
        RECT 71.980000 173.900000 72.180000 174.100000 ;
        RECT 71.980000 174.300000 72.180000 174.500000 ;
        RECT 71.980000 174.700000 72.180000 174.900000 ;
        RECT 71.980000 175.100000 72.180000 175.300000 ;
        RECT 71.980000 175.500000 72.180000 175.700000 ;
        RECT 71.980000 175.900000 72.180000 176.100000 ;
        RECT 71.980000 176.300000 72.180000 176.500000 ;
        RECT 71.980000 176.700000 72.180000 176.900000 ;
        RECT 71.980000 177.100000 72.180000 177.300000 ;
        RECT 71.980000 177.500000 72.180000 177.700000 ;
        RECT 71.980000 177.900000 72.180000 178.100000 ;
        RECT 71.980000 178.300000 72.180000 178.500000 ;
        RECT 71.980000 178.700000 72.180000 178.900000 ;
        RECT 71.980000 179.100000 72.180000 179.300000 ;
        RECT 71.980000 179.500000 72.180000 179.700000 ;
        RECT 71.980000 179.900000 72.180000 180.100000 ;
        RECT 71.980000 180.300000 72.180000 180.500000 ;
        RECT 71.980000 180.700000 72.180000 180.900000 ;
        RECT 71.980000 181.100000 72.180000 181.300000 ;
        RECT 71.980000 181.505000 72.180000 181.705000 ;
        RECT 71.980000 181.910000 72.180000 182.110000 ;
        RECT 71.980000 182.315000 72.180000 182.515000 ;
        RECT 71.980000 182.720000 72.180000 182.920000 ;
        RECT 71.980000 183.125000 72.180000 183.325000 ;
        RECT 71.980000 183.530000 72.180000 183.730000 ;
        RECT 71.980000 183.935000 72.180000 184.135000 ;
        RECT 71.980000 184.340000 72.180000 184.540000 ;
        RECT 71.980000 184.745000 72.180000 184.945000 ;
        RECT 71.980000 185.150000 72.180000 185.350000 ;
        RECT 71.980000 185.555000 72.180000 185.755000 ;
        RECT 71.980000 185.960000 72.180000 186.160000 ;
        RECT 71.980000 186.365000 72.180000 186.565000 ;
        RECT 71.980000 186.770000 72.180000 186.970000 ;
        RECT 71.980000 187.175000 72.180000 187.375000 ;
        RECT 71.980000 187.580000 72.180000 187.780000 ;
        RECT 71.980000 187.985000 72.180000 188.185000 ;
        RECT 71.980000 188.390000 72.180000 188.590000 ;
        RECT 71.980000 188.795000 72.180000 188.995000 ;
        RECT 71.980000 189.200000 72.180000 189.400000 ;
        RECT 71.980000 189.605000 72.180000 189.805000 ;
        RECT 71.980000 190.010000 72.180000 190.210000 ;
        RECT 71.980000 190.415000 72.180000 190.615000 ;
        RECT 71.980000 190.820000 72.180000 191.020000 ;
        RECT 71.980000 191.225000 72.180000 191.425000 ;
        RECT 71.980000 191.630000 72.180000 191.830000 ;
        RECT 71.980000 192.035000 72.180000 192.235000 ;
        RECT 71.980000 192.440000 72.180000 192.640000 ;
        RECT 71.980000 192.845000 72.180000 193.045000 ;
        RECT 71.980000 193.250000 72.180000 193.450000 ;
        RECT 71.980000 193.655000 72.180000 193.855000 ;
        RECT 71.980000 194.060000 72.180000 194.260000 ;
        RECT 71.980000 194.465000 72.180000 194.665000 ;
        RECT 71.980000 194.870000 72.180000 195.070000 ;
        RECT 71.980000 195.275000 72.180000 195.475000 ;
        RECT 71.980000 195.680000 72.180000 195.880000 ;
        RECT 71.980000 196.085000 72.180000 196.285000 ;
        RECT 71.980000 196.490000 72.180000 196.690000 ;
        RECT 71.980000 196.895000 72.180000 197.095000 ;
        RECT 71.980000 197.300000 72.180000 197.500000 ;
        RECT 71.980000 197.705000 72.180000 197.905000 ;
        RECT 72.380000  23.910000 72.580000  24.110000 ;
        RECT 72.380000  24.340000 72.580000  24.540000 ;
        RECT 72.380000  24.770000 72.580000  24.970000 ;
        RECT 72.380000  25.200000 72.580000  25.400000 ;
        RECT 72.380000  25.630000 72.580000  25.830000 ;
        RECT 72.380000  26.060000 72.580000  26.260000 ;
        RECT 72.380000  26.490000 72.580000  26.690000 ;
        RECT 72.380000  26.920000 72.580000  27.120000 ;
        RECT 72.380000  27.350000 72.580000  27.550000 ;
        RECT 72.380000  27.780000 72.580000  27.980000 ;
        RECT 72.380000  28.210000 72.580000  28.410000 ;
        RECT 72.390000 173.900000 72.590000 174.100000 ;
        RECT 72.390000 174.300000 72.590000 174.500000 ;
        RECT 72.390000 174.700000 72.590000 174.900000 ;
        RECT 72.390000 175.100000 72.590000 175.300000 ;
        RECT 72.390000 175.500000 72.590000 175.700000 ;
        RECT 72.390000 175.900000 72.590000 176.100000 ;
        RECT 72.390000 176.300000 72.590000 176.500000 ;
        RECT 72.390000 176.700000 72.590000 176.900000 ;
        RECT 72.390000 177.100000 72.590000 177.300000 ;
        RECT 72.390000 177.500000 72.590000 177.700000 ;
        RECT 72.390000 177.900000 72.590000 178.100000 ;
        RECT 72.390000 178.300000 72.590000 178.500000 ;
        RECT 72.390000 178.700000 72.590000 178.900000 ;
        RECT 72.390000 179.100000 72.590000 179.300000 ;
        RECT 72.390000 179.500000 72.590000 179.700000 ;
        RECT 72.390000 179.900000 72.590000 180.100000 ;
        RECT 72.390000 180.300000 72.590000 180.500000 ;
        RECT 72.390000 180.700000 72.590000 180.900000 ;
        RECT 72.390000 181.100000 72.590000 181.300000 ;
        RECT 72.390000 181.505000 72.590000 181.705000 ;
        RECT 72.390000 181.910000 72.590000 182.110000 ;
        RECT 72.390000 182.315000 72.590000 182.515000 ;
        RECT 72.390000 182.720000 72.590000 182.920000 ;
        RECT 72.390000 183.125000 72.590000 183.325000 ;
        RECT 72.390000 183.530000 72.590000 183.730000 ;
        RECT 72.390000 183.935000 72.590000 184.135000 ;
        RECT 72.390000 184.340000 72.590000 184.540000 ;
        RECT 72.390000 184.745000 72.590000 184.945000 ;
        RECT 72.390000 185.150000 72.590000 185.350000 ;
        RECT 72.390000 185.555000 72.590000 185.755000 ;
        RECT 72.390000 185.960000 72.590000 186.160000 ;
        RECT 72.390000 186.365000 72.590000 186.565000 ;
        RECT 72.390000 186.770000 72.590000 186.970000 ;
        RECT 72.390000 187.175000 72.590000 187.375000 ;
        RECT 72.390000 187.580000 72.590000 187.780000 ;
        RECT 72.390000 187.985000 72.590000 188.185000 ;
        RECT 72.390000 188.390000 72.590000 188.590000 ;
        RECT 72.390000 188.795000 72.590000 188.995000 ;
        RECT 72.390000 189.200000 72.590000 189.400000 ;
        RECT 72.390000 189.605000 72.590000 189.805000 ;
        RECT 72.390000 190.010000 72.590000 190.210000 ;
        RECT 72.390000 190.415000 72.590000 190.615000 ;
        RECT 72.390000 190.820000 72.590000 191.020000 ;
        RECT 72.390000 191.225000 72.590000 191.425000 ;
        RECT 72.390000 191.630000 72.590000 191.830000 ;
        RECT 72.390000 192.035000 72.590000 192.235000 ;
        RECT 72.390000 192.440000 72.590000 192.640000 ;
        RECT 72.390000 192.845000 72.590000 193.045000 ;
        RECT 72.390000 193.250000 72.590000 193.450000 ;
        RECT 72.390000 193.655000 72.590000 193.855000 ;
        RECT 72.390000 194.060000 72.590000 194.260000 ;
        RECT 72.390000 194.465000 72.590000 194.665000 ;
        RECT 72.390000 194.870000 72.590000 195.070000 ;
        RECT 72.390000 195.275000 72.590000 195.475000 ;
        RECT 72.390000 195.680000 72.590000 195.880000 ;
        RECT 72.390000 196.085000 72.590000 196.285000 ;
        RECT 72.390000 196.490000 72.590000 196.690000 ;
        RECT 72.390000 196.895000 72.590000 197.095000 ;
        RECT 72.390000 197.300000 72.590000 197.500000 ;
        RECT 72.390000 197.705000 72.590000 197.905000 ;
        RECT 72.785000  23.910000 72.985000  24.110000 ;
        RECT 72.785000  24.340000 72.985000  24.540000 ;
        RECT 72.785000  24.770000 72.985000  24.970000 ;
        RECT 72.785000  25.200000 72.985000  25.400000 ;
        RECT 72.785000  25.630000 72.985000  25.830000 ;
        RECT 72.785000  26.060000 72.985000  26.260000 ;
        RECT 72.785000  26.490000 72.985000  26.690000 ;
        RECT 72.785000  26.920000 72.985000  27.120000 ;
        RECT 72.785000  27.350000 72.985000  27.550000 ;
        RECT 72.785000  27.780000 72.985000  27.980000 ;
        RECT 72.785000  28.210000 72.985000  28.410000 ;
        RECT 72.800000 173.900000 73.000000 174.100000 ;
        RECT 72.800000 174.300000 73.000000 174.500000 ;
        RECT 72.800000 174.700000 73.000000 174.900000 ;
        RECT 72.800000 175.100000 73.000000 175.300000 ;
        RECT 72.800000 175.500000 73.000000 175.700000 ;
        RECT 72.800000 175.900000 73.000000 176.100000 ;
        RECT 72.800000 176.300000 73.000000 176.500000 ;
        RECT 72.800000 176.700000 73.000000 176.900000 ;
        RECT 72.800000 177.100000 73.000000 177.300000 ;
        RECT 72.800000 177.500000 73.000000 177.700000 ;
        RECT 72.800000 177.900000 73.000000 178.100000 ;
        RECT 72.800000 178.300000 73.000000 178.500000 ;
        RECT 72.800000 178.700000 73.000000 178.900000 ;
        RECT 72.800000 179.100000 73.000000 179.300000 ;
        RECT 72.800000 179.500000 73.000000 179.700000 ;
        RECT 72.800000 179.900000 73.000000 180.100000 ;
        RECT 72.800000 180.300000 73.000000 180.500000 ;
        RECT 72.800000 180.700000 73.000000 180.900000 ;
        RECT 72.800000 181.100000 73.000000 181.300000 ;
        RECT 72.800000 181.505000 73.000000 181.705000 ;
        RECT 72.800000 181.910000 73.000000 182.110000 ;
        RECT 72.800000 182.315000 73.000000 182.515000 ;
        RECT 72.800000 182.720000 73.000000 182.920000 ;
        RECT 72.800000 183.125000 73.000000 183.325000 ;
        RECT 72.800000 183.530000 73.000000 183.730000 ;
        RECT 72.800000 183.935000 73.000000 184.135000 ;
        RECT 72.800000 184.340000 73.000000 184.540000 ;
        RECT 72.800000 184.745000 73.000000 184.945000 ;
        RECT 72.800000 185.150000 73.000000 185.350000 ;
        RECT 72.800000 185.555000 73.000000 185.755000 ;
        RECT 72.800000 185.960000 73.000000 186.160000 ;
        RECT 72.800000 186.365000 73.000000 186.565000 ;
        RECT 72.800000 186.770000 73.000000 186.970000 ;
        RECT 72.800000 187.175000 73.000000 187.375000 ;
        RECT 72.800000 187.580000 73.000000 187.780000 ;
        RECT 72.800000 187.985000 73.000000 188.185000 ;
        RECT 72.800000 188.390000 73.000000 188.590000 ;
        RECT 72.800000 188.795000 73.000000 188.995000 ;
        RECT 72.800000 189.200000 73.000000 189.400000 ;
        RECT 72.800000 189.605000 73.000000 189.805000 ;
        RECT 72.800000 190.010000 73.000000 190.210000 ;
        RECT 72.800000 190.415000 73.000000 190.615000 ;
        RECT 72.800000 190.820000 73.000000 191.020000 ;
        RECT 72.800000 191.225000 73.000000 191.425000 ;
        RECT 72.800000 191.630000 73.000000 191.830000 ;
        RECT 72.800000 192.035000 73.000000 192.235000 ;
        RECT 72.800000 192.440000 73.000000 192.640000 ;
        RECT 72.800000 192.845000 73.000000 193.045000 ;
        RECT 72.800000 193.250000 73.000000 193.450000 ;
        RECT 72.800000 193.655000 73.000000 193.855000 ;
        RECT 72.800000 194.060000 73.000000 194.260000 ;
        RECT 72.800000 194.465000 73.000000 194.665000 ;
        RECT 72.800000 194.870000 73.000000 195.070000 ;
        RECT 72.800000 195.275000 73.000000 195.475000 ;
        RECT 72.800000 195.680000 73.000000 195.880000 ;
        RECT 72.800000 196.085000 73.000000 196.285000 ;
        RECT 72.800000 196.490000 73.000000 196.690000 ;
        RECT 72.800000 196.895000 73.000000 197.095000 ;
        RECT 72.800000 197.300000 73.000000 197.500000 ;
        RECT 72.800000 197.705000 73.000000 197.905000 ;
        RECT 73.190000  23.910000 73.390000  24.110000 ;
        RECT 73.190000  24.340000 73.390000  24.540000 ;
        RECT 73.190000  24.770000 73.390000  24.970000 ;
        RECT 73.190000  25.200000 73.390000  25.400000 ;
        RECT 73.190000  25.630000 73.390000  25.830000 ;
        RECT 73.190000  26.060000 73.390000  26.260000 ;
        RECT 73.190000  26.490000 73.390000  26.690000 ;
        RECT 73.190000  26.920000 73.390000  27.120000 ;
        RECT 73.190000  27.350000 73.390000  27.550000 ;
        RECT 73.190000  27.780000 73.390000  27.980000 ;
        RECT 73.190000  28.210000 73.390000  28.410000 ;
        RECT 73.210000 173.900000 73.410000 174.100000 ;
        RECT 73.210000 174.300000 73.410000 174.500000 ;
        RECT 73.210000 174.700000 73.410000 174.900000 ;
        RECT 73.210000 175.100000 73.410000 175.300000 ;
        RECT 73.210000 175.500000 73.410000 175.700000 ;
        RECT 73.210000 175.900000 73.410000 176.100000 ;
        RECT 73.210000 176.300000 73.410000 176.500000 ;
        RECT 73.210000 176.700000 73.410000 176.900000 ;
        RECT 73.210000 177.100000 73.410000 177.300000 ;
        RECT 73.210000 177.500000 73.410000 177.700000 ;
        RECT 73.210000 177.900000 73.410000 178.100000 ;
        RECT 73.210000 178.300000 73.410000 178.500000 ;
        RECT 73.210000 178.700000 73.410000 178.900000 ;
        RECT 73.210000 179.100000 73.410000 179.300000 ;
        RECT 73.210000 179.500000 73.410000 179.700000 ;
        RECT 73.210000 179.900000 73.410000 180.100000 ;
        RECT 73.210000 180.300000 73.410000 180.500000 ;
        RECT 73.210000 180.700000 73.410000 180.900000 ;
        RECT 73.210000 181.100000 73.410000 181.300000 ;
        RECT 73.210000 181.505000 73.410000 181.705000 ;
        RECT 73.210000 181.910000 73.410000 182.110000 ;
        RECT 73.210000 182.315000 73.410000 182.515000 ;
        RECT 73.210000 182.720000 73.410000 182.920000 ;
        RECT 73.210000 183.125000 73.410000 183.325000 ;
        RECT 73.210000 183.530000 73.410000 183.730000 ;
        RECT 73.210000 183.935000 73.410000 184.135000 ;
        RECT 73.210000 184.340000 73.410000 184.540000 ;
        RECT 73.210000 184.745000 73.410000 184.945000 ;
        RECT 73.210000 185.150000 73.410000 185.350000 ;
        RECT 73.210000 185.555000 73.410000 185.755000 ;
        RECT 73.210000 185.960000 73.410000 186.160000 ;
        RECT 73.210000 186.365000 73.410000 186.565000 ;
        RECT 73.210000 186.770000 73.410000 186.970000 ;
        RECT 73.210000 187.175000 73.410000 187.375000 ;
        RECT 73.210000 187.580000 73.410000 187.780000 ;
        RECT 73.210000 187.985000 73.410000 188.185000 ;
        RECT 73.210000 188.390000 73.410000 188.590000 ;
        RECT 73.210000 188.795000 73.410000 188.995000 ;
        RECT 73.210000 189.200000 73.410000 189.400000 ;
        RECT 73.210000 189.605000 73.410000 189.805000 ;
        RECT 73.210000 190.010000 73.410000 190.210000 ;
        RECT 73.210000 190.415000 73.410000 190.615000 ;
        RECT 73.210000 190.820000 73.410000 191.020000 ;
        RECT 73.210000 191.225000 73.410000 191.425000 ;
        RECT 73.210000 191.630000 73.410000 191.830000 ;
        RECT 73.210000 192.035000 73.410000 192.235000 ;
        RECT 73.210000 192.440000 73.410000 192.640000 ;
        RECT 73.210000 192.845000 73.410000 193.045000 ;
        RECT 73.210000 193.250000 73.410000 193.450000 ;
        RECT 73.210000 193.655000 73.410000 193.855000 ;
        RECT 73.210000 194.060000 73.410000 194.260000 ;
        RECT 73.210000 194.465000 73.410000 194.665000 ;
        RECT 73.210000 194.870000 73.410000 195.070000 ;
        RECT 73.210000 195.275000 73.410000 195.475000 ;
        RECT 73.210000 195.680000 73.410000 195.880000 ;
        RECT 73.210000 196.085000 73.410000 196.285000 ;
        RECT 73.210000 196.490000 73.410000 196.690000 ;
        RECT 73.210000 196.895000 73.410000 197.095000 ;
        RECT 73.210000 197.300000 73.410000 197.500000 ;
        RECT 73.210000 197.705000 73.410000 197.905000 ;
        RECT 73.595000  23.910000 73.795000  24.110000 ;
        RECT 73.595000  24.340000 73.795000  24.540000 ;
        RECT 73.595000  24.770000 73.795000  24.970000 ;
        RECT 73.595000  25.200000 73.795000  25.400000 ;
        RECT 73.595000  25.630000 73.795000  25.830000 ;
        RECT 73.595000  26.060000 73.795000  26.260000 ;
        RECT 73.595000  26.490000 73.795000  26.690000 ;
        RECT 73.595000  26.920000 73.795000  27.120000 ;
        RECT 73.595000  27.350000 73.795000  27.550000 ;
        RECT 73.595000  27.780000 73.795000  27.980000 ;
        RECT 73.595000  28.210000 73.795000  28.410000 ;
        RECT 73.620000 173.900000 73.820000 174.100000 ;
        RECT 73.620000 174.300000 73.820000 174.500000 ;
        RECT 73.620000 174.700000 73.820000 174.900000 ;
        RECT 73.620000 175.100000 73.820000 175.300000 ;
        RECT 73.620000 175.500000 73.820000 175.700000 ;
        RECT 73.620000 175.900000 73.820000 176.100000 ;
        RECT 73.620000 176.300000 73.820000 176.500000 ;
        RECT 73.620000 176.700000 73.820000 176.900000 ;
        RECT 73.620000 177.100000 73.820000 177.300000 ;
        RECT 73.620000 177.500000 73.820000 177.700000 ;
        RECT 73.620000 177.900000 73.820000 178.100000 ;
        RECT 73.620000 178.300000 73.820000 178.500000 ;
        RECT 73.620000 178.700000 73.820000 178.900000 ;
        RECT 73.620000 179.100000 73.820000 179.300000 ;
        RECT 73.620000 179.500000 73.820000 179.700000 ;
        RECT 73.620000 179.900000 73.820000 180.100000 ;
        RECT 73.620000 180.300000 73.820000 180.500000 ;
        RECT 73.620000 180.700000 73.820000 180.900000 ;
        RECT 73.620000 181.100000 73.820000 181.300000 ;
        RECT 73.620000 181.505000 73.820000 181.705000 ;
        RECT 73.620000 181.910000 73.820000 182.110000 ;
        RECT 73.620000 182.315000 73.820000 182.515000 ;
        RECT 73.620000 182.720000 73.820000 182.920000 ;
        RECT 73.620000 183.125000 73.820000 183.325000 ;
        RECT 73.620000 183.530000 73.820000 183.730000 ;
        RECT 73.620000 183.935000 73.820000 184.135000 ;
        RECT 73.620000 184.340000 73.820000 184.540000 ;
        RECT 73.620000 184.745000 73.820000 184.945000 ;
        RECT 73.620000 185.150000 73.820000 185.350000 ;
        RECT 73.620000 185.555000 73.820000 185.755000 ;
        RECT 73.620000 185.960000 73.820000 186.160000 ;
        RECT 73.620000 186.365000 73.820000 186.565000 ;
        RECT 73.620000 186.770000 73.820000 186.970000 ;
        RECT 73.620000 187.175000 73.820000 187.375000 ;
        RECT 73.620000 187.580000 73.820000 187.780000 ;
        RECT 73.620000 187.985000 73.820000 188.185000 ;
        RECT 73.620000 188.390000 73.820000 188.590000 ;
        RECT 73.620000 188.795000 73.820000 188.995000 ;
        RECT 73.620000 189.200000 73.820000 189.400000 ;
        RECT 73.620000 189.605000 73.820000 189.805000 ;
        RECT 73.620000 190.010000 73.820000 190.210000 ;
        RECT 73.620000 190.415000 73.820000 190.615000 ;
        RECT 73.620000 190.820000 73.820000 191.020000 ;
        RECT 73.620000 191.225000 73.820000 191.425000 ;
        RECT 73.620000 191.630000 73.820000 191.830000 ;
        RECT 73.620000 192.035000 73.820000 192.235000 ;
        RECT 73.620000 192.440000 73.820000 192.640000 ;
        RECT 73.620000 192.845000 73.820000 193.045000 ;
        RECT 73.620000 193.250000 73.820000 193.450000 ;
        RECT 73.620000 193.655000 73.820000 193.855000 ;
        RECT 73.620000 194.060000 73.820000 194.260000 ;
        RECT 73.620000 194.465000 73.820000 194.665000 ;
        RECT 73.620000 194.870000 73.820000 195.070000 ;
        RECT 73.620000 195.275000 73.820000 195.475000 ;
        RECT 73.620000 195.680000 73.820000 195.880000 ;
        RECT 73.620000 196.085000 73.820000 196.285000 ;
        RECT 73.620000 196.490000 73.820000 196.690000 ;
        RECT 73.620000 196.895000 73.820000 197.095000 ;
        RECT 73.620000 197.300000 73.820000 197.500000 ;
        RECT 73.620000 197.705000 73.820000 197.905000 ;
        RECT 74.000000  23.910000 74.200000  24.110000 ;
        RECT 74.000000  24.340000 74.200000  24.540000 ;
        RECT 74.000000  24.770000 74.200000  24.970000 ;
        RECT 74.000000  25.200000 74.200000  25.400000 ;
        RECT 74.000000  25.630000 74.200000  25.830000 ;
        RECT 74.000000  26.060000 74.200000  26.260000 ;
        RECT 74.000000  26.490000 74.200000  26.690000 ;
        RECT 74.000000  26.920000 74.200000  27.120000 ;
        RECT 74.000000  27.350000 74.200000  27.550000 ;
        RECT 74.000000  27.780000 74.200000  27.980000 ;
        RECT 74.000000  28.210000 74.200000  28.410000 ;
        RECT 74.030000 173.900000 74.230000 174.100000 ;
        RECT 74.030000 174.300000 74.230000 174.500000 ;
        RECT 74.030000 174.700000 74.230000 174.900000 ;
        RECT 74.030000 175.100000 74.230000 175.300000 ;
        RECT 74.030000 175.500000 74.230000 175.700000 ;
        RECT 74.030000 175.900000 74.230000 176.100000 ;
        RECT 74.030000 176.300000 74.230000 176.500000 ;
        RECT 74.030000 176.700000 74.230000 176.900000 ;
        RECT 74.030000 177.100000 74.230000 177.300000 ;
        RECT 74.030000 177.500000 74.230000 177.700000 ;
        RECT 74.030000 177.900000 74.230000 178.100000 ;
        RECT 74.030000 178.300000 74.230000 178.500000 ;
        RECT 74.030000 178.700000 74.230000 178.900000 ;
        RECT 74.030000 179.100000 74.230000 179.300000 ;
        RECT 74.030000 179.500000 74.230000 179.700000 ;
        RECT 74.030000 179.900000 74.230000 180.100000 ;
        RECT 74.030000 180.300000 74.230000 180.500000 ;
        RECT 74.030000 180.700000 74.230000 180.900000 ;
        RECT 74.030000 181.100000 74.230000 181.300000 ;
        RECT 74.030000 181.505000 74.230000 181.705000 ;
        RECT 74.030000 181.910000 74.230000 182.110000 ;
        RECT 74.030000 182.315000 74.230000 182.515000 ;
        RECT 74.030000 182.720000 74.230000 182.920000 ;
        RECT 74.030000 183.125000 74.230000 183.325000 ;
        RECT 74.030000 183.530000 74.230000 183.730000 ;
        RECT 74.030000 183.935000 74.230000 184.135000 ;
        RECT 74.030000 184.340000 74.230000 184.540000 ;
        RECT 74.030000 184.745000 74.230000 184.945000 ;
        RECT 74.030000 185.150000 74.230000 185.350000 ;
        RECT 74.030000 185.555000 74.230000 185.755000 ;
        RECT 74.030000 185.960000 74.230000 186.160000 ;
        RECT 74.030000 186.365000 74.230000 186.565000 ;
        RECT 74.030000 186.770000 74.230000 186.970000 ;
        RECT 74.030000 187.175000 74.230000 187.375000 ;
        RECT 74.030000 187.580000 74.230000 187.780000 ;
        RECT 74.030000 187.985000 74.230000 188.185000 ;
        RECT 74.030000 188.390000 74.230000 188.590000 ;
        RECT 74.030000 188.795000 74.230000 188.995000 ;
        RECT 74.030000 189.200000 74.230000 189.400000 ;
        RECT 74.030000 189.605000 74.230000 189.805000 ;
        RECT 74.030000 190.010000 74.230000 190.210000 ;
        RECT 74.030000 190.415000 74.230000 190.615000 ;
        RECT 74.030000 190.820000 74.230000 191.020000 ;
        RECT 74.030000 191.225000 74.230000 191.425000 ;
        RECT 74.030000 191.630000 74.230000 191.830000 ;
        RECT 74.030000 192.035000 74.230000 192.235000 ;
        RECT 74.030000 192.440000 74.230000 192.640000 ;
        RECT 74.030000 192.845000 74.230000 193.045000 ;
        RECT 74.030000 193.250000 74.230000 193.450000 ;
        RECT 74.030000 193.655000 74.230000 193.855000 ;
        RECT 74.030000 194.060000 74.230000 194.260000 ;
        RECT 74.030000 194.465000 74.230000 194.665000 ;
        RECT 74.030000 194.870000 74.230000 195.070000 ;
        RECT 74.030000 195.275000 74.230000 195.475000 ;
        RECT 74.030000 195.680000 74.230000 195.880000 ;
        RECT 74.030000 196.085000 74.230000 196.285000 ;
        RECT 74.030000 196.490000 74.230000 196.690000 ;
        RECT 74.030000 196.895000 74.230000 197.095000 ;
        RECT 74.030000 197.300000 74.230000 197.500000 ;
        RECT 74.030000 197.705000 74.230000 197.905000 ;
        RECT 74.440000 173.900000 74.640000 174.100000 ;
        RECT 74.440000 174.300000 74.640000 174.500000 ;
        RECT 74.440000 174.700000 74.640000 174.900000 ;
        RECT 74.440000 175.100000 74.640000 175.300000 ;
        RECT 74.440000 175.500000 74.640000 175.700000 ;
        RECT 74.440000 175.900000 74.640000 176.100000 ;
        RECT 74.440000 176.300000 74.640000 176.500000 ;
        RECT 74.440000 176.700000 74.640000 176.900000 ;
        RECT 74.440000 177.100000 74.640000 177.300000 ;
        RECT 74.440000 177.500000 74.640000 177.700000 ;
        RECT 74.440000 177.900000 74.640000 178.100000 ;
        RECT 74.440000 178.300000 74.640000 178.500000 ;
        RECT 74.440000 178.700000 74.640000 178.900000 ;
        RECT 74.440000 179.100000 74.640000 179.300000 ;
        RECT 74.440000 179.500000 74.640000 179.700000 ;
        RECT 74.440000 179.900000 74.640000 180.100000 ;
        RECT 74.440000 180.300000 74.640000 180.500000 ;
        RECT 74.440000 180.700000 74.640000 180.900000 ;
        RECT 74.440000 181.100000 74.640000 181.300000 ;
        RECT 74.440000 181.505000 74.640000 181.705000 ;
        RECT 74.440000 181.910000 74.640000 182.110000 ;
        RECT 74.440000 182.315000 74.640000 182.515000 ;
        RECT 74.440000 182.720000 74.640000 182.920000 ;
        RECT 74.440000 183.125000 74.640000 183.325000 ;
        RECT 74.440000 183.530000 74.640000 183.730000 ;
        RECT 74.440000 183.935000 74.640000 184.135000 ;
        RECT 74.440000 184.340000 74.640000 184.540000 ;
        RECT 74.440000 184.745000 74.640000 184.945000 ;
        RECT 74.440000 185.150000 74.640000 185.350000 ;
        RECT 74.440000 185.555000 74.640000 185.755000 ;
        RECT 74.440000 185.960000 74.640000 186.160000 ;
        RECT 74.440000 186.365000 74.640000 186.565000 ;
        RECT 74.440000 186.770000 74.640000 186.970000 ;
        RECT 74.440000 187.175000 74.640000 187.375000 ;
        RECT 74.440000 187.580000 74.640000 187.780000 ;
        RECT 74.440000 187.985000 74.640000 188.185000 ;
        RECT 74.440000 188.390000 74.640000 188.590000 ;
        RECT 74.440000 188.795000 74.640000 188.995000 ;
        RECT 74.440000 189.200000 74.640000 189.400000 ;
        RECT 74.440000 189.605000 74.640000 189.805000 ;
        RECT 74.440000 190.010000 74.640000 190.210000 ;
        RECT 74.440000 190.415000 74.640000 190.615000 ;
        RECT 74.440000 190.820000 74.640000 191.020000 ;
        RECT 74.440000 191.225000 74.640000 191.425000 ;
        RECT 74.440000 191.630000 74.640000 191.830000 ;
        RECT 74.440000 192.035000 74.640000 192.235000 ;
        RECT 74.440000 192.440000 74.640000 192.640000 ;
        RECT 74.440000 192.845000 74.640000 193.045000 ;
        RECT 74.440000 193.250000 74.640000 193.450000 ;
        RECT 74.440000 193.655000 74.640000 193.855000 ;
        RECT 74.440000 194.060000 74.640000 194.260000 ;
        RECT 74.440000 194.465000 74.640000 194.665000 ;
        RECT 74.440000 194.870000 74.640000 195.070000 ;
        RECT 74.440000 195.275000 74.640000 195.475000 ;
        RECT 74.440000 195.680000 74.640000 195.880000 ;
        RECT 74.440000 196.085000 74.640000 196.285000 ;
        RECT 74.440000 196.490000 74.640000 196.690000 ;
        RECT 74.440000 196.895000 74.640000 197.095000 ;
        RECT 74.440000 197.300000 74.640000 197.500000 ;
        RECT 74.440000 197.705000 74.640000 197.905000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.500000 56.240000 24.400000 60.680000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 56.240000 74.290000 60.680000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 24.375000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.590000 56.310000  0.790000 56.510000 ;
        RECT  0.590000 56.720000  0.790000 56.920000 ;
        RECT  0.590000 57.130000  0.790000 57.330000 ;
        RECT  0.590000 57.540000  0.790000 57.740000 ;
        RECT  0.590000 57.950000  0.790000 58.150000 ;
        RECT  0.590000 58.360000  0.790000 58.560000 ;
        RECT  0.590000 58.770000  0.790000 58.970000 ;
        RECT  0.590000 59.180000  0.790000 59.380000 ;
        RECT  0.590000 59.590000  0.790000 59.790000 ;
        RECT  0.590000 60.000000  0.790000 60.200000 ;
        RECT  0.590000 60.410000  0.790000 60.610000 ;
        RECT  1.000000 56.310000  1.200000 56.510000 ;
        RECT  1.000000 56.720000  1.200000 56.920000 ;
        RECT  1.000000 57.130000  1.200000 57.330000 ;
        RECT  1.000000 57.540000  1.200000 57.740000 ;
        RECT  1.000000 57.950000  1.200000 58.150000 ;
        RECT  1.000000 58.360000  1.200000 58.560000 ;
        RECT  1.000000 58.770000  1.200000 58.970000 ;
        RECT  1.000000 59.180000  1.200000 59.380000 ;
        RECT  1.000000 59.590000  1.200000 59.790000 ;
        RECT  1.000000 60.000000  1.200000 60.200000 ;
        RECT  1.000000 60.410000  1.200000 60.610000 ;
        RECT  1.410000 56.310000  1.610000 56.510000 ;
        RECT  1.410000 56.720000  1.610000 56.920000 ;
        RECT  1.410000 57.130000  1.610000 57.330000 ;
        RECT  1.410000 57.540000  1.610000 57.740000 ;
        RECT  1.410000 57.950000  1.610000 58.150000 ;
        RECT  1.410000 58.360000  1.610000 58.560000 ;
        RECT  1.410000 58.770000  1.610000 58.970000 ;
        RECT  1.410000 59.180000  1.610000 59.380000 ;
        RECT  1.410000 59.590000  1.610000 59.790000 ;
        RECT  1.410000 60.000000  1.610000 60.200000 ;
        RECT  1.410000 60.410000  1.610000 60.610000 ;
        RECT  1.820000 56.310000  2.020000 56.510000 ;
        RECT  1.820000 56.720000  2.020000 56.920000 ;
        RECT  1.820000 57.130000  2.020000 57.330000 ;
        RECT  1.820000 57.540000  2.020000 57.740000 ;
        RECT  1.820000 57.950000  2.020000 58.150000 ;
        RECT  1.820000 58.360000  2.020000 58.560000 ;
        RECT  1.820000 58.770000  2.020000 58.970000 ;
        RECT  1.820000 59.180000  2.020000 59.380000 ;
        RECT  1.820000 59.590000  2.020000 59.790000 ;
        RECT  1.820000 60.000000  2.020000 60.200000 ;
        RECT  1.820000 60.410000  2.020000 60.610000 ;
        RECT  2.230000 56.310000  2.430000 56.510000 ;
        RECT  2.230000 56.720000  2.430000 56.920000 ;
        RECT  2.230000 57.130000  2.430000 57.330000 ;
        RECT  2.230000 57.540000  2.430000 57.740000 ;
        RECT  2.230000 57.950000  2.430000 58.150000 ;
        RECT  2.230000 58.360000  2.430000 58.560000 ;
        RECT  2.230000 58.770000  2.430000 58.970000 ;
        RECT  2.230000 59.180000  2.430000 59.380000 ;
        RECT  2.230000 59.590000  2.430000 59.790000 ;
        RECT  2.230000 60.000000  2.430000 60.200000 ;
        RECT  2.230000 60.410000  2.430000 60.610000 ;
        RECT  2.640000 56.310000  2.840000 56.510000 ;
        RECT  2.640000 56.720000  2.840000 56.920000 ;
        RECT  2.640000 57.130000  2.840000 57.330000 ;
        RECT  2.640000 57.540000  2.840000 57.740000 ;
        RECT  2.640000 57.950000  2.840000 58.150000 ;
        RECT  2.640000 58.360000  2.840000 58.560000 ;
        RECT  2.640000 58.770000  2.840000 58.970000 ;
        RECT  2.640000 59.180000  2.840000 59.380000 ;
        RECT  2.640000 59.590000  2.840000 59.790000 ;
        RECT  2.640000 60.000000  2.840000 60.200000 ;
        RECT  2.640000 60.410000  2.840000 60.610000 ;
        RECT  3.050000 56.310000  3.250000 56.510000 ;
        RECT  3.050000 56.720000  3.250000 56.920000 ;
        RECT  3.050000 57.130000  3.250000 57.330000 ;
        RECT  3.050000 57.540000  3.250000 57.740000 ;
        RECT  3.050000 57.950000  3.250000 58.150000 ;
        RECT  3.050000 58.360000  3.250000 58.560000 ;
        RECT  3.050000 58.770000  3.250000 58.970000 ;
        RECT  3.050000 59.180000  3.250000 59.380000 ;
        RECT  3.050000 59.590000  3.250000 59.790000 ;
        RECT  3.050000 60.000000  3.250000 60.200000 ;
        RECT  3.050000 60.410000  3.250000 60.610000 ;
        RECT  3.455000 56.310000  3.655000 56.510000 ;
        RECT  3.455000 56.720000  3.655000 56.920000 ;
        RECT  3.455000 57.130000  3.655000 57.330000 ;
        RECT  3.455000 57.540000  3.655000 57.740000 ;
        RECT  3.455000 57.950000  3.655000 58.150000 ;
        RECT  3.455000 58.360000  3.655000 58.560000 ;
        RECT  3.455000 58.770000  3.655000 58.970000 ;
        RECT  3.455000 59.180000  3.655000 59.380000 ;
        RECT  3.455000 59.590000  3.655000 59.790000 ;
        RECT  3.455000 60.000000  3.655000 60.200000 ;
        RECT  3.455000 60.410000  3.655000 60.610000 ;
        RECT  3.860000 56.310000  4.060000 56.510000 ;
        RECT  3.860000 56.720000  4.060000 56.920000 ;
        RECT  3.860000 57.130000  4.060000 57.330000 ;
        RECT  3.860000 57.540000  4.060000 57.740000 ;
        RECT  3.860000 57.950000  4.060000 58.150000 ;
        RECT  3.860000 58.360000  4.060000 58.560000 ;
        RECT  3.860000 58.770000  4.060000 58.970000 ;
        RECT  3.860000 59.180000  4.060000 59.380000 ;
        RECT  3.860000 59.590000  4.060000 59.790000 ;
        RECT  3.860000 60.000000  4.060000 60.200000 ;
        RECT  3.860000 60.410000  4.060000 60.610000 ;
        RECT  4.265000 56.310000  4.465000 56.510000 ;
        RECT  4.265000 56.720000  4.465000 56.920000 ;
        RECT  4.265000 57.130000  4.465000 57.330000 ;
        RECT  4.265000 57.540000  4.465000 57.740000 ;
        RECT  4.265000 57.950000  4.465000 58.150000 ;
        RECT  4.265000 58.360000  4.465000 58.560000 ;
        RECT  4.265000 58.770000  4.465000 58.970000 ;
        RECT  4.265000 59.180000  4.465000 59.380000 ;
        RECT  4.265000 59.590000  4.465000 59.790000 ;
        RECT  4.265000 60.000000  4.465000 60.200000 ;
        RECT  4.265000 60.410000  4.465000 60.610000 ;
        RECT  4.670000 56.310000  4.870000 56.510000 ;
        RECT  4.670000 56.720000  4.870000 56.920000 ;
        RECT  4.670000 57.130000  4.870000 57.330000 ;
        RECT  4.670000 57.540000  4.870000 57.740000 ;
        RECT  4.670000 57.950000  4.870000 58.150000 ;
        RECT  4.670000 58.360000  4.870000 58.560000 ;
        RECT  4.670000 58.770000  4.870000 58.970000 ;
        RECT  4.670000 59.180000  4.870000 59.380000 ;
        RECT  4.670000 59.590000  4.870000 59.790000 ;
        RECT  4.670000 60.000000  4.870000 60.200000 ;
        RECT  4.670000 60.410000  4.870000 60.610000 ;
        RECT  5.075000 56.310000  5.275000 56.510000 ;
        RECT  5.075000 56.720000  5.275000 56.920000 ;
        RECT  5.075000 57.130000  5.275000 57.330000 ;
        RECT  5.075000 57.540000  5.275000 57.740000 ;
        RECT  5.075000 57.950000  5.275000 58.150000 ;
        RECT  5.075000 58.360000  5.275000 58.560000 ;
        RECT  5.075000 58.770000  5.275000 58.970000 ;
        RECT  5.075000 59.180000  5.275000 59.380000 ;
        RECT  5.075000 59.590000  5.275000 59.790000 ;
        RECT  5.075000 60.000000  5.275000 60.200000 ;
        RECT  5.075000 60.410000  5.275000 60.610000 ;
        RECT  5.480000 56.310000  5.680000 56.510000 ;
        RECT  5.480000 56.720000  5.680000 56.920000 ;
        RECT  5.480000 57.130000  5.680000 57.330000 ;
        RECT  5.480000 57.540000  5.680000 57.740000 ;
        RECT  5.480000 57.950000  5.680000 58.150000 ;
        RECT  5.480000 58.360000  5.680000 58.560000 ;
        RECT  5.480000 58.770000  5.680000 58.970000 ;
        RECT  5.480000 59.180000  5.680000 59.380000 ;
        RECT  5.480000 59.590000  5.680000 59.790000 ;
        RECT  5.480000 60.000000  5.680000 60.200000 ;
        RECT  5.480000 60.410000  5.680000 60.610000 ;
        RECT  5.885000 56.310000  6.085000 56.510000 ;
        RECT  5.885000 56.720000  6.085000 56.920000 ;
        RECT  5.885000 57.130000  6.085000 57.330000 ;
        RECT  5.885000 57.540000  6.085000 57.740000 ;
        RECT  5.885000 57.950000  6.085000 58.150000 ;
        RECT  5.885000 58.360000  6.085000 58.560000 ;
        RECT  5.885000 58.770000  6.085000 58.970000 ;
        RECT  5.885000 59.180000  6.085000 59.380000 ;
        RECT  5.885000 59.590000  6.085000 59.790000 ;
        RECT  5.885000 60.000000  6.085000 60.200000 ;
        RECT  5.885000 60.410000  6.085000 60.610000 ;
        RECT  6.290000 56.310000  6.490000 56.510000 ;
        RECT  6.290000 56.720000  6.490000 56.920000 ;
        RECT  6.290000 57.130000  6.490000 57.330000 ;
        RECT  6.290000 57.540000  6.490000 57.740000 ;
        RECT  6.290000 57.950000  6.490000 58.150000 ;
        RECT  6.290000 58.360000  6.490000 58.560000 ;
        RECT  6.290000 58.770000  6.490000 58.970000 ;
        RECT  6.290000 59.180000  6.490000 59.380000 ;
        RECT  6.290000 59.590000  6.490000 59.790000 ;
        RECT  6.290000 60.000000  6.490000 60.200000 ;
        RECT  6.290000 60.410000  6.490000 60.610000 ;
        RECT  6.695000 56.310000  6.895000 56.510000 ;
        RECT  6.695000 56.720000  6.895000 56.920000 ;
        RECT  6.695000 57.130000  6.895000 57.330000 ;
        RECT  6.695000 57.540000  6.895000 57.740000 ;
        RECT  6.695000 57.950000  6.895000 58.150000 ;
        RECT  6.695000 58.360000  6.895000 58.560000 ;
        RECT  6.695000 58.770000  6.895000 58.970000 ;
        RECT  6.695000 59.180000  6.895000 59.380000 ;
        RECT  6.695000 59.590000  6.895000 59.790000 ;
        RECT  6.695000 60.000000  6.895000 60.200000 ;
        RECT  6.695000 60.410000  6.895000 60.610000 ;
        RECT  7.100000 56.310000  7.300000 56.510000 ;
        RECT  7.100000 56.720000  7.300000 56.920000 ;
        RECT  7.100000 57.130000  7.300000 57.330000 ;
        RECT  7.100000 57.540000  7.300000 57.740000 ;
        RECT  7.100000 57.950000  7.300000 58.150000 ;
        RECT  7.100000 58.360000  7.300000 58.560000 ;
        RECT  7.100000 58.770000  7.300000 58.970000 ;
        RECT  7.100000 59.180000  7.300000 59.380000 ;
        RECT  7.100000 59.590000  7.300000 59.790000 ;
        RECT  7.100000 60.000000  7.300000 60.200000 ;
        RECT  7.100000 60.410000  7.300000 60.610000 ;
        RECT  7.505000 56.310000  7.705000 56.510000 ;
        RECT  7.505000 56.720000  7.705000 56.920000 ;
        RECT  7.505000 57.130000  7.705000 57.330000 ;
        RECT  7.505000 57.540000  7.705000 57.740000 ;
        RECT  7.505000 57.950000  7.705000 58.150000 ;
        RECT  7.505000 58.360000  7.705000 58.560000 ;
        RECT  7.505000 58.770000  7.705000 58.970000 ;
        RECT  7.505000 59.180000  7.705000 59.380000 ;
        RECT  7.505000 59.590000  7.705000 59.790000 ;
        RECT  7.505000 60.000000  7.705000 60.200000 ;
        RECT  7.505000 60.410000  7.705000 60.610000 ;
        RECT  7.910000 56.310000  8.110000 56.510000 ;
        RECT  7.910000 56.720000  8.110000 56.920000 ;
        RECT  7.910000 57.130000  8.110000 57.330000 ;
        RECT  7.910000 57.540000  8.110000 57.740000 ;
        RECT  7.910000 57.950000  8.110000 58.150000 ;
        RECT  7.910000 58.360000  8.110000 58.560000 ;
        RECT  7.910000 58.770000  8.110000 58.970000 ;
        RECT  7.910000 59.180000  8.110000 59.380000 ;
        RECT  7.910000 59.590000  8.110000 59.790000 ;
        RECT  7.910000 60.000000  8.110000 60.200000 ;
        RECT  7.910000 60.410000  8.110000 60.610000 ;
        RECT  8.315000 56.310000  8.515000 56.510000 ;
        RECT  8.315000 56.720000  8.515000 56.920000 ;
        RECT  8.315000 57.130000  8.515000 57.330000 ;
        RECT  8.315000 57.540000  8.515000 57.740000 ;
        RECT  8.315000 57.950000  8.515000 58.150000 ;
        RECT  8.315000 58.360000  8.515000 58.560000 ;
        RECT  8.315000 58.770000  8.515000 58.970000 ;
        RECT  8.315000 59.180000  8.515000 59.380000 ;
        RECT  8.315000 59.590000  8.515000 59.790000 ;
        RECT  8.315000 60.000000  8.515000 60.200000 ;
        RECT  8.315000 60.410000  8.515000 60.610000 ;
        RECT  8.720000 56.310000  8.920000 56.510000 ;
        RECT  8.720000 56.720000  8.920000 56.920000 ;
        RECT  8.720000 57.130000  8.920000 57.330000 ;
        RECT  8.720000 57.540000  8.920000 57.740000 ;
        RECT  8.720000 57.950000  8.920000 58.150000 ;
        RECT  8.720000 58.360000  8.920000 58.560000 ;
        RECT  8.720000 58.770000  8.920000 58.970000 ;
        RECT  8.720000 59.180000  8.920000 59.380000 ;
        RECT  8.720000 59.590000  8.920000 59.790000 ;
        RECT  8.720000 60.000000  8.920000 60.200000 ;
        RECT  8.720000 60.410000  8.920000 60.610000 ;
        RECT  9.125000 56.310000  9.325000 56.510000 ;
        RECT  9.125000 56.720000  9.325000 56.920000 ;
        RECT  9.125000 57.130000  9.325000 57.330000 ;
        RECT  9.125000 57.540000  9.325000 57.740000 ;
        RECT  9.125000 57.950000  9.325000 58.150000 ;
        RECT  9.125000 58.360000  9.325000 58.560000 ;
        RECT  9.125000 58.770000  9.325000 58.970000 ;
        RECT  9.125000 59.180000  9.325000 59.380000 ;
        RECT  9.125000 59.590000  9.325000 59.790000 ;
        RECT  9.125000 60.000000  9.325000 60.200000 ;
        RECT  9.125000 60.410000  9.325000 60.610000 ;
        RECT  9.530000 56.310000  9.730000 56.510000 ;
        RECT  9.530000 56.720000  9.730000 56.920000 ;
        RECT  9.530000 57.130000  9.730000 57.330000 ;
        RECT  9.530000 57.540000  9.730000 57.740000 ;
        RECT  9.530000 57.950000  9.730000 58.150000 ;
        RECT  9.530000 58.360000  9.730000 58.560000 ;
        RECT  9.530000 58.770000  9.730000 58.970000 ;
        RECT  9.530000 59.180000  9.730000 59.380000 ;
        RECT  9.530000 59.590000  9.730000 59.790000 ;
        RECT  9.530000 60.000000  9.730000 60.200000 ;
        RECT  9.530000 60.410000  9.730000 60.610000 ;
        RECT  9.935000 56.310000 10.135000 56.510000 ;
        RECT  9.935000 56.720000 10.135000 56.920000 ;
        RECT  9.935000 57.130000 10.135000 57.330000 ;
        RECT  9.935000 57.540000 10.135000 57.740000 ;
        RECT  9.935000 57.950000 10.135000 58.150000 ;
        RECT  9.935000 58.360000 10.135000 58.560000 ;
        RECT  9.935000 58.770000 10.135000 58.970000 ;
        RECT  9.935000 59.180000 10.135000 59.380000 ;
        RECT  9.935000 59.590000 10.135000 59.790000 ;
        RECT  9.935000 60.000000 10.135000 60.200000 ;
        RECT  9.935000 60.410000 10.135000 60.610000 ;
        RECT 10.340000 56.310000 10.540000 56.510000 ;
        RECT 10.340000 56.720000 10.540000 56.920000 ;
        RECT 10.340000 57.130000 10.540000 57.330000 ;
        RECT 10.340000 57.540000 10.540000 57.740000 ;
        RECT 10.340000 57.950000 10.540000 58.150000 ;
        RECT 10.340000 58.360000 10.540000 58.560000 ;
        RECT 10.340000 58.770000 10.540000 58.970000 ;
        RECT 10.340000 59.180000 10.540000 59.380000 ;
        RECT 10.340000 59.590000 10.540000 59.790000 ;
        RECT 10.340000 60.000000 10.540000 60.200000 ;
        RECT 10.340000 60.410000 10.540000 60.610000 ;
        RECT 10.745000 56.310000 10.945000 56.510000 ;
        RECT 10.745000 56.720000 10.945000 56.920000 ;
        RECT 10.745000 57.130000 10.945000 57.330000 ;
        RECT 10.745000 57.540000 10.945000 57.740000 ;
        RECT 10.745000 57.950000 10.945000 58.150000 ;
        RECT 10.745000 58.360000 10.945000 58.560000 ;
        RECT 10.745000 58.770000 10.945000 58.970000 ;
        RECT 10.745000 59.180000 10.945000 59.380000 ;
        RECT 10.745000 59.590000 10.945000 59.790000 ;
        RECT 10.745000 60.000000 10.945000 60.200000 ;
        RECT 10.745000 60.410000 10.945000 60.610000 ;
        RECT 11.150000 56.310000 11.350000 56.510000 ;
        RECT 11.150000 56.720000 11.350000 56.920000 ;
        RECT 11.150000 57.130000 11.350000 57.330000 ;
        RECT 11.150000 57.540000 11.350000 57.740000 ;
        RECT 11.150000 57.950000 11.350000 58.150000 ;
        RECT 11.150000 58.360000 11.350000 58.560000 ;
        RECT 11.150000 58.770000 11.350000 58.970000 ;
        RECT 11.150000 59.180000 11.350000 59.380000 ;
        RECT 11.150000 59.590000 11.350000 59.790000 ;
        RECT 11.150000 60.000000 11.350000 60.200000 ;
        RECT 11.150000 60.410000 11.350000 60.610000 ;
        RECT 11.555000 56.310000 11.755000 56.510000 ;
        RECT 11.555000 56.720000 11.755000 56.920000 ;
        RECT 11.555000 57.130000 11.755000 57.330000 ;
        RECT 11.555000 57.540000 11.755000 57.740000 ;
        RECT 11.555000 57.950000 11.755000 58.150000 ;
        RECT 11.555000 58.360000 11.755000 58.560000 ;
        RECT 11.555000 58.770000 11.755000 58.970000 ;
        RECT 11.555000 59.180000 11.755000 59.380000 ;
        RECT 11.555000 59.590000 11.755000 59.790000 ;
        RECT 11.555000 60.000000 11.755000 60.200000 ;
        RECT 11.555000 60.410000 11.755000 60.610000 ;
        RECT 11.960000 56.310000 12.160000 56.510000 ;
        RECT 11.960000 56.720000 12.160000 56.920000 ;
        RECT 11.960000 57.130000 12.160000 57.330000 ;
        RECT 11.960000 57.540000 12.160000 57.740000 ;
        RECT 11.960000 57.950000 12.160000 58.150000 ;
        RECT 11.960000 58.360000 12.160000 58.560000 ;
        RECT 11.960000 58.770000 12.160000 58.970000 ;
        RECT 11.960000 59.180000 12.160000 59.380000 ;
        RECT 11.960000 59.590000 12.160000 59.790000 ;
        RECT 11.960000 60.000000 12.160000 60.200000 ;
        RECT 11.960000 60.410000 12.160000 60.610000 ;
        RECT 12.365000 56.310000 12.565000 56.510000 ;
        RECT 12.365000 56.720000 12.565000 56.920000 ;
        RECT 12.365000 57.130000 12.565000 57.330000 ;
        RECT 12.365000 57.540000 12.565000 57.740000 ;
        RECT 12.365000 57.950000 12.565000 58.150000 ;
        RECT 12.365000 58.360000 12.565000 58.560000 ;
        RECT 12.365000 58.770000 12.565000 58.970000 ;
        RECT 12.365000 59.180000 12.565000 59.380000 ;
        RECT 12.365000 59.590000 12.565000 59.790000 ;
        RECT 12.365000 60.000000 12.565000 60.200000 ;
        RECT 12.365000 60.410000 12.565000 60.610000 ;
        RECT 12.770000 56.310000 12.970000 56.510000 ;
        RECT 12.770000 56.720000 12.970000 56.920000 ;
        RECT 12.770000 57.130000 12.970000 57.330000 ;
        RECT 12.770000 57.540000 12.970000 57.740000 ;
        RECT 12.770000 57.950000 12.970000 58.150000 ;
        RECT 12.770000 58.360000 12.970000 58.560000 ;
        RECT 12.770000 58.770000 12.970000 58.970000 ;
        RECT 12.770000 59.180000 12.970000 59.380000 ;
        RECT 12.770000 59.590000 12.970000 59.790000 ;
        RECT 12.770000 60.000000 12.970000 60.200000 ;
        RECT 12.770000 60.410000 12.970000 60.610000 ;
        RECT 13.175000 56.310000 13.375000 56.510000 ;
        RECT 13.175000 56.720000 13.375000 56.920000 ;
        RECT 13.175000 57.130000 13.375000 57.330000 ;
        RECT 13.175000 57.540000 13.375000 57.740000 ;
        RECT 13.175000 57.950000 13.375000 58.150000 ;
        RECT 13.175000 58.360000 13.375000 58.560000 ;
        RECT 13.175000 58.770000 13.375000 58.970000 ;
        RECT 13.175000 59.180000 13.375000 59.380000 ;
        RECT 13.175000 59.590000 13.375000 59.790000 ;
        RECT 13.175000 60.000000 13.375000 60.200000 ;
        RECT 13.175000 60.410000 13.375000 60.610000 ;
        RECT 13.580000 56.310000 13.780000 56.510000 ;
        RECT 13.580000 56.720000 13.780000 56.920000 ;
        RECT 13.580000 57.130000 13.780000 57.330000 ;
        RECT 13.580000 57.540000 13.780000 57.740000 ;
        RECT 13.580000 57.950000 13.780000 58.150000 ;
        RECT 13.580000 58.360000 13.780000 58.560000 ;
        RECT 13.580000 58.770000 13.780000 58.970000 ;
        RECT 13.580000 59.180000 13.780000 59.380000 ;
        RECT 13.580000 59.590000 13.780000 59.790000 ;
        RECT 13.580000 60.000000 13.780000 60.200000 ;
        RECT 13.580000 60.410000 13.780000 60.610000 ;
        RECT 13.985000 56.310000 14.185000 56.510000 ;
        RECT 13.985000 56.720000 14.185000 56.920000 ;
        RECT 13.985000 57.130000 14.185000 57.330000 ;
        RECT 13.985000 57.540000 14.185000 57.740000 ;
        RECT 13.985000 57.950000 14.185000 58.150000 ;
        RECT 13.985000 58.360000 14.185000 58.560000 ;
        RECT 13.985000 58.770000 14.185000 58.970000 ;
        RECT 13.985000 59.180000 14.185000 59.380000 ;
        RECT 13.985000 59.590000 14.185000 59.790000 ;
        RECT 13.985000 60.000000 14.185000 60.200000 ;
        RECT 13.985000 60.410000 14.185000 60.610000 ;
        RECT 14.390000 56.310000 14.590000 56.510000 ;
        RECT 14.390000 56.720000 14.590000 56.920000 ;
        RECT 14.390000 57.130000 14.590000 57.330000 ;
        RECT 14.390000 57.540000 14.590000 57.740000 ;
        RECT 14.390000 57.950000 14.590000 58.150000 ;
        RECT 14.390000 58.360000 14.590000 58.560000 ;
        RECT 14.390000 58.770000 14.590000 58.970000 ;
        RECT 14.390000 59.180000 14.590000 59.380000 ;
        RECT 14.390000 59.590000 14.590000 59.790000 ;
        RECT 14.390000 60.000000 14.590000 60.200000 ;
        RECT 14.390000 60.410000 14.590000 60.610000 ;
        RECT 14.795000 56.310000 14.995000 56.510000 ;
        RECT 14.795000 56.720000 14.995000 56.920000 ;
        RECT 14.795000 57.130000 14.995000 57.330000 ;
        RECT 14.795000 57.540000 14.995000 57.740000 ;
        RECT 14.795000 57.950000 14.995000 58.150000 ;
        RECT 14.795000 58.360000 14.995000 58.560000 ;
        RECT 14.795000 58.770000 14.995000 58.970000 ;
        RECT 14.795000 59.180000 14.995000 59.380000 ;
        RECT 14.795000 59.590000 14.995000 59.790000 ;
        RECT 14.795000 60.000000 14.995000 60.200000 ;
        RECT 14.795000 60.410000 14.995000 60.610000 ;
        RECT 15.200000 56.310000 15.400000 56.510000 ;
        RECT 15.200000 56.720000 15.400000 56.920000 ;
        RECT 15.200000 57.130000 15.400000 57.330000 ;
        RECT 15.200000 57.540000 15.400000 57.740000 ;
        RECT 15.200000 57.950000 15.400000 58.150000 ;
        RECT 15.200000 58.360000 15.400000 58.560000 ;
        RECT 15.200000 58.770000 15.400000 58.970000 ;
        RECT 15.200000 59.180000 15.400000 59.380000 ;
        RECT 15.200000 59.590000 15.400000 59.790000 ;
        RECT 15.200000 60.000000 15.400000 60.200000 ;
        RECT 15.200000 60.410000 15.400000 60.610000 ;
        RECT 15.605000 56.310000 15.805000 56.510000 ;
        RECT 15.605000 56.720000 15.805000 56.920000 ;
        RECT 15.605000 57.130000 15.805000 57.330000 ;
        RECT 15.605000 57.540000 15.805000 57.740000 ;
        RECT 15.605000 57.950000 15.805000 58.150000 ;
        RECT 15.605000 58.360000 15.805000 58.560000 ;
        RECT 15.605000 58.770000 15.805000 58.970000 ;
        RECT 15.605000 59.180000 15.805000 59.380000 ;
        RECT 15.605000 59.590000 15.805000 59.790000 ;
        RECT 15.605000 60.000000 15.805000 60.200000 ;
        RECT 15.605000 60.410000 15.805000 60.610000 ;
        RECT 16.010000 56.310000 16.210000 56.510000 ;
        RECT 16.010000 56.720000 16.210000 56.920000 ;
        RECT 16.010000 57.130000 16.210000 57.330000 ;
        RECT 16.010000 57.540000 16.210000 57.740000 ;
        RECT 16.010000 57.950000 16.210000 58.150000 ;
        RECT 16.010000 58.360000 16.210000 58.560000 ;
        RECT 16.010000 58.770000 16.210000 58.970000 ;
        RECT 16.010000 59.180000 16.210000 59.380000 ;
        RECT 16.010000 59.590000 16.210000 59.790000 ;
        RECT 16.010000 60.000000 16.210000 60.200000 ;
        RECT 16.010000 60.410000 16.210000 60.610000 ;
        RECT 16.415000 56.310000 16.615000 56.510000 ;
        RECT 16.415000 56.720000 16.615000 56.920000 ;
        RECT 16.415000 57.130000 16.615000 57.330000 ;
        RECT 16.415000 57.540000 16.615000 57.740000 ;
        RECT 16.415000 57.950000 16.615000 58.150000 ;
        RECT 16.415000 58.360000 16.615000 58.560000 ;
        RECT 16.415000 58.770000 16.615000 58.970000 ;
        RECT 16.415000 59.180000 16.615000 59.380000 ;
        RECT 16.415000 59.590000 16.615000 59.790000 ;
        RECT 16.415000 60.000000 16.615000 60.200000 ;
        RECT 16.415000 60.410000 16.615000 60.610000 ;
        RECT 16.820000 56.310000 17.020000 56.510000 ;
        RECT 16.820000 56.720000 17.020000 56.920000 ;
        RECT 16.820000 57.130000 17.020000 57.330000 ;
        RECT 16.820000 57.540000 17.020000 57.740000 ;
        RECT 16.820000 57.950000 17.020000 58.150000 ;
        RECT 16.820000 58.360000 17.020000 58.560000 ;
        RECT 16.820000 58.770000 17.020000 58.970000 ;
        RECT 16.820000 59.180000 17.020000 59.380000 ;
        RECT 16.820000 59.590000 17.020000 59.790000 ;
        RECT 16.820000 60.000000 17.020000 60.200000 ;
        RECT 16.820000 60.410000 17.020000 60.610000 ;
        RECT 17.225000 56.310000 17.425000 56.510000 ;
        RECT 17.225000 56.720000 17.425000 56.920000 ;
        RECT 17.225000 57.130000 17.425000 57.330000 ;
        RECT 17.225000 57.540000 17.425000 57.740000 ;
        RECT 17.225000 57.950000 17.425000 58.150000 ;
        RECT 17.225000 58.360000 17.425000 58.560000 ;
        RECT 17.225000 58.770000 17.425000 58.970000 ;
        RECT 17.225000 59.180000 17.425000 59.380000 ;
        RECT 17.225000 59.590000 17.425000 59.790000 ;
        RECT 17.225000 60.000000 17.425000 60.200000 ;
        RECT 17.225000 60.410000 17.425000 60.610000 ;
        RECT 17.630000 56.310000 17.830000 56.510000 ;
        RECT 17.630000 56.720000 17.830000 56.920000 ;
        RECT 17.630000 57.130000 17.830000 57.330000 ;
        RECT 17.630000 57.540000 17.830000 57.740000 ;
        RECT 17.630000 57.950000 17.830000 58.150000 ;
        RECT 17.630000 58.360000 17.830000 58.560000 ;
        RECT 17.630000 58.770000 17.830000 58.970000 ;
        RECT 17.630000 59.180000 17.830000 59.380000 ;
        RECT 17.630000 59.590000 17.830000 59.790000 ;
        RECT 17.630000 60.000000 17.830000 60.200000 ;
        RECT 17.630000 60.410000 17.830000 60.610000 ;
        RECT 18.035000 56.310000 18.235000 56.510000 ;
        RECT 18.035000 56.720000 18.235000 56.920000 ;
        RECT 18.035000 57.130000 18.235000 57.330000 ;
        RECT 18.035000 57.540000 18.235000 57.740000 ;
        RECT 18.035000 57.950000 18.235000 58.150000 ;
        RECT 18.035000 58.360000 18.235000 58.560000 ;
        RECT 18.035000 58.770000 18.235000 58.970000 ;
        RECT 18.035000 59.180000 18.235000 59.380000 ;
        RECT 18.035000 59.590000 18.235000 59.790000 ;
        RECT 18.035000 60.000000 18.235000 60.200000 ;
        RECT 18.035000 60.410000 18.235000 60.610000 ;
        RECT 18.440000 56.310000 18.640000 56.510000 ;
        RECT 18.440000 56.720000 18.640000 56.920000 ;
        RECT 18.440000 57.130000 18.640000 57.330000 ;
        RECT 18.440000 57.540000 18.640000 57.740000 ;
        RECT 18.440000 57.950000 18.640000 58.150000 ;
        RECT 18.440000 58.360000 18.640000 58.560000 ;
        RECT 18.440000 58.770000 18.640000 58.970000 ;
        RECT 18.440000 59.180000 18.640000 59.380000 ;
        RECT 18.440000 59.590000 18.640000 59.790000 ;
        RECT 18.440000 60.000000 18.640000 60.200000 ;
        RECT 18.440000 60.410000 18.640000 60.610000 ;
        RECT 18.845000 56.310000 19.045000 56.510000 ;
        RECT 18.845000 56.720000 19.045000 56.920000 ;
        RECT 18.845000 57.130000 19.045000 57.330000 ;
        RECT 18.845000 57.540000 19.045000 57.740000 ;
        RECT 18.845000 57.950000 19.045000 58.150000 ;
        RECT 18.845000 58.360000 19.045000 58.560000 ;
        RECT 18.845000 58.770000 19.045000 58.970000 ;
        RECT 18.845000 59.180000 19.045000 59.380000 ;
        RECT 18.845000 59.590000 19.045000 59.790000 ;
        RECT 18.845000 60.000000 19.045000 60.200000 ;
        RECT 18.845000 60.410000 19.045000 60.610000 ;
        RECT 19.250000 56.310000 19.450000 56.510000 ;
        RECT 19.250000 56.720000 19.450000 56.920000 ;
        RECT 19.250000 57.130000 19.450000 57.330000 ;
        RECT 19.250000 57.540000 19.450000 57.740000 ;
        RECT 19.250000 57.950000 19.450000 58.150000 ;
        RECT 19.250000 58.360000 19.450000 58.560000 ;
        RECT 19.250000 58.770000 19.450000 58.970000 ;
        RECT 19.250000 59.180000 19.450000 59.380000 ;
        RECT 19.250000 59.590000 19.450000 59.790000 ;
        RECT 19.250000 60.000000 19.450000 60.200000 ;
        RECT 19.250000 60.410000 19.450000 60.610000 ;
        RECT 19.655000 56.310000 19.855000 56.510000 ;
        RECT 19.655000 56.720000 19.855000 56.920000 ;
        RECT 19.655000 57.130000 19.855000 57.330000 ;
        RECT 19.655000 57.540000 19.855000 57.740000 ;
        RECT 19.655000 57.950000 19.855000 58.150000 ;
        RECT 19.655000 58.360000 19.855000 58.560000 ;
        RECT 19.655000 58.770000 19.855000 58.970000 ;
        RECT 19.655000 59.180000 19.855000 59.380000 ;
        RECT 19.655000 59.590000 19.855000 59.790000 ;
        RECT 19.655000 60.000000 19.855000 60.200000 ;
        RECT 19.655000 60.410000 19.855000 60.610000 ;
        RECT 20.060000 56.310000 20.260000 56.510000 ;
        RECT 20.060000 56.720000 20.260000 56.920000 ;
        RECT 20.060000 57.130000 20.260000 57.330000 ;
        RECT 20.060000 57.540000 20.260000 57.740000 ;
        RECT 20.060000 57.950000 20.260000 58.150000 ;
        RECT 20.060000 58.360000 20.260000 58.560000 ;
        RECT 20.060000 58.770000 20.260000 58.970000 ;
        RECT 20.060000 59.180000 20.260000 59.380000 ;
        RECT 20.060000 59.590000 20.260000 59.790000 ;
        RECT 20.060000 60.000000 20.260000 60.200000 ;
        RECT 20.060000 60.410000 20.260000 60.610000 ;
        RECT 20.465000 56.310000 20.665000 56.510000 ;
        RECT 20.465000 56.720000 20.665000 56.920000 ;
        RECT 20.465000 57.130000 20.665000 57.330000 ;
        RECT 20.465000 57.540000 20.665000 57.740000 ;
        RECT 20.465000 57.950000 20.665000 58.150000 ;
        RECT 20.465000 58.360000 20.665000 58.560000 ;
        RECT 20.465000 58.770000 20.665000 58.970000 ;
        RECT 20.465000 59.180000 20.665000 59.380000 ;
        RECT 20.465000 59.590000 20.665000 59.790000 ;
        RECT 20.465000 60.000000 20.665000 60.200000 ;
        RECT 20.465000 60.410000 20.665000 60.610000 ;
        RECT 20.870000 56.310000 21.070000 56.510000 ;
        RECT 20.870000 56.720000 21.070000 56.920000 ;
        RECT 20.870000 57.130000 21.070000 57.330000 ;
        RECT 20.870000 57.540000 21.070000 57.740000 ;
        RECT 20.870000 57.950000 21.070000 58.150000 ;
        RECT 20.870000 58.360000 21.070000 58.560000 ;
        RECT 20.870000 58.770000 21.070000 58.970000 ;
        RECT 20.870000 59.180000 21.070000 59.380000 ;
        RECT 20.870000 59.590000 21.070000 59.790000 ;
        RECT 20.870000 60.000000 21.070000 60.200000 ;
        RECT 20.870000 60.410000 21.070000 60.610000 ;
        RECT 21.275000 56.310000 21.475000 56.510000 ;
        RECT 21.275000 56.720000 21.475000 56.920000 ;
        RECT 21.275000 57.130000 21.475000 57.330000 ;
        RECT 21.275000 57.540000 21.475000 57.740000 ;
        RECT 21.275000 57.950000 21.475000 58.150000 ;
        RECT 21.275000 58.360000 21.475000 58.560000 ;
        RECT 21.275000 58.770000 21.475000 58.970000 ;
        RECT 21.275000 59.180000 21.475000 59.380000 ;
        RECT 21.275000 59.590000 21.475000 59.790000 ;
        RECT 21.275000 60.000000 21.475000 60.200000 ;
        RECT 21.275000 60.410000 21.475000 60.610000 ;
        RECT 21.680000 56.310000 21.880000 56.510000 ;
        RECT 21.680000 56.720000 21.880000 56.920000 ;
        RECT 21.680000 57.130000 21.880000 57.330000 ;
        RECT 21.680000 57.540000 21.880000 57.740000 ;
        RECT 21.680000 57.950000 21.880000 58.150000 ;
        RECT 21.680000 58.360000 21.880000 58.560000 ;
        RECT 21.680000 58.770000 21.880000 58.970000 ;
        RECT 21.680000 59.180000 21.880000 59.380000 ;
        RECT 21.680000 59.590000 21.880000 59.790000 ;
        RECT 21.680000 60.000000 21.880000 60.200000 ;
        RECT 21.680000 60.410000 21.880000 60.610000 ;
        RECT 22.085000 56.310000 22.285000 56.510000 ;
        RECT 22.085000 56.720000 22.285000 56.920000 ;
        RECT 22.085000 57.130000 22.285000 57.330000 ;
        RECT 22.085000 57.540000 22.285000 57.740000 ;
        RECT 22.085000 57.950000 22.285000 58.150000 ;
        RECT 22.085000 58.360000 22.285000 58.560000 ;
        RECT 22.085000 58.770000 22.285000 58.970000 ;
        RECT 22.085000 59.180000 22.285000 59.380000 ;
        RECT 22.085000 59.590000 22.285000 59.790000 ;
        RECT 22.085000 60.000000 22.285000 60.200000 ;
        RECT 22.085000 60.410000 22.285000 60.610000 ;
        RECT 22.490000 56.310000 22.690000 56.510000 ;
        RECT 22.490000 56.720000 22.690000 56.920000 ;
        RECT 22.490000 57.130000 22.690000 57.330000 ;
        RECT 22.490000 57.540000 22.690000 57.740000 ;
        RECT 22.490000 57.950000 22.690000 58.150000 ;
        RECT 22.490000 58.360000 22.690000 58.560000 ;
        RECT 22.490000 58.770000 22.690000 58.970000 ;
        RECT 22.490000 59.180000 22.690000 59.380000 ;
        RECT 22.490000 59.590000 22.690000 59.790000 ;
        RECT 22.490000 60.000000 22.690000 60.200000 ;
        RECT 22.490000 60.410000 22.690000 60.610000 ;
        RECT 22.895000 56.310000 23.095000 56.510000 ;
        RECT 22.895000 56.720000 23.095000 56.920000 ;
        RECT 22.895000 57.130000 23.095000 57.330000 ;
        RECT 22.895000 57.540000 23.095000 57.740000 ;
        RECT 22.895000 57.950000 23.095000 58.150000 ;
        RECT 22.895000 58.360000 23.095000 58.560000 ;
        RECT 22.895000 58.770000 23.095000 58.970000 ;
        RECT 22.895000 59.180000 23.095000 59.380000 ;
        RECT 22.895000 59.590000 23.095000 59.790000 ;
        RECT 22.895000 60.000000 23.095000 60.200000 ;
        RECT 22.895000 60.410000 23.095000 60.610000 ;
        RECT 23.300000 56.310000 23.500000 56.510000 ;
        RECT 23.300000 56.720000 23.500000 56.920000 ;
        RECT 23.300000 57.130000 23.500000 57.330000 ;
        RECT 23.300000 57.540000 23.500000 57.740000 ;
        RECT 23.300000 57.950000 23.500000 58.150000 ;
        RECT 23.300000 58.360000 23.500000 58.560000 ;
        RECT 23.300000 58.770000 23.500000 58.970000 ;
        RECT 23.300000 59.180000 23.500000 59.380000 ;
        RECT 23.300000 59.590000 23.500000 59.790000 ;
        RECT 23.300000 60.000000 23.500000 60.200000 ;
        RECT 23.300000 60.410000 23.500000 60.610000 ;
        RECT 23.705000 56.310000 23.905000 56.510000 ;
        RECT 23.705000 56.720000 23.905000 56.920000 ;
        RECT 23.705000 57.130000 23.905000 57.330000 ;
        RECT 23.705000 57.540000 23.905000 57.740000 ;
        RECT 23.705000 57.950000 23.905000 58.150000 ;
        RECT 23.705000 58.360000 23.905000 58.560000 ;
        RECT 23.705000 58.770000 23.905000 58.970000 ;
        RECT 23.705000 59.180000 23.905000 59.380000 ;
        RECT 23.705000 59.590000 23.905000 59.790000 ;
        RECT 23.705000 60.000000 23.905000 60.200000 ;
        RECT 23.705000 60.410000 23.905000 60.610000 ;
        RECT 24.110000 56.310000 24.310000 56.510000 ;
        RECT 24.110000 56.720000 24.310000 56.920000 ;
        RECT 24.110000 57.130000 24.310000 57.330000 ;
        RECT 24.110000 57.540000 24.310000 57.740000 ;
        RECT 24.110000 57.950000 24.310000 58.150000 ;
        RECT 24.110000 58.360000 24.310000 58.560000 ;
        RECT 24.110000 58.770000 24.310000 58.970000 ;
        RECT 24.110000 59.180000 24.310000 59.380000 ;
        RECT 24.110000 59.590000 24.310000 59.790000 ;
        RECT 24.110000 60.000000 24.310000 60.200000 ;
        RECT 24.110000 60.410000 24.310000 60.610000 ;
        RECT 50.845000 56.310000 51.045000 56.510000 ;
        RECT 50.845000 56.720000 51.045000 56.920000 ;
        RECT 50.845000 57.130000 51.045000 57.330000 ;
        RECT 50.845000 57.540000 51.045000 57.740000 ;
        RECT 50.845000 57.950000 51.045000 58.150000 ;
        RECT 50.845000 58.360000 51.045000 58.560000 ;
        RECT 50.845000 58.770000 51.045000 58.970000 ;
        RECT 50.845000 59.180000 51.045000 59.380000 ;
        RECT 50.845000 59.590000 51.045000 59.790000 ;
        RECT 50.845000 60.000000 51.045000 60.200000 ;
        RECT 50.845000 60.410000 51.045000 60.610000 ;
        RECT 51.255000 56.310000 51.455000 56.510000 ;
        RECT 51.255000 56.720000 51.455000 56.920000 ;
        RECT 51.255000 57.130000 51.455000 57.330000 ;
        RECT 51.255000 57.540000 51.455000 57.740000 ;
        RECT 51.255000 57.950000 51.455000 58.150000 ;
        RECT 51.255000 58.360000 51.455000 58.560000 ;
        RECT 51.255000 58.770000 51.455000 58.970000 ;
        RECT 51.255000 59.180000 51.455000 59.380000 ;
        RECT 51.255000 59.590000 51.455000 59.790000 ;
        RECT 51.255000 60.000000 51.455000 60.200000 ;
        RECT 51.255000 60.410000 51.455000 60.610000 ;
        RECT 51.665000 56.310000 51.865000 56.510000 ;
        RECT 51.665000 56.720000 51.865000 56.920000 ;
        RECT 51.665000 57.130000 51.865000 57.330000 ;
        RECT 51.665000 57.540000 51.865000 57.740000 ;
        RECT 51.665000 57.950000 51.865000 58.150000 ;
        RECT 51.665000 58.360000 51.865000 58.560000 ;
        RECT 51.665000 58.770000 51.865000 58.970000 ;
        RECT 51.665000 59.180000 51.865000 59.380000 ;
        RECT 51.665000 59.590000 51.865000 59.790000 ;
        RECT 51.665000 60.000000 51.865000 60.200000 ;
        RECT 51.665000 60.410000 51.865000 60.610000 ;
        RECT 52.075000 56.310000 52.275000 56.510000 ;
        RECT 52.075000 56.720000 52.275000 56.920000 ;
        RECT 52.075000 57.130000 52.275000 57.330000 ;
        RECT 52.075000 57.540000 52.275000 57.740000 ;
        RECT 52.075000 57.950000 52.275000 58.150000 ;
        RECT 52.075000 58.360000 52.275000 58.560000 ;
        RECT 52.075000 58.770000 52.275000 58.970000 ;
        RECT 52.075000 59.180000 52.275000 59.380000 ;
        RECT 52.075000 59.590000 52.275000 59.790000 ;
        RECT 52.075000 60.000000 52.275000 60.200000 ;
        RECT 52.075000 60.410000 52.275000 60.610000 ;
        RECT 52.485000 56.310000 52.685000 56.510000 ;
        RECT 52.485000 56.720000 52.685000 56.920000 ;
        RECT 52.485000 57.130000 52.685000 57.330000 ;
        RECT 52.485000 57.540000 52.685000 57.740000 ;
        RECT 52.485000 57.950000 52.685000 58.150000 ;
        RECT 52.485000 58.360000 52.685000 58.560000 ;
        RECT 52.485000 58.770000 52.685000 58.970000 ;
        RECT 52.485000 59.180000 52.685000 59.380000 ;
        RECT 52.485000 59.590000 52.685000 59.790000 ;
        RECT 52.485000 60.000000 52.685000 60.200000 ;
        RECT 52.485000 60.410000 52.685000 60.610000 ;
        RECT 52.895000 56.310000 53.095000 56.510000 ;
        RECT 52.895000 56.720000 53.095000 56.920000 ;
        RECT 52.895000 57.130000 53.095000 57.330000 ;
        RECT 52.895000 57.540000 53.095000 57.740000 ;
        RECT 52.895000 57.950000 53.095000 58.150000 ;
        RECT 52.895000 58.360000 53.095000 58.560000 ;
        RECT 52.895000 58.770000 53.095000 58.970000 ;
        RECT 52.895000 59.180000 53.095000 59.380000 ;
        RECT 52.895000 59.590000 53.095000 59.790000 ;
        RECT 52.895000 60.000000 53.095000 60.200000 ;
        RECT 52.895000 60.410000 53.095000 60.610000 ;
        RECT 53.305000 56.310000 53.505000 56.510000 ;
        RECT 53.305000 56.720000 53.505000 56.920000 ;
        RECT 53.305000 57.130000 53.505000 57.330000 ;
        RECT 53.305000 57.540000 53.505000 57.740000 ;
        RECT 53.305000 57.950000 53.505000 58.150000 ;
        RECT 53.305000 58.360000 53.505000 58.560000 ;
        RECT 53.305000 58.770000 53.505000 58.970000 ;
        RECT 53.305000 59.180000 53.505000 59.380000 ;
        RECT 53.305000 59.590000 53.505000 59.790000 ;
        RECT 53.305000 60.000000 53.505000 60.200000 ;
        RECT 53.305000 60.410000 53.505000 60.610000 ;
        RECT 53.715000 56.310000 53.915000 56.510000 ;
        RECT 53.715000 56.720000 53.915000 56.920000 ;
        RECT 53.715000 57.130000 53.915000 57.330000 ;
        RECT 53.715000 57.540000 53.915000 57.740000 ;
        RECT 53.715000 57.950000 53.915000 58.150000 ;
        RECT 53.715000 58.360000 53.915000 58.560000 ;
        RECT 53.715000 58.770000 53.915000 58.970000 ;
        RECT 53.715000 59.180000 53.915000 59.380000 ;
        RECT 53.715000 59.590000 53.915000 59.790000 ;
        RECT 53.715000 60.000000 53.915000 60.200000 ;
        RECT 53.715000 60.410000 53.915000 60.610000 ;
        RECT 54.125000 56.310000 54.325000 56.510000 ;
        RECT 54.125000 56.720000 54.325000 56.920000 ;
        RECT 54.125000 57.130000 54.325000 57.330000 ;
        RECT 54.125000 57.540000 54.325000 57.740000 ;
        RECT 54.125000 57.950000 54.325000 58.150000 ;
        RECT 54.125000 58.360000 54.325000 58.560000 ;
        RECT 54.125000 58.770000 54.325000 58.970000 ;
        RECT 54.125000 59.180000 54.325000 59.380000 ;
        RECT 54.125000 59.590000 54.325000 59.790000 ;
        RECT 54.125000 60.000000 54.325000 60.200000 ;
        RECT 54.125000 60.410000 54.325000 60.610000 ;
        RECT 54.535000 56.310000 54.735000 56.510000 ;
        RECT 54.535000 56.720000 54.735000 56.920000 ;
        RECT 54.535000 57.130000 54.735000 57.330000 ;
        RECT 54.535000 57.540000 54.735000 57.740000 ;
        RECT 54.535000 57.950000 54.735000 58.150000 ;
        RECT 54.535000 58.360000 54.735000 58.560000 ;
        RECT 54.535000 58.770000 54.735000 58.970000 ;
        RECT 54.535000 59.180000 54.735000 59.380000 ;
        RECT 54.535000 59.590000 54.735000 59.790000 ;
        RECT 54.535000 60.000000 54.735000 60.200000 ;
        RECT 54.535000 60.410000 54.735000 60.610000 ;
        RECT 54.945000 56.310000 55.145000 56.510000 ;
        RECT 54.945000 56.720000 55.145000 56.920000 ;
        RECT 54.945000 57.130000 55.145000 57.330000 ;
        RECT 54.945000 57.540000 55.145000 57.740000 ;
        RECT 54.945000 57.950000 55.145000 58.150000 ;
        RECT 54.945000 58.360000 55.145000 58.560000 ;
        RECT 54.945000 58.770000 55.145000 58.970000 ;
        RECT 54.945000 59.180000 55.145000 59.380000 ;
        RECT 54.945000 59.590000 55.145000 59.790000 ;
        RECT 54.945000 60.000000 55.145000 60.200000 ;
        RECT 54.945000 60.410000 55.145000 60.610000 ;
        RECT 55.355000 56.310000 55.555000 56.510000 ;
        RECT 55.355000 56.720000 55.555000 56.920000 ;
        RECT 55.355000 57.130000 55.555000 57.330000 ;
        RECT 55.355000 57.540000 55.555000 57.740000 ;
        RECT 55.355000 57.950000 55.555000 58.150000 ;
        RECT 55.355000 58.360000 55.555000 58.560000 ;
        RECT 55.355000 58.770000 55.555000 58.970000 ;
        RECT 55.355000 59.180000 55.555000 59.380000 ;
        RECT 55.355000 59.590000 55.555000 59.790000 ;
        RECT 55.355000 60.000000 55.555000 60.200000 ;
        RECT 55.355000 60.410000 55.555000 60.610000 ;
        RECT 55.765000 56.310000 55.965000 56.510000 ;
        RECT 55.765000 56.720000 55.965000 56.920000 ;
        RECT 55.765000 57.130000 55.965000 57.330000 ;
        RECT 55.765000 57.540000 55.965000 57.740000 ;
        RECT 55.765000 57.950000 55.965000 58.150000 ;
        RECT 55.765000 58.360000 55.965000 58.560000 ;
        RECT 55.765000 58.770000 55.965000 58.970000 ;
        RECT 55.765000 59.180000 55.965000 59.380000 ;
        RECT 55.765000 59.590000 55.965000 59.790000 ;
        RECT 55.765000 60.000000 55.965000 60.200000 ;
        RECT 55.765000 60.410000 55.965000 60.610000 ;
        RECT 56.175000 56.310000 56.375000 56.510000 ;
        RECT 56.175000 56.720000 56.375000 56.920000 ;
        RECT 56.175000 57.130000 56.375000 57.330000 ;
        RECT 56.175000 57.540000 56.375000 57.740000 ;
        RECT 56.175000 57.950000 56.375000 58.150000 ;
        RECT 56.175000 58.360000 56.375000 58.560000 ;
        RECT 56.175000 58.770000 56.375000 58.970000 ;
        RECT 56.175000 59.180000 56.375000 59.380000 ;
        RECT 56.175000 59.590000 56.375000 59.790000 ;
        RECT 56.175000 60.000000 56.375000 60.200000 ;
        RECT 56.175000 60.410000 56.375000 60.610000 ;
        RECT 56.585000 56.310000 56.785000 56.510000 ;
        RECT 56.585000 56.720000 56.785000 56.920000 ;
        RECT 56.585000 57.130000 56.785000 57.330000 ;
        RECT 56.585000 57.540000 56.785000 57.740000 ;
        RECT 56.585000 57.950000 56.785000 58.150000 ;
        RECT 56.585000 58.360000 56.785000 58.560000 ;
        RECT 56.585000 58.770000 56.785000 58.970000 ;
        RECT 56.585000 59.180000 56.785000 59.380000 ;
        RECT 56.585000 59.590000 56.785000 59.790000 ;
        RECT 56.585000 60.000000 56.785000 60.200000 ;
        RECT 56.585000 60.410000 56.785000 60.610000 ;
        RECT 56.990000 56.310000 57.190000 56.510000 ;
        RECT 56.990000 56.720000 57.190000 56.920000 ;
        RECT 56.990000 57.130000 57.190000 57.330000 ;
        RECT 56.990000 57.540000 57.190000 57.740000 ;
        RECT 56.990000 57.950000 57.190000 58.150000 ;
        RECT 56.990000 58.360000 57.190000 58.560000 ;
        RECT 56.990000 58.770000 57.190000 58.970000 ;
        RECT 56.990000 59.180000 57.190000 59.380000 ;
        RECT 56.990000 59.590000 57.190000 59.790000 ;
        RECT 56.990000 60.000000 57.190000 60.200000 ;
        RECT 56.990000 60.410000 57.190000 60.610000 ;
        RECT 57.395000 56.310000 57.595000 56.510000 ;
        RECT 57.395000 56.720000 57.595000 56.920000 ;
        RECT 57.395000 57.130000 57.595000 57.330000 ;
        RECT 57.395000 57.540000 57.595000 57.740000 ;
        RECT 57.395000 57.950000 57.595000 58.150000 ;
        RECT 57.395000 58.360000 57.595000 58.560000 ;
        RECT 57.395000 58.770000 57.595000 58.970000 ;
        RECT 57.395000 59.180000 57.595000 59.380000 ;
        RECT 57.395000 59.590000 57.595000 59.790000 ;
        RECT 57.395000 60.000000 57.595000 60.200000 ;
        RECT 57.395000 60.410000 57.595000 60.610000 ;
        RECT 57.800000 56.310000 58.000000 56.510000 ;
        RECT 57.800000 56.720000 58.000000 56.920000 ;
        RECT 57.800000 57.130000 58.000000 57.330000 ;
        RECT 57.800000 57.540000 58.000000 57.740000 ;
        RECT 57.800000 57.950000 58.000000 58.150000 ;
        RECT 57.800000 58.360000 58.000000 58.560000 ;
        RECT 57.800000 58.770000 58.000000 58.970000 ;
        RECT 57.800000 59.180000 58.000000 59.380000 ;
        RECT 57.800000 59.590000 58.000000 59.790000 ;
        RECT 57.800000 60.000000 58.000000 60.200000 ;
        RECT 57.800000 60.410000 58.000000 60.610000 ;
        RECT 58.205000 56.310000 58.405000 56.510000 ;
        RECT 58.205000 56.720000 58.405000 56.920000 ;
        RECT 58.205000 57.130000 58.405000 57.330000 ;
        RECT 58.205000 57.540000 58.405000 57.740000 ;
        RECT 58.205000 57.950000 58.405000 58.150000 ;
        RECT 58.205000 58.360000 58.405000 58.560000 ;
        RECT 58.205000 58.770000 58.405000 58.970000 ;
        RECT 58.205000 59.180000 58.405000 59.380000 ;
        RECT 58.205000 59.590000 58.405000 59.790000 ;
        RECT 58.205000 60.000000 58.405000 60.200000 ;
        RECT 58.205000 60.410000 58.405000 60.610000 ;
        RECT 58.610000 56.310000 58.810000 56.510000 ;
        RECT 58.610000 56.720000 58.810000 56.920000 ;
        RECT 58.610000 57.130000 58.810000 57.330000 ;
        RECT 58.610000 57.540000 58.810000 57.740000 ;
        RECT 58.610000 57.950000 58.810000 58.150000 ;
        RECT 58.610000 58.360000 58.810000 58.560000 ;
        RECT 58.610000 58.770000 58.810000 58.970000 ;
        RECT 58.610000 59.180000 58.810000 59.380000 ;
        RECT 58.610000 59.590000 58.810000 59.790000 ;
        RECT 58.610000 60.000000 58.810000 60.200000 ;
        RECT 58.610000 60.410000 58.810000 60.610000 ;
        RECT 59.015000 56.310000 59.215000 56.510000 ;
        RECT 59.015000 56.720000 59.215000 56.920000 ;
        RECT 59.015000 57.130000 59.215000 57.330000 ;
        RECT 59.015000 57.540000 59.215000 57.740000 ;
        RECT 59.015000 57.950000 59.215000 58.150000 ;
        RECT 59.015000 58.360000 59.215000 58.560000 ;
        RECT 59.015000 58.770000 59.215000 58.970000 ;
        RECT 59.015000 59.180000 59.215000 59.380000 ;
        RECT 59.015000 59.590000 59.215000 59.790000 ;
        RECT 59.015000 60.000000 59.215000 60.200000 ;
        RECT 59.015000 60.410000 59.215000 60.610000 ;
        RECT 59.420000 56.310000 59.620000 56.510000 ;
        RECT 59.420000 56.720000 59.620000 56.920000 ;
        RECT 59.420000 57.130000 59.620000 57.330000 ;
        RECT 59.420000 57.540000 59.620000 57.740000 ;
        RECT 59.420000 57.950000 59.620000 58.150000 ;
        RECT 59.420000 58.360000 59.620000 58.560000 ;
        RECT 59.420000 58.770000 59.620000 58.970000 ;
        RECT 59.420000 59.180000 59.620000 59.380000 ;
        RECT 59.420000 59.590000 59.620000 59.790000 ;
        RECT 59.420000 60.000000 59.620000 60.200000 ;
        RECT 59.420000 60.410000 59.620000 60.610000 ;
        RECT 59.825000 56.310000 60.025000 56.510000 ;
        RECT 59.825000 56.720000 60.025000 56.920000 ;
        RECT 59.825000 57.130000 60.025000 57.330000 ;
        RECT 59.825000 57.540000 60.025000 57.740000 ;
        RECT 59.825000 57.950000 60.025000 58.150000 ;
        RECT 59.825000 58.360000 60.025000 58.560000 ;
        RECT 59.825000 58.770000 60.025000 58.970000 ;
        RECT 59.825000 59.180000 60.025000 59.380000 ;
        RECT 59.825000 59.590000 60.025000 59.790000 ;
        RECT 59.825000 60.000000 60.025000 60.200000 ;
        RECT 59.825000 60.410000 60.025000 60.610000 ;
        RECT 60.230000 56.310000 60.430000 56.510000 ;
        RECT 60.230000 56.720000 60.430000 56.920000 ;
        RECT 60.230000 57.130000 60.430000 57.330000 ;
        RECT 60.230000 57.540000 60.430000 57.740000 ;
        RECT 60.230000 57.950000 60.430000 58.150000 ;
        RECT 60.230000 58.360000 60.430000 58.560000 ;
        RECT 60.230000 58.770000 60.430000 58.970000 ;
        RECT 60.230000 59.180000 60.430000 59.380000 ;
        RECT 60.230000 59.590000 60.430000 59.790000 ;
        RECT 60.230000 60.000000 60.430000 60.200000 ;
        RECT 60.230000 60.410000 60.430000 60.610000 ;
        RECT 60.635000 56.310000 60.835000 56.510000 ;
        RECT 60.635000 56.720000 60.835000 56.920000 ;
        RECT 60.635000 57.130000 60.835000 57.330000 ;
        RECT 60.635000 57.540000 60.835000 57.740000 ;
        RECT 60.635000 57.950000 60.835000 58.150000 ;
        RECT 60.635000 58.360000 60.835000 58.560000 ;
        RECT 60.635000 58.770000 60.835000 58.970000 ;
        RECT 60.635000 59.180000 60.835000 59.380000 ;
        RECT 60.635000 59.590000 60.835000 59.790000 ;
        RECT 60.635000 60.000000 60.835000 60.200000 ;
        RECT 60.635000 60.410000 60.835000 60.610000 ;
        RECT 61.040000 56.310000 61.240000 56.510000 ;
        RECT 61.040000 56.720000 61.240000 56.920000 ;
        RECT 61.040000 57.130000 61.240000 57.330000 ;
        RECT 61.040000 57.540000 61.240000 57.740000 ;
        RECT 61.040000 57.950000 61.240000 58.150000 ;
        RECT 61.040000 58.360000 61.240000 58.560000 ;
        RECT 61.040000 58.770000 61.240000 58.970000 ;
        RECT 61.040000 59.180000 61.240000 59.380000 ;
        RECT 61.040000 59.590000 61.240000 59.790000 ;
        RECT 61.040000 60.000000 61.240000 60.200000 ;
        RECT 61.040000 60.410000 61.240000 60.610000 ;
        RECT 61.445000 56.310000 61.645000 56.510000 ;
        RECT 61.445000 56.720000 61.645000 56.920000 ;
        RECT 61.445000 57.130000 61.645000 57.330000 ;
        RECT 61.445000 57.540000 61.645000 57.740000 ;
        RECT 61.445000 57.950000 61.645000 58.150000 ;
        RECT 61.445000 58.360000 61.645000 58.560000 ;
        RECT 61.445000 58.770000 61.645000 58.970000 ;
        RECT 61.445000 59.180000 61.645000 59.380000 ;
        RECT 61.445000 59.590000 61.645000 59.790000 ;
        RECT 61.445000 60.000000 61.645000 60.200000 ;
        RECT 61.445000 60.410000 61.645000 60.610000 ;
        RECT 61.850000 56.310000 62.050000 56.510000 ;
        RECT 61.850000 56.720000 62.050000 56.920000 ;
        RECT 61.850000 57.130000 62.050000 57.330000 ;
        RECT 61.850000 57.540000 62.050000 57.740000 ;
        RECT 61.850000 57.950000 62.050000 58.150000 ;
        RECT 61.850000 58.360000 62.050000 58.560000 ;
        RECT 61.850000 58.770000 62.050000 58.970000 ;
        RECT 61.850000 59.180000 62.050000 59.380000 ;
        RECT 61.850000 59.590000 62.050000 59.790000 ;
        RECT 61.850000 60.000000 62.050000 60.200000 ;
        RECT 61.850000 60.410000 62.050000 60.610000 ;
        RECT 62.255000 56.310000 62.455000 56.510000 ;
        RECT 62.255000 56.720000 62.455000 56.920000 ;
        RECT 62.255000 57.130000 62.455000 57.330000 ;
        RECT 62.255000 57.540000 62.455000 57.740000 ;
        RECT 62.255000 57.950000 62.455000 58.150000 ;
        RECT 62.255000 58.360000 62.455000 58.560000 ;
        RECT 62.255000 58.770000 62.455000 58.970000 ;
        RECT 62.255000 59.180000 62.455000 59.380000 ;
        RECT 62.255000 59.590000 62.455000 59.790000 ;
        RECT 62.255000 60.000000 62.455000 60.200000 ;
        RECT 62.255000 60.410000 62.455000 60.610000 ;
        RECT 62.660000 56.310000 62.860000 56.510000 ;
        RECT 62.660000 56.720000 62.860000 56.920000 ;
        RECT 62.660000 57.130000 62.860000 57.330000 ;
        RECT 62.660000 57.540000 62.860000 57.740000 ;
        RECT 62.660000 57.950000 62.860000 58.150000 ;
        RECT 62.660000 58.360000 62.860000 58.560000 ;
        RECT 62.660000 58.770000 62.860000 58.970000 ;
        RECT 62.660000 59.180000 62.860000 59.380000 ;
        RECT 62.660000 59.590000 62.860000 59.790000 ;
        RECT 62.660000 60.000000 62.860000 60.200000 ;
        RECT 62.660000 60.410000 62.860000 60.610000 ;
        RECT 63.065000 56.310000 63.265000 56.510000 ;
        RECT 63.065000 56.720000 63.265000 56.920000 ;
        RECT 63.065000 57.130000 63.265000 57.330000 ;
        RECT 63.065000 57.540000 63.265000 57.740000 ;
        RECT 63.065000 57.950000 63.265000 58.150000 ;
        RECT 63.065000 58.360000 63.265000 58.560000 ;
        RECT 63.065000 58.770000 63.265000 58.970000 ;
        RECT 63.065000 59.180000 63.265000 59.380000 ;
        RECT 63.065000 59.590000 63.265000 59.790000 ;
        RECT 63.065000 60.000000 63.265000 60.200000 ;
        RECT 63.065000 60.410000 63.265000 60.610000 ;
        RECT 63.470000 56.310000 63.670000 56.510000 ;
        RECT 63.470000 56.720000 63.670000 56.920000 ;
        RECT 63.470000 57.130000 63.670000 57.330000 ;
        RECT 63.470000 57.540000 63.670000 57.740000 ;
        RECT 63.470000 57.950000 63.670000 58.150000 ;
        RECT 63.470000 58.360000 63.670000 58.560000 ;
        RECT 63.470000 58.770000 63.670000 58.970000 ;
        RECT 63.470000 59.180000 63.670000 59.380000 ;
        RECT 63.470000 59.590000 63.670000 59.790000 ;
        RECT 63.470000 60.000000 63.670000 60.200000 ;
        RECT 63.470000 60.410000 63.670000 60.610000 ;
        RECT 63.875000 56.310000 64.075000 56.510000 ;
        RECT 63.875000 56.720000 64.075000 56.920000 ;
        RECT 63.875000 57.130000 64.075000 57.330000 ;
        RECT 63.875000 57.540000 64.075000 57.740000 ;
        RECT 63.875000 57.950000 64.075000 58.150000 ;
        RECT 63.875000 58.360000 64.075000 58.560000 ;
        RECT 63.875000 58.770000 64.075000 58.970000 ;
        RECT 63.875000 59.180000 64.075000 59.380000 ;
        RECT 63.875000 59.590000 64.075000 59.790000 ;
        RECT 63.875000 60.000000 64.075000 60.200000 ;
        RECT 63.875000 60.410000 64.075000 60.610000 ;
        RECT 64.280000 56.310000 64.480000 56.510000 ;
        RECT 64.280000 56.720000 64.480000 56.920000 ;
        RECT 64.280000 57.130000 64.480000 57.330000 ;
        RECT 64.280000 57.540000 64.480000 57.740000 ;
        RECT 64.280000 57.950000 64.480000 58.150000 ;
        RECT 64.280000 58.360000 64.480000 58.560000 ;
        RECT 64.280000 58.770000 64.480000 58.970000 ;
        RECT 64.280000 59.180000 64.480000 59.380000 ;
        RECT 64.280000 59.590000 64.480000 59.790000 ;
        RECT 64.280000 60.000000 64.480000 60.200000 ;
        RECT 64.280000 60.410000 64.480000 60.610000 ;
        RECT 64.685000 56.310000 64.885000 56.510000 ;
        RECT 64.685000 56.720000 64.885000 56.920000 ;
        RECT 64.685000 57.130000 64.885000 57.330000 ;
        RECT 64.685000 57.540000 64.885000 57.740000 ;
        RECT 64.685000 57.950000 64.885000 58.150000 ;
        RECT 64.685000 58.360000 64.885000 58.560000 ;
        RECT 64.685000 58.770000 64.885000 58.970000 ;
        RECT 64.685000 59.180000 64.885000 59.380000 ;
        RECT 64.685000 59.590000 64.885000 59.790000 ;
        RECT 64.685000 60.000000 64.885000 60.200000 ;
        RECT 64.685000 60.410000 64.885000 60.610000 ;
        RECT 65.090000 56.310000 65.290000 56.510000 ;
        RECT 65.090000 56.720000 65.290000 56.920000 ;
        RECT 65.090000 57.130000 65.290000 57.330000 ;
        RECT 65.090000 57.540000 65.290000 57.740000 ;
        RECT 65.090000 57.950000 65.290000 58.150000 ;
        RECT 65.090000 58.360000 65.290000 58.560000 ;
        RECT 65.090000 58.770000 65.290000 58.970000 ;
        RECT 65.090000 59.180000 65.290000 59.380000 ;
        RECT 65.090000 59.590000 65.290000 59.790000 ;
        RECT 65.090000 60.000000 65.290000 60.200000 ;
        RECT 65.090000 60.410000 65.290000 60.610000 ;
        RECT 65.495000 56.310000 65.695000 56.510000 ;
        RECT 65.495000 56.720000 65.695000 56.920000 ;
        RECT 65.495000 57.130000 65.695000 57.330000 ;
        RECT 65.495000 57.540000 65.695000 57.740000 ;
        RECT 65.495000 57.950000 65.695000 58.150000 ;
        RECT 65.495000 58.360000 65.695000 58.560000 ;
        RECT 65.495000 58.770000 65.695000 58.970000 ;
        RECT 65.495000 59.180000 65.695000 59.380000 ;
        RECT 65.495000 59.590000 65.695000 59.790000 ;
        RECT 65.495000 60.000000 65.695000 60.200000 ;
        RECT 65.495000 60.410000 65.695000 60.610000 ;
        RECT 65.900000 56.310000 66.100000 56.510000 ;
        RECT 65.900000 56.720000 66.100000 56.920000 ;
        RECT 65.900000 57.130000 66.100000 57.330000 ;
        RECT 65.900000 57.540000 66.100000 57.740000 ;
        RECT 65.900000 57.950000 66.100000 58.150000 ;
        RECT 65.900000 58.360000 66.100000 58.560000 ;
        RECT 65.900000 58.770000 66.100000 58.970000 ;
        RECT 65.900000 59.180000 66.100000 59.380000 ;
        RECT 65.900000 59.590000 66.100000 59.790000 ;
        RECT 65.900000 60.000000 66.100000 60.200000 ;
        RECT 65.900000 60.410000 66.100000 60.610000 ;
        RECT 66.305000 56.310000 66.505000 56.510000 ;
        RECT 66.305000 56.720000 66.505000 56.920000 ;
        RECT 66.305000 57.130000 66.505000 57.330000 ;
        RECT 66.305000 57.540000 66.505000 57.740000 ;
        RECT 66.305000 57.950000 66.505000 58.150000 ;
        RECT 66.305000 58.360000 66.505000 58.560000 ;
        RECT 66.305000 58.770000 66.505000 58.970000 ;
        RECT 66.305000 59.180000 66.505000 59.380000 ;
        RECT 66.305000 59.590000 66.505000 59.790000 ;
        RECT 66.305000 60.000000 66.505000 60.200000 ;
        RECT 66.305000 60.410000 66.505000 60.610000 ;
        RECT 66.710000 56.310000 66.910000 56.510000 ;
        RECT 66.710000 56.720000 66.910000 56.920000 ;
        RECT 66.710000 57.130000 66.910000 57.330000 ;
        RECT 66.710000 57.540000 66.910000 57.740000 ;
        RECT 66.710000 57.950000 66.910000 58.150000 ;
        RECT 66.710000 58.360000 66.910000 58.560000 ;
        RECT 66.710000 58.770000 66.910000 58.970000 ;
        RECT 66.710000 59.180000 66.910000 59.380000 ;
        RECT 66.710000 59.590000 66.910000 59.790000 ;
        RECT 66.710000 60.000000 66.910000 60.200000 ;
        RECT 66.710000 60.410000 66.910000 60.610000 ;
        RECT 67.115000 56.310000 67.315000 56.510000 ;
        RECT 67.115000 56.720000 67.315000 56.920000 ;
        RECT 67.115000 57.130000 67.315000 57.330000 ;
        RECT 67.115000 57.540000 67.315000 57.740000 ;
        RECT 67.115000 57.950000 67.315000 58.150000 ;
        RECT 67.115000 58.360000 67.315000 58.560000 ;
        RECT 67.115000 58.770000 67.315000 58.970000 ;
        RECT 67.115000 59.180000 67.315000 59.380000 ;
        RECT 67.115000 59.590000 67.315000 59.790000 ;
        RECT 67.115000 60.000000 67.315000 60.200000 ;
        RECT 67.115000 60.410000 67.315000 60.610000 ;
        RECT 67.520000 56.310000 67.720000 56.510000 ;
        RECT 67.520000 56.720000 67.720000 56.920000 ;
        RECT 67.520000 57.130000 67.720000 57.330000 ;
        RECT 67.520000 57.540000 67.720000 57.740000 ;
        RECT 67.520000 57.950000 67.720000 58.150000 ;
        RECT 67.520000 58.360000 67.720000 58.560000 ;
        RECT 67.520000 58.770000 67.720000 58.970000 ;
        RECT 67.520000 59.180000 67.720000 59.380000 ;
        RECT 67.520000 59.590000 67.720000 59.790000 ;
        RECT 67.520000 60.000000 67.720000 60.200000 ;
        RECT 67.520000 60.410000 67.720000 60.610000 ;
        RECT 67.925000 56.310000 68.125000 56.510000 ;
        RECT 67.925000 56.720000 68.125000 56.920000 ;
        RECT 67.925000 57.130000 68.125000 57.330000 ;
        RECT 67.925000 57.540000 68.125000 57.740000 ;
        RECT 67.925000 57.950000 68.125000 58.150000 ;
        RECT 67.925000 58.360000 68.125000 58.560000 ;
        RECT 67.925000 58.770000 68.125000 58.970000 ;
        RECT 67.925000 59.180000 68.125000 59.380000 ;
        RECT 67.925000 59.590000 68.125000 59.790000 ;
        RECT 67.925000 60.000000 68.125000 60.200000 ;
        RECT 67.925000 60.410000 68.125000 60.610000 ;
        RECT 68.330000 56.310000 68.530000 56.510000 ;
        RECT 68.330000 56.720000 68.530000 56.920000 ;
        RECT 68.330000 57.130000 68.530000 57.330000 ;
        RECT 68.330000 57.540000 68.530000 57.740000 ;
        RECT 68.330000 57.950000 68.530000 58.150000 ;
        RECT 68.330000 58.360000 68.530000 58.560000 ;
        RECT 68.330000 58.770000 68.530000 58.970000 ;
        RECT 68.330000 59.180000 68.530000 59.380000 ;
        RECT 68.330000 59.590000 68.530000 59.790000 ;
        RECT 68.330000 60.000000 68.530000 60.200000 ;
        RECT 68.330000 60.410000 68.530000 60.610000 ;
        RECT 68.735000 56.310000 68.935000 56.510000 ;
        RECT 68.735000 56.720000 68.935000 56.920000 ;
        RECT 68.735000 57.130000 68.935000 57.330000 ;
        RECT 68.735000 57.540000 68.935000 57.740000 ;
        RECT 68.735000 57.950000 68.935000 58.150000 ;
        RECT 68.735000 58.360000 68.935000 58.560000 ;
        RECT 68.735000 58.770000 68.935000 58.970000 ;
        RECT 68.735000 59.180000 68.935000 59.380000 ;
        RECT 68.735000 59.590000 68.935000 59.790000 ;
        RECT 68.735000 60.000000 68.935000 60.200000 ;
        RECT 68.735000 60.410000 68.935000 60.610000 ;
        RECT 69.140000 56.310000 69.340000 56.510000 ;
        RECT 69.140000 56.720000 69.340000 56.920000 ;
        RECT 69.140000 57.130000 69.340000 57.330000 ;
        RECT 69.140000 57.540000 69.340000 57.740000 ;
        RECT 69.140000 57.950000 69.340000 58.150000 ;
        RECT 69.140000 58.360000 69.340000 58.560000 ;
        RECT 69.140000 58.770000 69.340000 58.970000 ;
        RECT 69.140000 59.180000 69.340000 59.380000 ;
        RECT 69.140000 59.590000 69.340000 59.790000 ;
        RECT 69.140000 60.000000 69.340000 60.200000 ;
        RECT 69.140000 60.410000 69.340000 60.610000 ;
        RECT 69.545000 56.310000 69.745000 56.510000 ;
        RECT 69.545000 56.720000 69.745000 56.920000 ;
        RECT 69.545000 57.130000 69.745000 57.330000 ;
        RECT 69.545000 57.540000 69.745000 57.740000 ;
        RECT 69.545000 57.950000 69.745000 58.150000 ;
        RECT 69.545000 58.360000 69.745000 58.560000 ;
        RECT 69.545000 58.770000 69.745000 58.970000 ;
        RECT 69.545000 59.180000 69.745000 59.380000 ;
        RECT 69.545000 59.590000 69.745000 59.790000 ;
        RECT 69.545000 60.000000 69.745000 60.200000 ;
        RECT 69.545000 60.410000 69.745000 60.610000 ;
        RECT 69.950000 56.310000 70.150000 56.510000 ;
        RECT 69.950000 56.720000 70.150000 56.920000 ;
        RECT 69.950000 57.130000 70.150000 57.330000 ;
        RECT 69.950000 57.540000 70.150000 57.740000 ;
        RECT 69.950000 57.950000 70.150000 58.150000 ;
        RECT 69.950000 58.360000 70.150000 58.560000 ;
        RECT 69.950000 58.770000 70.150000 58.970000 ;
        RECT 69.950000 59.180000 70.150000 59.380000 ;
        RECT 69.950000 59.590000 70.150000 59.790000 ;
        RECT 69.950000 60.000000 70.150000 60.200000 ;
        RECT 69.950000 60.410000 70.150000 60.610000 ;
        RECT 70.355000 56.310000 70.555000 56.510000 ;
        RECT 70.355000 56.720000 70.555000 56.920000 ;
        RECT 70.355000 57.130000 70.555000 57.330000 ;
        RECT 70.355000 57.540000 70.555000 57.740000 ;
        RECT 70.355000 57.950000 70.555000 58.150000 ;
        RECT 70.355000 58.360000 70.555000 58.560000 ;
        RECT 70.355000 58.770000 70.555000 58.970000 ;
        RECT 70.355000 59.180000 70.555000 59.380000 ;
        RECT 70.355000 59.590000 70.555000 59.790000 ;
        RECT 70.355000 60.000000 70.555000 60.200000 ;
        RECT 70.355000 60.410000 70.555000 60.610000 ;
        RECT 70.760000 56.310000 70.960000 56.510000 ;
        RECT 70.760000 56.720000 70.960000 56.920000 ;
        RECT 70.760000 57.130000 70.960000 57.330000 ;
        RECT 70.760000 57.540000 70.960000 57.740000 ;
        RECT 70.760000 57.950000 70.960000 58.150000 ;
        RECT 70.760000 58.360000 70.960000 58.560000 ;
        RECT 70.760000 58.770000 70.960000 58.970000 ;
        RECT 70.760000 59.180000 70.960000 59.380000 ;
        RECT 70.760000 59.590000 70.960000 59.790000 ;
        RECT 70.760000 60.000000 70.960000 60.200000 ;
        RECT 70.760000 60.410000 70.960000 60.610000 ;
        RECT 71.165000 56.310000 71.365000 56.510000 ;
        RECT 71.165000 56.720000 71.365000 56.920000 ;
        RECT 71.165000 57.130000 71.365000 57.330000 ;
        RECT 71.165000 57.540000 71.365000 57.740000 ;
        RECT 71.165000 57.950000 71.365000 58.150000 ;
        RECT 71.165000 58.360000 71.365000 58.560000 ;
        RECT 71.165000 58.770000 71.365000 58.970000 ;
        RECT 71.165000 59.180000 71.365000 59.380000 ;
        RECT 71.165000 59.590000 71.365000 59.790000 ;
        RECT 71.165000 60.000000 71.365000 60.200000 ;
        RECT 71.165000 60.410000 71.365000 60.610000 ;
        RECT 71.570000 56.310000 71.770000 56.510000 ;
        RECT 71.570000 56.720000 71.770000 56.920000 ;
        RECT 71.570000 57.130000 71.770000 57.330000 ;
        RECT 71.570000 57.540000 71.770000 57.740000 ;
        RECT 71.570000 57.950000 71.770000 58.150000 ;
        RECT 71.570000 58.360000 71.770000 58.560000 ;
        RECT 71.570000 58.770000 71.770000 58.970000 ;
        RECT 71.570000 59.180000 71.770000 59.380000 ;
        RECT 71.570000 59.590000 71.770000 59.790000 ;
        RECT 71.570000 60.000000 71.770000 60.200000 ;
        RECT 71.570000 60.410000 71.770000 60.610000 ;
        RECT 71.975000 56.310000 72.175000 56.510000 ;
        RECT 71.975000 56.720000 72.175000 56.920000 ;
        RECT 71.975000 57.130000 72.175000 57.330000 ;
        RECT 71.975000 57.540000 72.175000 57.740000 ;
        RECT 71.975000 57.950000 72.175000 58.150000 ;
        RECT 71.975000 58.360000 72.175000 58.560000 ;
        RECT 71.975000 58.770000 72.175000 58.970000 ;
        RECT 71.975000 59.180000 72.175000 59.380000 ;
        RECT 71.975000 59.590000 72.175000 59.790000 ;
        RECT 71.975000 60.000000 72.175000 60.200000 ;
        RECT 71.975000 60.410000 72.175000 60.610000 ;
        RECT 72.380000 56.310000 72.580000 56.510000 ;
        RECT 72.380000 56.720000 72.580000 56.920000 ;
        RECT 72.380000 57.130000 72.580000 57.330000 ;
        RECT 72.380000 57.540000 72.580000 57.740000 ;
        RECT 72.380000 57.950000 72.580000 58.150000 ;
        RECT 72.380000 58.360000 72.580000 58.560000 ;
        RECT 72.380000 58.770000 72.580000 58.970000 ;
        RECT 72.380000 59.180000 72.580000 59.380000 ;
        RECT 72.380000 59.590000 72.580000 59.790000 ;
        RECT 72.380000 60.000000 72.580000 60.200000 ;
        RECT 72.380000 60.410000 72.580000 60.610000 ;
        RECT 72.785000 56.310000 72.985000 56.510000 ;
        RECT 72.785000 56.720000 72.985000 56.920000 ;
        RECT 72.785000 57.130000 72.985000 57.330000 ;
        RECT 72.785000 57.540000 72.985000 57.740000 ;
        RECT 72.785000 57.950000 72.985000 58.150000 ;
        RECT 72.785000 58.360000 72.985000 58.560000 ;
        RECT 72.785000 58.770000 72.985000 58.970000 ;
        RECT 72.785000 59.180000 72.985000 59.380000 ;
        RECT 72.785000 59.590000 72.985000 59.790000 ;
        RECT 72.785000 60.000000 72.985000 60.200000 ;
        RECT 72.785000 60.410000 72.985000 60.610000 ;
        RECT 73.190000 56.310000 73.390000 56.510000 ;
        RECT 73.190000 56.720000 73.390000 56.920000 ;
        RECT 73.190000 57.130000 73.390000 57.330000 ;
        RECT 73.190000 57.540000 73.390000 57.740000 ;
        RECT 73.190000 57.950000 73.390000 58.150000 ;
        RECT 73.190000 58.360000 73.390000 58.560000 ;
        RECT 73.190000 58.770000 73.390000 58.970000 ;
        RECT 73.190000 59.180000 73.390000 59.380000 ;
        RECT 73.190000 59.590000 73.390000 59.790000 ;
        RECT 73.190000 60.000000 73.390000 60.200000 ;
        RECT 73.190000 60.410000 73.390000 60.610000 ;
        RECT 73.595000 56.310000 73.795000 56.510000 ;
        RECT 73.595000 56.720000 73.795000 56.920000 ;
        RECT 73.595000 57.130000 73.795000 57.330000 ;
        RECT 73.595000 57.540000 73.795000 57.740000 ;
        RECT 73.595000 57.950000 73.795000 58.150000 ;
        RECT 73.595000 58.360000 73.795000 58.560000 ;
        RECT 73.595000 58.770000 73.795000 58.970000 ;
        RECT 73.595000 59.180000 73.795000 59.380000 ;
        RECT 73.595000 59.590000 73.795000 59.790000 ;
        RECT 73.595000 60.000000 73.795000 60.200000 ;
        RECT 73.595000 60.410000 73.795000 60.610000 ;
        RECT 74.000000 56.310000 74.200000 56.510000 ;
        RECT 74.000000 56.720000 74.200000 56.920000 ;
        RECT 74.000000 57.130000 74.200000 57.330000 ;
        RECT 74.000000 57.540000 74.200000 57.740000 ;
        RECT 74.000000 57.950000 74.200000 58.150000 ;
        RECT 74.000000 58.360000 74.200000 58.560000 ;
        RECT 74.000000 58.770000 74.200000 58.970000 ;
        RECT 74.000000 59.180000 74.200000 59.380000 ;
        RECT 74.000000 59.590000 74.200000 59.790000 ;
        RECT 74.000000 60.000000 74.200000 60.200000 ;
        RECT 74.000000 60.410000 74.200000 60.610000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000 75.000000  23.440000 ;
      RECT  0.000000  28.880000 75.000000  55.840000 ;
      RECT  0.000000  61.080000 75.000000 170.795000 ;
      RECT 13.300000 170.795000 61.645000 198.000000 ;
      RECT 24.800000  23.440000 50.355000  28.880000 ;
      RECT 24.800000  55.840000 50.355000  61.080000 ;
      RECT 74.690000  23.440000 75.000000  28.880000 ;
      RECT 74.690000  55.840000 75.000000  61.080000 ;
    LAYER met4 ;
      RECT  0.000000   5.885000  1.670000   6.485000 ;
      RECT  0.000000  11.935000  1.365000  12.535000 ;
      RECT  0.000000  16.785000  1.365000  17.385000 ;
      RECT  0.000000  22.835000  1.670000  23.435000 ;
      RECT  0.000000  28.885000  1.670000  29.485000 ;
      RECT  0.000000  33.735000  1.670000  34.335000 ;
      RECT  0.000000  38.585000  1.670000  39.185000 ;
      RECT  0.000000  44.635000  1.670000  45.335000 ;
      RECT  0.000000  55.135000  1.670000  55.835000 ;
      RECT  0.000000  61.085000  1.670000  61.685000 ;
      RECT  0.000000  66.935000  1.670000  67.635000 ;
      RECT  0.000000  93.400000 75.000000 173.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.670000   0.000000 73.330000  11.935000 ;
      RECT  1.670000   0.000000 73.330000  23.435000 ;
      RECT  1.670000   0.000000 73.330000  23.435000 ;
      RECT  1.670000   0.000000 73.330000  23.435000 ;
      RECT  1.670000  17.385000 73.330000  23.435000 ;
      RECT  1.670000  28.885000 73.330000  55.835000 ;
      RECT  1.670000  28.885000 73.330000  55.835000 ;
      RECT  1.670000  28.885000 73.330000  55.835000 ;
      RECT  1.670000  28.885000 73.330000  55.835000 ;
      RECT  1.670000  28.885000 73.330000  55.835000 ;
      RECT  1.670000  61.085000 73.330000  93.400000 ;
      RECT  1.670000  61.085000 73.330000 173.435000 ;
      RECT  1.670000  61.085000 73.330000 173.435000 ;
      RECT  1.670000  61.085000 73.330000 173.435000 ;
      RECT  1.670000 173.385000 73.330000 173.435000 ;
      RECT 13.300000  61.085000 61.675000 198.000000 ;
      RECT 13.300000 173.435000 61.675000 198.000000 ;
      RECT 24.775000   0.000000 50.380000  61.085000 ;
      RECT 24.775000   0.000000 50.380000 198.000000 ;
      RECT 24.775000  23.435000 50.380000  28.885000 ;
      RECT 24.775000  55.835000 50.380000  61.085000 ;
      RECT 73.330000   5.885000 75.000000   6.485000 ;
      RECT 73.330000  22.835000 75.000000  23.435000 ;
      RECT 73.330000  28.885000 75.000000  29.485000 ;
      RECT 73.330000  33.735000 75.000000  34.335000 ;
      RECT 73.330000  38.585000 75.000000  39.185000 ;
      RECT 73.330000  44.635000 75.000000  45.335000 ;
      RECT 73.330000  55.135000 75.000000  55.835000 ;
      RECT 73.330000  61.085000 75.000000  61.685000 ;
      RECT 73.330000  66.935000 75.000000  67.635000 ;
      RECT 73.635000  11.935000 75.000000  12.535000 ;
      RECT 73.635000  16.785000 75.000000  17.385000 ;
    LAYER met5 ;
      RECT 0.000000  93.785000 75.000000 172.985000 ;
      RECT 1.765000  12.235000 73.235000  17.085000 ;
      RECT 2.070000   0.000000 72.930000  12.235000 ;
      RECT 2.070000  17.085000 72.930000  93.785000 ;
      RECT 2.070000 172.985000 72.930000 198.000000 ;
  END
END sky130_fd_io__overlay_vssio_lvc


MACRO sky130_fd_io__overlay_vddio_lvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.595000 68.035000 24.495000 82.665000 ;
        RECT 0.595000 82.665000 24.345000 82.815000 ;
        RECT 0.595000 82.815000 24.195000 82.965000 ;
        RECT 0.595000 82.965000 24.045000 83.115000 ;
        RECT 0.595000 83.115000 23.895000 83.265000 ;
        RECT 0.595000 83.265000 23.745000 83.415000 ;
        RECT 0.595000 83.415000 23.595000 83.565000 ;
        RECT 0.595000 83.565000 23.445000 83.715000 ;
        RECT 0.595000 83.715000 23.295000 83.865000 ;
        RECT 0.595000 83.865000 23.145000 84.015000 ;
        RECT 0.595000 84.015000 22.995000 84.165000 ;
        RECT 0.595000 84.165000 22.845000 84.315000 ;
        RECT 0.595000 84.315000 22.695000 84.465000 ;
        RECT 0.595000 84.465000 22.545000 84.615000 ;
        RECT 0.595000 84.615000 22.395000 84.765000 ;
        RECT 0.595000 84.765000 22.245000 84.915000 ;
        RECT 0.595000 84.915000 22.095000 85.065000 ;
        RECT 0.595000 85.065000 21.945000 85.215000 ;
        RECT 0.595000 85.215000 21.795000 85.365000 ;
        RECT 0.595000 85.365000 21.645000 85.515000 ;
        RECT 0.595000 85.515000 21.495000 85.665000 ;
        RECT 0.595000 85.665000 21.345000 85.815000 ;
        RECT 0.595000 85.815000 21.195000 85.965000 ;
        RECT 0.595000 85.965000 21.045000 86.115000 ;
        RECT 0.595000 86.115000 20.895000 86.265000 ;
        RECT 0.595000 86.265000 20.745000 86.415000 ;
        RECT 0.595000 86.415000 20.595000 86.565000 ;
        RECT 0.595000 86.565000 20.445000 86.715000 ;
        RECT 0.595000 86.715000 20.295000 86.865000 ;
        RECT 0.595000 86.865000 20.145000 87.015000 ;
        RECT 0.595000 87.015000 19.995000 87.165000 ;
        RECT 0.595000 87.165000 19.845000 87.315000 ;
        RECT 0.595000 87.315000 19.695000 87.465000 ;
        RECT 0.595000 87.465000 19.545000 87.615000 ;
        RECT 0.595000 87.615000 19.395000 87.765000 ;
        RECT 0.595000 87.765000 19.245000 87.915000 ;
        RECT 0.595000 87.915000 19.095000 88.065000 ;
        RECT 0.595000 88.065000 18.945000 88.215000 ;
        RECT 0.595000 88.215000 18.795000 88.365000 ;
        RECT 0.595000 88.365000 18.645000 88.515000 ;
        RECT 0.595000 88.515000 18.495000 88.665000 ;
        RECT 0.595000 88.665000 18.345000 88.815000 ;
        RECT 0.595000 88.815000 18.195000 88.965000 ;
        RECT 0.595000 88.965000 18.045000 89.115000 ;
        RECT 0.595000 89.115000 17.895000 89.265000 ;
        RECT 0.595000 89.265000 17.745000 89.415000 ;
        RECT 0.595000 89.415000 17.595000 89.565000 ;
        RECT 0.595000 89.565000 17.445000 89.715000 ;
        RECT 0.595000 89.715000 17.295000 89.865000 ;
        RECT 0.595000 89.865000 17.145000 90.015000 ;
        RECT 0.595000 90.015000 16.995000 90.165000 ;
        RECT 0.595000 90.165000 16.845000 90.315000 ;
        RECT 0.595000 90.315000 16.695000 90.465000 ;
        RECT 0.595000 90.465000 16.545000 90.615000 ;
        RECT 0.595000 90.615000 16.395000 90.765000 ;
        RECT 0.595000 90.765000 16.245000 90.915000 ;
        RECT 0.595000 90.915000 16.095000 91.065000 ;
        RECT 0.595000 91.065000 15.945000 91.215000 ;
        RECT 0.595000 91.215000 15.795000 91.365000 ;
        RECT 0.595000 91.365000 15.645000 91.515000 ;
        RECT 0.595000 91.515000 15.495000 91.665000 ;
        RECT 0.595000 91.665000 15.345000 91.815000 ;
        RECT 0.595000 91.815000 15.195000 91.965000 ;
        RECT 0.595000 91.965000 15.045000 92.115000 ;
        RECT 0.595000 92.115000 14.895000 92.265000 ;
        RECT 0.595000 92.265000 14.745000 92.415000 ;
        RECT 0.595000 92.415000 14.595000 92.565000 ;
        RECT 0.595000 92.565000 14.445000 92.715000 ;
        RECT 0.595000 92.715000 14.295000 92.865000 ;
        RECT 0.595000 92.865000 14.205000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.600000 17.790000 24.500000 22.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 17.790000 74.655000 22.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.760000 68.035000 74.660000 82.665000 ;
        RECT 50.910000 82.665000 74.660000 82.815000 ;
        RECT 51.060000 82.815000 74.660000 82.965000 ;
        RECT 51.210000 82.965000 74.660000 83.115000 ;
        RECT 51.360000 83.115000 74.660000 83.265000 ;
        RECT 51.510000 83.265000 74.660000 83.415000 ;
        RECT 51.660000 83.415000 74.660000 83.565000 ;
        RECT 51.810000 83.565000 74.660000 83.715000 ;
        RECT 51.960000 83.715000 74.660000 83.865000 ;
        RECT 52.110000 83.865000 74.660000 84.015000 ;
        RECT 52.260000 84.015000 74.660000 84.165000 ;
        RECT 52.410000 84.165000 74.660000 84.315000 ;
        RECT 52.560000 84.315000 74.660000 84.465000 ;
        RECT 52.710000 84.465000 74.660000 84.615000 ;
        RECT 52.860000 84.615000 74.660000 84.765000 ;
        RECT 53.010000 84.765000 74.660000 84.915000 ;
        RECT 53.160000 84.915000 74.660000 85.065000 ;
        RECT 53.310000 85.065000 74.660000 85.215000 ;
        RECT 53.460000 85.215000 74.660000 85.365000 ;
        RECT 53.610000 85.365000 74.660000 85.515000 ;
        RECT 53.760000 85.515000 74.660000 85.665000 ;
        RECT 53.910000 85.665000 74.660000 85.815000 ;
        RECT 54.060000 85.815000 74.660000 85.965000 ;
        RECT 54.210000 85.965000 74.660000 86.115000 ;
        RECT 54.360000 86.115000 74.660000 86.265000 ;
        RECT 54.510000 86.265000 74.660000 86.415000 ;
        RECT 54.660000 86.415000 74.660000 86.565000 ;
        RECT 54.810000 86.565000 74.660000 86.715000 ;
        RECT 54.960000 86.715000 74.660000 86.865000 ;
        RECT 55.110000 86.865000 74.660000 87.015000 ;
        RECT 55.260000 87.015000 74.660000 87.165000 ;
        RECT 55.410000 87.165000 74.660000 87.315000 ;
        RECT 55.560000 87.315000 74.660000 87.465000 ;
        RECT 55.710000 87.465000 74.660000 87.615000 ;
        RECT 55.860000 87.615000 74.660000 87.765000 ;
        RECT 56.010000 87.765000 74.660000 87.915000 ;
        RECT 56.160000 87.915000 74.660000 88.065000 ;
        RECT 56.310000 88.065000 74.660000 88.215000 ;
        RECT 56.460000 88.215000 74.660000 88.365000 ;
        RECT 56.610000 88.365000 74.660000 88.515000 ;
        RECT 56.760000 88.515000 74.660000 88.665000 ;
        RECT 56.910000 88.665000 74.660000 88.815000 ;
        RECT 57.060000 88.815000 74.660000 88.965000 ;
        RECT 57.210000 88.965000 74.660000 89.115000 ;
        RECT 57.360000 89.115000 74.660000 89.265000 ;
        RECT 57.510000 89.265000 74.660000 89.415000 ;
        RECT 57.660000 89.415000 74.660000 89.565000 ;
        RECT 57.810000 89.565000 74.660000 89.715000 ;
        RECT 57.960000 89.715000 74.660000 89.865000 ;
        RECT 58.110000 89.865000 74.660000 90.015000 ;
        RECT 58.260000 90.015000 74.660000 90.165000 ;
        RECT 58.410000 90.165000 74.660000 90.315000 ;
        RECT 58.560000 90.315000 74.660000 90.465000 ;
        RECT 58.710000 90.465000 74.660000 90.615000 ;
        RECT 58.860000 90.615000 74.660000 90.765000 ;
        RECT 59.010000 90.765000 74.660000 90.915000 ;
        RECT 59.160000 90.915000 74.660000 91.065000 ;
        RECT 59.310000 91.065000 74.660000 91.215000 ;
        RECT 59.460000 91.215000 74.660000 91.365000 ;
        RECT 59.610000 91.365000 74.660000 91.515000 ;
        RECT 59.760000 91.515000 74.660000 91.665000 ;
        RECT 59.910000 91.665000 74.660000 91.815000 ;
        RECT 60.060000 91.815000 74.660000 91.965000 ;
        RECT 60.210000 91.965000 74.660000 92.115000 ;
        RECT 60.360000 92.115000 74.660000 92.265000 ;
        RECT 60.510000 92.265000 74.660000 92.415000 ;
        RECT 60.660000 92.415000 74.660000 92.565000 ;
        RECT 60.810000 92.565000 74.660000 92.715000 ;
        RECT 60.960000 92.715000 74.660000 92.865000 ;
        RECT 61.055000 92.865000 74.660000 92.960000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 24.475000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000  1.270000 68.060000 ;
        RECT 0.000000 68.060000 24.500000 82.625000 ;
        RECT 0.000000 82.625000  1.270000 82.790000 ;
        RECT 0.000000 82.790000 14.105000 92.960000 ;
        RECT 0.000000 92.960000  1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.255000 90.950000 15.365000 91.710000 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.270000 88.345000 16.250000 90.820000 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.375000 82.990000 18.855000 88.140000 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.415000 88.365000 17.525000 89.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 18.995000 85.810000 20.065000 87.015000 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.170000 82.945000 21.450000 85.590000 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.650000 82.855000 22.770000 84.285000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.755000 68.060000 75.000000 82.625000 ;
        RECT 61.150000 82.785000 75.000000 92.965000 ;
        RECT 73.730000 68.035000 75.000000 68.060000 ;
        RECT 73.730000 82.625000 75.000000 82.785000 ;
        RECT 73.730000 92.965000 75.000000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 52.485000 82.855000 53.605000 84.285000 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.805000 82.945000 56.085000 85.590000 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.190000 85.810000 56.260000 87.015000 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.400000 82.990000 60.880000 88.140000 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.730000 88.365000 58.840000 89.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.005000 88.345000 60.985000 90.820000 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.890000 90.950000 61.000000 91.710000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.690000 17.860000  0.890000 18.060000 ;
        RECT  0.690000 18.290000  0.890000 18.490000 ;
        RECT  0.690000 18.720000  0.890000 18.920000 ;
        RECT  0.690000 19.150000  0.890000 19.350000 ;
        RECT  0.690000 19.580000  0.890000 19.780000 ;
        RECT  0.690000 20.010000  0.890000 20.210000 ;
        RECT  0.690000 20.440000  0.890000 20.640000 ;
        RECT  0.690000 20.870000  0.890000 21.070000 ;
        RECT  0.690000 21.300000  0.890000 21.500000 ;
        RECT  0.690000 21.730000  0.890000 21.930000 ;
        RECT  0.690000 22.160000  0.890000 22.360000 ;
        RECT  0.735000 82.855000  0.935000 83.055000 ;
        RECT  0.735000 83.265000  0.935000 83.465000 ;
        RECT  0.735000 83.675000  0.935000 83.875000 ;
        RECT  0.735000 84.085000  0.935000 84.285000 ;
        RECT  0.735000 84.495000  0.935000 84.695000 ;
        RECT  0.735000 84.905000  0.935000 85.105000 ;
        RECT  0.735000 85.315000  0.935000 85.515000 ;
        RECT  0.735000 85.725000  0.935000 85.925000 ;
        RECT  0.735000 86.135000  0.935000 86.335000 ;
        RECT  0.735000 86.545000  0.935000 86.745000 ;
        RECT  0.735000 86.955000  0.935000 87.155000 ;
        RECT  0.735000 87.365000  0.935000 87.565000 ;
        RECT  0.735000 87.775000  0.935000 87.975000 ;
        RECT  0.735000 88.185000  0.935000 88.385000 ;
        RECT  0.735000 88.595000  0.935000 88.795000 ;
        RECT  0.735000 89.005000  0.935000 89.205000 ;
        RECT  0.735000 89.415000  0.935000 89.615000 ;
        RECT  0.735000 89.825000  0.935000 90.025000 ;
        RECT  0.735000 90.235000  0.935000 90.435000 ;
        RECT  0.735000 90.645000  0.935000 90.845000 ;
        RECT  0.735000 91.055000  0.935000 91.255000 ;
        RECT  0.735000 91.465000  0.935000 91.665000 ;
        RECT  0.735000 91.875000  0.935000 92.075000 ;
        RECT  0.735000 92.285000  0.935000 92.485000 ;
        RECT  0.735000 92.695000  0.935000 92.895000 ;
        RECT  0.845000 68.125000  1.045000 68.325000 ;
        RECT  0.845000 68.535000  1.045000 68.735000 ;
        RECT  0.845000 68.945000  1.045000 69.145000 ;
        RECT  0.845000 69.355000  1.045000 69.555000 ;
        RECT  0.845000 69.765000  1.045000 69.965000 ;
        RECT  0.845000 70.175000  1.045000 70.375000 ;
        RECT  0.845000 70.585000  1.045000 70.785000 ;
        RECT  0.845000 70.995000  1.045000 71.195000 ;
        RECT  0.845000 71.405000  1.045000 71.605000 ;
        RECT  0.845000 71.815000  1.045000 72.015000 ;
        RECT  0.845000 72.225000  1.045000 72.425000 ;
        RECT  0.845000 72.635000  1.045000 72.835000 ;
        RECT  0.845000 73.045000  1.045000 73.245000 ;
        RECT  0.845000 73.450000  1.045000 73.650000 ;
        RECT  0.845000 73.855000  1.045000 74.055000 ;
        RECT  0.845000 74.260000  1.045000 74.460000 ;
        RECT  0.845000 74.665000  1.045000 74.865000 ;
        RECT  0.845000 75.070000  1.045000 75.270000 ;
        RECT  0.845000 75.475000  1.045000 75.675000 ;
        RECT  0.845000 75.880000  1.045000 76.080000 ;
        RECT  0.845000 76.285000  1.045000 76.485000 ;
        RECT  0.845000 76.690000  1.045000 76.890000 ;
        RECT  0.845000 77.095000  1.045000 77.295000 ;
        RECT  0.845000 77.500000  1.045000 77.700000 ;
        RECT  0.845000 77.905000  1.045000 78.105000 ;
        RECT  0.845000 78.310000  1.045000 78.510000 ;
        RECT  0.845000 78.715000  1.045000 78.915000 ;
        RECT  0.845000 79.120000  1.045000 79.320000 ;
        RECT  0.845000 79.525000  1.045000 79.725000 ;
        RECT  0.845000 79.930000  1.045000 80.130000 ;
        RECT  0.845000 80.335000  1.045000 80.535000 ;
        RECT  0.845000 80.740000  1.045000 80.940000 ;
        RECT  0.845000 81.145000  1.045000 81.345000 ;
        RECT  0.845000 81.550000  1.045000 81.750000 ;
        RECT  0.845000 81.955000  1.045000 82.155000 ;
        RECT  0.845000 82.360000  1.045000 82.560000 ;
        RECT  1.095000 17.860000  1.295000 18.060000 ;
        RECT  1.095000 18.290000  1.295000 18.490000 ;
        RECT  1.095000 18.720000  1.295000 18.920000 ;
        RECT  1.095000 19.150000  1.295000 19.350000 ;
        RECT  1.095000 19.580000  1.295000 19.780000 ;
        RECT  1.095000 20.010000  1.295000 20.210000 ;
        RECT  1.095000 20.440000  1.295000 20.640000 ;
        RECT  1.095000 20.870000  1.295000 21.070000 ;
        RECT  1.095000 21.300000  1.295000 21.500000 ;
        RECT  1.095000 21.730000  1.295000 21.930000 ;
        RECT  1.095000 22.160000  1.295000 22.360000 ;
        RECT  1.145000 82.855000  1.345000 83.055000 ;
        RECT  1.145000 83.265000  1.345000 83.465000 ;
        RECT  1.145000 83.675000  1.345000 83.875000 ;
        RECT  1.145000 84.085000  1.345000 84.285000 ;
        RECT  1.145000 84.495000  1.345000 84.695000 ;
        RECT  1.145000 84.905000  1.345000 85.105000 ;
        RECT  1.145000 85.315000  1.345000 85.515000 ;
        RECT  1.145000 85.725000  1.345000 85.925000 ;
        RECT  1.145000 86.135000  1.345000 86.335000 ;
        RECT  1.145000 86.545000  1.345000 86.745000 ;
        RECT  1.145000 86.955000  1.345000 87.155000 ;
        RECT  1.145000 87.365000  1.345000 87.565000 ;
        RECT  1.145000 87.775000  1.345000 87.975000 ;
        RECT  1.145000 88.185000  1.345000 88.385000 ;
        RECT  1.145000 88.595000  1.345000 88.795000 ;
        RECT  1.145000 89.005000  1.345000 89.205000 ;
        RECT  1.145000 89.415000  1.345000 89.615000 ;
        RECT  1.145000 89.825000  1.345000 90.025000 ;
        RECT  1.145000 90.235000  1.345000 90.435000 ;
        RECT  1.145000 90.645000  1.345000 90.845000 ;
        RECT  1.145000 91.055000  1.345000 91.255000 ;
        RECT  1.145000 91.465000  1.345000 91.665000 ;
        RECT  1.145000 91.875000  1.345000 92.075000 ;
        RECT  1.145000 92.285000  1.345000 92.485000 ;
        RECT  1.145000 92.695000  1.345000 92.895000 ;
        RECT  1.245000 68.125000  1.445000 68.325000 ;
        RECT  1.245000 68.535000  1.445000 68.735000 ;
        RECT  1.245000 68.945000  1.445000 69.145000 ;
        RECT  1.245000 69.355000  1.445000 69.555000 ;
        RECT  1.245000 69.765000  1.445000 69.965000 ;
        RECT  1.245000 70.175000  1.445000 70.375000 ;
        RECT  1.245000 70.585000  1.445000 70.785000 ;
        RECT  1.245000 70.995000  1.445000 71.195000 ;
        RECT  1.245000 71.405000  1.445000 71.605000 ;
        RECT  1.245000 71.815000  1.445000 72.015000 ;
        RECT  1.245000 72.225000  1.445000 72.425000 ;
        RECT  1.245000 72.635000  1.445000 72.835000 ;
        RECT  1.245000 73.045000  1.445000 73.245000 ;
        RECT  1.245000 73.450000  1.445000 73.650000 ;
        RECT  1.245000 73.855000  1.445000 74.055000 ;
        RECT  1.245000 74.260000  1.445000 74.460000 ;
        RECT  1.245000 74.665000  1.445000 74.865000 ;
        RECT  1.245000 75.070000  1.445000 75.270000 ;
        RECT  1.245000 75.475000  1.445000 75.675000 ;
        RECT  1.245000 75.880000  1.445000 76.080000 ;
        RECT  1.245000 76.285000  1.445000 76.485000 ;
        RECT  1.245000 76.690000  1.445000 76.890000 ;
        RECT  1.245000 77.095000  1.445000 77.295000 ;
        RECT  1.245000 77.500000  1.445000 77.700000 ;
        RECT  1.245000 77.905000  1.445000 78.105000 ;
        RECT  1.245000 78.310000  1.445000 78.510000 ;
        RECT  1.245000 78.715000  1.445000 78.915000 ;
        RECT  1.245000 79.120000  1.445000 79.320000 ;
        RECT  1.245000 79.525000  1.445000 79.725000 ;
        RECT  1.245000 79.930000  1.445000 80.130000 ;
        RECT  1.245000 80.335000  1.445000 80.535000 ;
        RECT  1.245000 80.740000  1.445000 80.940000 ;
        RECT  1.245000 81.145000  1.445000 81.345000 ;
        RECT  1.245000 81.550000  1.445000 81.750000 ;
        RECT  1.245000 81.955000  1.445000 82.155000 ;
        RECT  1.245000 82.360000  1.445000 82.560000 ;
        RECT  1.500000 17.860000  1.700000 18.060000 ;
        RECT  1.500000 18.290000  1.700000 18.490000 ;
        RECT  1.500000 18.720000  1.700000 18.920000 ;
        RECT  1.500000 19.150000  1.700000 19.350000 ;
        RECT  1.500000 19.580000  1.700000 19.780000 ;
        RECT  1.500000 20.010000  1.700000 20.210000 ;
        RECT  1.500000 20.440000  1.700000 20.640000 ;
        RECT  1.500000 20.870000  1.700000 21.070000 ;
        RECT  1.500000 21.300000  1.700000 21.500000 ;
        RECT  1.500000 21.730000  1.700000 21.930000 ;
        RECT  1.500000 22.160000  1.700000 22.360000 ;
        RECT  1.555000 82.855000  1.755000 83.055000 ;
        RECT  1.555000 83.265000  1.755000 83.465000 ;
        RECT  1.555000 83.675000  1.755000 83.875000 ;
        RECT  1.555000 84.085000  1.755000 84.285000 ;
        RECT  1.555000 84.495000  1.755000 84.695000 ;
        RECT  1.555000 84.905000  1.755000 85.105000 ;
        RECT  1.555000 85.315000  1.755000 85.515000 ;
        RECT  1.555000 85.725000  1.755000 85.925000 ;
        RECT  1.555000 86.135000  1.755000 86.335000 ;
        RECT  1.555000 86.545000  1.755000 86.745000 ;
        RECT  1.555000 86.955000  1.755000 87.155000 ;
        RECT  1.555000 87.365000  1.755000 87.565000 ;
        RECT  1.555000 87.775000  1.755000 87.975000 ;
        RECT  1.555000 88.185000  1.755000 88.385000 ;
        RECT  1.555000 88.595000  1.755000 88.795000 ;
        RECT  1.555000 89.005000  1.755000 89.205000 ;
        RECT  1.555000 89.415000  1.755000 89.615000 ;
        RECT  1.555000 89.825000  1.755000 90.025000 ;
        RECT  1.555000 90.235000  1.755000 90.435000 ;
        RECT  1.555000 90.645000  1.755000 90.845000 ;
        RECT  1.555000 91.055000  1.755000 91.255000 ;
        RECT  1.555000 91.465000  1.755000 91.665000 ;
        RECT  1.555000 91.875000  1.755000 92.075000 ;
        RECT  1.555000 92.285000  1.755000 92.485000 ;
        RECT  1.555000 92.695000  1.755000 92.895000 ;
        RECT  1.645000 68.125000  1.845000 68.325000 ;
        RECT  1.645000 68.535000  1.845000 68.735000 ;
        RECT  1.645000 68.945000  1.845000 69.145000 ;
        RECT  1.645000 69.355000  1.845000 69.555000 ;
        RECT  1.645000 69.765000  1.845000 69.965000 ;
        RECT  1.645000 70.175000  1.845000 70.375000 ;
        RECT  1.645000 70.585000  1.845000 70.785000 ;
        RECT  1.645000 70.995000  1.845000 71.195000 ;
        RECT  1.645000 71.405000  1.845000 71.605000 ;
        RECT  1.645000 71.815000  1.845000 72.015000 ;
        RECT  1.645000 72.225000  1.845000 72.425000 ;
        RECT  1.645000 72.635000  1.845000 72.835000 ;
        RECT  1.645000 73.045000  1.845000 73.245000 ;
        RECT  1.645000 73.450000  1.845000 73.650000 ;
        RECT  1.645000 73.855000  1.845000 74.055000 ;
        RECT  1.645000 74.260000  1.845000 74.460000 ;
        RECT  1.645000 74.665000  1.845000 74.865000 ;
        RECT  1.645000 75.070000  1.845000 75.270000 ;
        RECT  1.645000 75.475000  1.845000 75.675000 ;
        RECT  1.645000 75.880000  1.845000 76.080000 ;
        RECT  1.645000 76.285000  1.845000 76.485000 ;
        RECT  1.645000 76.690000  1.845000 76.890000 ;
        RECT  1.645000 77.095000  1.845000 77.295000 ;
        RECT  1.645000 77.500000  1.845000 77.700000 ;
        RECT  1.645000 77.905000  1.845000 78.105000 ;
        RECT  1.645000 78.310000  1.845000 78.510000 ;
        RECT  1.645000 78.715000  1.845000 78.915000 ;
        RECT  1.645000 79.120000  1.845000 79.320000 ;
        RECT  1.645000 79.525000  1.845000 79.725000 ;
        RECT  1.645000 79.930000  1.845000 80.130000 ;
        RECT  1.645000 80.335000  1.845000 80.535000 ;
        RECT  1.645000 80.740000  1.845000 80.940000 ;
        RECT  1.645000 81.145000  1.845000 81.345000 ;
        RECT  1.645000 81.550000  1.845000 81.750000 ;
        RECT  1.645000 81.955000  1.845000 82.155000 ;
        RECT  1.645000 82.360000  1.845000 82.560000 ;
        RECT  1.905000 17.860000  2.105000 18.060000 ;
        RECT  1.905000 18.290000  2.105000 18.490000 ;
        RECT  1.905000 18.720000  2.105000 18.920000 ;
        RECT  1.905000 19.150000  2.105000 19.350000 ;
        RECT  1.905000 19.580000  2.105000 19.780000 ;
        RECT  1.905000 20.010000  2.105000 20.210000 ;
        RECT  1.905000 20.440000  2.105000 20.640000 ;
        RECT  1.905000 20.870000  2.105000 21.070000 ;
        RECT  1.905000 21.300000  2.105000 21.500000 ;
        RECT  1.905000 21.730000  2.105000 21.930000 ;
        RECT  1.905000 22.160000  2.105000 22.360000 ;
        RECT  1.965000 82.855000  2.165000 83.055000 ;
        RECT  1.965000 83.265000  2.165000 83.465000 ;
        RECT  1.965000 83.675000  2.165000 83.875000 ;
        RECT  1.965000 84.085000  2.165000 84.285000 ;
        RECT  1.965000 84.495000  2.165000 84.695000 ;
        RECT  1.965000 84.905000  2.165000 85.105000 ;
        RECT  1.965000 85.315000  2.165000 85.515000 ;
        RECT  1.965000 85.725000  2.165000 85.925000 ;
        RECT  1.965000 86.135000  2.165000 86.335000 ;
        RECT  1.965000 86.545000  2.165000 86.745000 ;
        RECT  1.965000 86.955000  2.165000 87.155000 ;
        RECT  1.965000 87.365000  2.165000 87.565000 ;
        RECT  1.965000 87.775000  2.165000 87.975000 ;
        RECT  1.965000 88.185000  2.165000 88.385000 ;
        RECT  1.965000 88.595000  2.165000 88.795000 ;
        RECT  1.965000 89.005000  2.165000 89.205000 ;
        RECT  1.965000 89.415000  2.165000 89.615000 ;
        RECT  1.965000 89.825000  2.165000 90.025000 ;
        RECT  1.965000 90.235000  2.165000 90.435000 ;
        RECT  1.965000 90.645000  2.165000 90.845000 ;
        RECT  1.965000 91.055000  2.165000 91.255000 ;
        RECT  1.965000 91.465000  2.165000 91.665000 ;
        RECT  1.965000 91.875000  2.165000 92.075000 ;
        RECT  1.965000 92.285000  2.165000 92.485000 ;
        RECT  1.965000 92.695000  2.165000 92.895000 ;
        RECT  2.045000 68.125000  2.245000 68.325000 ;
        RECT  2.045000 68.535000  2.245000 68.735000 ;
        RECT  2.045000 68.945000  2.245000 69.145000 ;
        RECT  2.045000 69.355000  2.245000 69.555000 ;
        RECT  2.045000 69.765000  2.245000 69.965000 ;
        RECT  2.045000 70.175000  2.245000 70.375000 ;
        RECT  2.045000 70.585000  2.245000 70.785000 ;
        RECT  2.045000 70.995000  2.245000 71.195000 ;
        RECT  2.045000 71.405000  2.245000 71.605000 ;
        RECT  2.045000 71.815000  2.245000 72.015000 ;
        RECT  2.045000 72.225000  2.245000 72.425000 ;
        RECT  2.045000 72.635000  2.245000 72.835000 ;
        RECT  2.045000 73.045000  2.245000 73.245000 ;
        RECT  2.045000 73.450000  2.245000 73.650000 ;
        RECT  2.045000 73.855000  2.245000 74.055000 ;
        RECT  2.045000 74.260000  2.245000 74.460000 ;
        RECT  2.045000 74.665000  2.245000 74.865000 ;
        RECT  2.045000 75.070000  2.245000 75.270000 ;
        RECT  2.045000 75.475000  2.245000 75.675000 ;
        RECT  2.045000 75.880000  2.245000 76.080000 ;
        RECT  2.045000 76.285000  2.245000 76.485000 ;
        RECT  2.045000 76.690000  2.245000 76.890000 ;
        RECT  2.045000 77.095000  2.245000 77.295000 ;
        RECT  2.045000 77.500000  2.245000 77.700000 ;
        RECT  2.045000 77.905000  2.245000 78.105000 ;
        RECT  2.045000 78.310000  2.245000 78.510000 ;
        RECT  2.045000 78.715000  2.245000 78.915000 ;
        RECT  2.045000 79.120000  2.245000 79.320000 ;
        RECT  2.045000 79.525000  2.245000 79.725000 ;
        RECT  2.045000 79.930000  2.245000 80.130000 ;
        RECT  2.045000 80.335000  2.245000 80.535000 ;
        RECT  2.045000 80.740000  2.245000 80.940000 ;
        RECT  2.045000 81.145000  2.245000 81.345000 ;
        RECT  2.045000 81.550000  2.245000 81.750000 ;
        RECT  2.045000 81.955000  2.245000 82.155000 ;
        RECT  2.045000 82.360000  2.245000 82.560000 ;
        RECT  2.310000 17.860000  2.510000 18.060000 ;
        RECT  2.310000 18.290000  2.510000 18.490000 ;
        RECT  2.310000 18.720000  2.510000 18.920000 ;
        RECT  2.310000 19.150000  2.510000 19.350000 ;
        RECT  2.310000 19.580000  2.510000 19.780000 ;
        RECT  2.310000 20.010000  2.510000 20.210000 ;
        RECT  2.310000 20.440000  2.510000 20.640000 ;
        RECT  2.310000 20.870000  2.510000 21.070000 ;
        RECT  2.310000 21.300000  2.510000 21.500000 ;
        RECT  2.310000 21.730000  2.510000 21.930000 ;
        RECT  2.310000 22.160000  2.510000 22.360000 ;
        RECT  2.375000 82.855000  2.575000 83.055000 ;
        RECT  2.375000 83.265000  2.575000 83.465000 ;
        RECT  2.375000 83.675000  2.575000 83.875000 ;
        RECT  2.375000 84.085000  2.575000 84.285000 ;
        RECT  2.375000 84.495000  2.575000 84.695000 ;
        RECT  2.375000 84.905000  2.575000 85.105000 ;
        RECT  2.375000 85.315000  2.575000 85.515000 ;
        RECT  2.375000 85.725000  2.575000 85.925000 ;
        RECT  2.375000 86.135000  2.575000 86.335000 ;
        RECT  2.375000 86.545000  2.575000 86.745000 ;
        RECT  2.375000 86.955000  2.575000 87.155000 ;
        RECT  2.375000 87.365000  2.575000 87.565000 ;
        RECT  2.375000 87.775000  2.575000 87.975000 ;
        RECT  2.375000 88.185000  2.575000 88.385000 ;
        RECT  2.375000 88.595000  2.575000 88.795000 ;
        RECT  2.375000 89.005000  2.575000 89.205000 ;
        RECT  2.375000 89.415000  2.575000 89.615000 ;
        RECT  2.375000 89.825000  2.575000 90.025000 ;
        RECT  2.375000 90.235000  2.575000 90.435000 ;
        RECT  2.375000 90.645000  2.575000 90.845000 ;
        RECT  2.375000 91.055000  2.575000 91.255000 ;
        RECT  2.375000 91.465000  2.575000 91.665000 ;
        RECT  2.375000 91.875000  2.575000 92.075000 ;
        RECT  2.375000 92.285000  2.575000 92.485000 ;
        RECT  2.375000 92.695000  2.575000 92.895000 ;
        RECT  2.445000 68.125000  2.645000 68.325000 ;
        RECT  2.445000 68.535000  2.645000 68.735000 ;
        RECT  2.445000 68.945000  2.645000 69.145000 ;
        RECT  2.445000 69.355000  2.645000 69.555000 ;
        RECT  2.445000 69.765000  2.645000 69.965000 ;
        RECT  2.445000 70.175000  2.645000 70.375000 ;
        RECT  2.445000 70.585000  2.645000 70.785000 ;
        RECT  2.445000 70.995000  2.645000 71.195000 ;
        RECT  2.445000 71.405000  2.645000 71.605000 ;
        RECT  2.445000 71.815000  2.645000 72.015000 ;
        RECT  2.445000 72.225000  2.645000 72.425000 ;
        RECT  2.445000 72.635000  2.645000 72.835000 ;
        RECT  2.445000 73.045000  2.645000 73.245000 ;
        RECT  2.445000 73.450000  2.645000 73.650000 ;
        RECT  2.445000 73.855000  2.645000 74.055000 ;
        RECT  2.445000 74.260000  2.645000 74.460000 ;
        RECT  2.445000 74.665000  2.645000 74.865000 ;
        RECT  2.445000 75.070000  2.645000 75.270000 ;
        RECT  2.445000 75.475000  2.645000 75.675000 ;
        RECT  2.445000 75.880000  2.645000 76.080000 ;
        RECT  2.445000 76.285000  2.645000 76.485000 ;
        RECT  2.445000 76.690000  2.645000 76.890000 ;
        RECT  2.445000 77.095000  2.645000 77.295000 ;
        RECT  2.445000 77.500000  2.645000 77.700000 ;
        RECT  2.445000 77.905000  2.645000 78.105000 ;
        RECT  2.445000 78.310000  2.645000 78.510000 ;
        RECT  2.445000 78.715000  2.645000 78.915000 ;
        RECT  2.445000 79.120000  2.645000 79.320000 ;
        RECT  2.445000 79.525000  2.645000 79.725000 ;
        RECT  2.445000 79.930000  2.645000 80.130000 ;
        RECT  2.445000 80.335000  2.645000 80.535000 ;
        RECT  2.445000 80.740000  2.645000 80.940000 ;
        RECT  2.445000 81.145000  2.645000 81.345000 ;
        RECT  2.445000 81.550000  2.645000 81.750000 ;
        RECT  2.445000 81.955000  2.645000 82.155000 ;
        RECT  2.445000 82.360000  2.645000 82.560000 ;
        RECT  2.715000 17.860000  2.915000 18.060000 ;
        RECT  2.715000 18.290000  2.915000 18.490000 ;
        RECT  2.715000 18.720000  2.915000 18.920000 ;
        RECT  2.715000 19.150000  2.915000 19.350000 ;
        RECT  2.715000 19.580000  2.915000 19.780000 ;
        RECT  2.715000 20.010000  2.915000 20.210000 ;
        RECT  2.715000 20.440000  2.915000 20.640000 ;
        RECT  2.715000 20.870000  2.915000 21.070000 ;
        RECT  2.715000 21.300000  2.915000 21.500000 ;
        RECT  2.715000 21.730000  2.915000 21.930000 ;
        RECT  2.715000 22.160000  2.915000 22.360000 ;
        RECT  2.785000 82.855000  2.985000 83.055000 ;
        RECT  2.785000 83.265000  2.985000 83.465000 ;
        RECT  2.785000 83.675000  2.985000 83.875000 ;
        RECT  2.785000 84.085000  2.985000 84.285000 ;
        RECT  2.785000 84.495000  2.985000 84.695000 ;
        RECT  2.785000 84.905000  2.985000 85.105000 ;
        RECT  2.785000 85.315000  2.985000 85.515000 ;
        RECT  2.785000 85.725000  2.985000 85.925000 ;
        RECT  2.785000 86.135000  2.985000 86.335000 ;
        RECT  2.785000 86.545000  2.985000 86.745000 ;
        RECT  2.785000 86.955000  2.985000 87.155000 ;
        RECT  2.785000 87.365000  2.985000 87.565000 ;
        RECT  2.785000 87.775000  2.985000 87.975000 ;
        RECT  2.785000 88.185000  2.985000 88.385000 ;
        RECT  2.785000 88.595000  2.985000 88.795000 ;
        RECT  2.785000 89.005000  2.985000 89.205000 ;
        RECT  2.785000 89.415000  2.985000 89.615000 ;
        RECT  2.785000 89.825000  2.985000 90.025000 ;
        RECT  2.785000 90.235000  2.985000 90.435000 ;
        RECT  2.785000 90.645000  2.985000 90.845000 ;
        RECT  2.785000 91.055000  2.985000 91.255000 ;
        RECT  2.785000 91.465000  2.985000 91.665000 ;
        RECT  2.785000 91.875000  2.985000 92.075000 ;
        RECT  2.785000 92.285000  2.985000 92.485000 ;
        RECT  2.785000 92.695000  2.985000 92.895000 ;
        RECT  2.845000 68.125000  3.045000 68.325000 ;
        RECT  2.845000 68.535000  3.045000 68.735000 ;
        RECT  2.845000 68.945000  3.045000 69.145000 ;
        RECT  2.845000 69.355000  3.045000 69.555000 ;
        RECT  2.845000 69.765000  3.045000 69.965000 ;
        RECT  2.845000 70.175000  3.045000 70.375000 ;
        RECT  2.845000 70.585000  3.045000 70.785000 ;
        RECT  2.845000 70.995000  3.045000 71.195000 ;
        RECT  2.845000 71.405000  3.045000 71.605000 ;
        RECT  2.845000 71.815000  3.045000 72.015000 ;
        RECT  2.845000 72.225000  3.045000 72.425000 ;
        RECT  2.845000 72.635000  3.045000 72.835000 ;
        RECT  2.845000 73.045000  3.045000 73.245000 ;
        RECT  2.845000 73.450000  3.045000 73.650000 ;
        RECT  2.845000 73.855000  3.045000 74.055000 ;
        RECT  2.845000 74.260000  3.045000 74.460000 ;
        RECT  2.845000 74.665000  3.045000 74.865000 ;
        RECT  2.845000 75.070000  3.045000 75.270000 ;
        RECT  2.845000 75.475000  3.045000 75.675000 ;
        RECT  2.845000 75.880000  3.045000 76.080000 ;
        RECT  2.845000 76.285000  3.045000 76.485000 ;
        RECT  2.845000 76.690000  3.045000 76.890000 ;
        RECT  2.845000 77.095000  3.045000 77.295000 ;
        RECT  2.845000 77.500000  3.045000 77.700000 ;
        RECT  2.845000 77.905000  3.045000 78.105000 ;
        RECT  2.845000 78.310000  3.045000 78.510000 ;
        RECT  2.845000 78.715000  3.045000 78.915000 ;
        RECT  2.845000 79.120000  3.045000 79.320000 ;
        RECT  2.845000 79.525000  3.045000 79.725000 ;
        RECT  2.845000 79.930000  3.045000 80.130000 ;
        RECT  2.845000 80.335000  3.045000 80.535000 ;
        RECT  2.845000 80.740000  3.045000 80.940000 ;
        RECT  2.845000 81.145000  3.045000 81.345000 ;
        RECT  2.845000 81.550000  3.045000 81.750000 ;
        RECT  2.845000 81.955000  3.045000 82.155000 ;
        RECT  2.845000 82.360000  3.045000 82.560000 ;
        RECT  3.120000 17.860000  3.320000 18.060000 ;
        RECT  3.120000 18.290000  3.320000 18.490000 ;
        RECT  3.120000 18.720000  3.320000 18.920000 ;
        RECT  3.120000 19.150000  3.320000 19.350000 ;
        RECT  3.120000 19.580000  3.320000 19.780000 ;
        RECT  3.120000 20.010000  3.320000 20.210000 ;
        RECT  3.120000 20.440000  3.320000 20.640000 ;
        RECT  3.120000 20.870000  3.320000 21.070000 ;
        RECT  3.120000 21.300000  3.320000 21.500000 ;
        RECT  3.120000 21.730000  3.320000 21.930000 ;
        RECT  3.120000 22.160000  3.320000 22.360000 ;
        RECT  3.195000 82.855000  3.395000 83.055000 ;
        RECT  3.195000 83.265000  3.395000 83.465000 ;
        RECT  3.195000 83.675000  3.395000 83.875000 ;
        RECT  3.195000 84.085000  3.395000 84.285000 ;
        RECT  3.195000 84.495000  3.395000 84.695000 ;
        RECT  3.195000 84.905000  3.395000 85.105000 ;
        RECT  3.195000 85.315000  3.395000 85.515000 ;
        RECT  3.195000 85.725000  3.395000 85.925000 ;
        RECT  3.195000 86.135000  3.395000 86.335000 ;
        RECT  3.195000 86.545000  3.395000 86.745000 ;
        RECT  3.195000 86.955000  3.395000 87.155000 ;
        RECT  3.195000 87.365000  3.395000 87.565000 ;
        RECT  3.195000 87.775000  3.395000 87.975000 ;
        RECT  3.195000 88.185000  3.395000 88.385000 ;
        RECT  3.195000 88.595000  3.395000 88.795000 ;
        RECT  3.195000 89.005000  3.395000 89.205000 ;
        RECT  3.195000 89.415000  3.395000 89.615000 ;
        RECT  3.195000 89.825000  3.395000 90.025000 ;
        RECT  3.195000 90.235000  3.395000 90.435000 ;
        RECT  3.195000 90.645000  3.395000 90.845000 ;
        RECT  3.195000 91.055000  3.395000 91.255000 ;
        RECT  3.195000 91.465000  3.395000 91.665000 ;
        RECT  3.195000 91.875000  3.395000 92.075000 ;
        RECT  3.195000 92.285000  3.395000 92.485000 ;
        RECT  3.195000 92.695000  3.395000 92.895000 ;
        RECT  3.245000 68.125000  3.445000 68.325000 ;
        RECT  3.245000 68.535000  3.445000 68.735000 ;
        RECT  3.245000 68.945000  3.445000 69.145000 ;
        RECT  3.245000 69.355000  3.445000 69.555000 ;
        RECT  3.245000 69.765000  3.445000 69.965000 ;
        RECT  3.245000 70.175000  3.445000 70.375000 ;
        RECT  3.245000 70.585000  3.445000 70.785000 ;
        RECT  3.245000 70.995000  3.445000 71.195000 ;
        RECT  3.245000 71.405000  3.445000 71.605000 ;
        RECT  3.245000 71.815000  3.445000 72.015000 ;
        RECT  3.245000 72.225000  3.445000 72.425000 ;
        RECT  3.245000 72.635000  3.445000 72.835000 ;
        RECT  3.245000 73.045000  3.445000 73.245000 ;
        RECT  3.245000 73.450000  3.445000 73.650000 ;
        RECT  3.245000 73.855000  3.445000 74.055000 ;
        RECT  3.245000 74.260000  3.445000 74.460000 ;
        RECT  3.245000 74.665000  3.445000 74.865000 ;
        RECT  3.245000 75.070000  3.445000 75.270000 ;
        RECT  3.245000 75.475000  3.445000 75.675000 ;
        RECT  3.245000 75.880000  3.445000 76.080000 ;
        RECT  3.245000 76.285000  3.445000 76.485000 ;
        RECT  3.245000 76.690000  3.445000 76.890000 ;
        RECT  3.245000 77.095000  3.445000 77.295000 ;
        RECT  3.245000 77.500000  3.445000 77.700000 ;
        RECT  3.245000 77.905000  3.445000 78.105000 ;
        RECT  3.245000 78.310000  3.445000 78.510000 ;
        RECT  3.245000 78.715000  3.445000 78.915000 ;
        RECT  3.245000 79.120000  3.445000 79.320000 ;
        RECT  3.245000 79.525000  3.445000 79.725000 ;
        RECT  3.245000 79.930000  3.445000 80.130000 ;
        RECT  3.245000 80.335000  3.445000 80.535000 ;
        RECT  3.245000 80.740000  3.445000 80.940000 ;
        RECT  3.245000 81.145000  3.445000 81.345000 ;
        RECT  3.245000 81.550000  3.445000 81.750000 ;
        RECT  3.245000 81.955000  3.445000 82.155000 ;
        RECT  3.245000 82.360000  3.445000 82.560000 ;
        RECT  3.525000 17.860000  3.725000 18.060000 ;
        RECT  3.525000 18.290000  3.725000 18.490000 ;
        RECT  3.525000 18.720000  3.725000 18.920000 ;
        RECT  3.525000 19.150000  3.725000 19.350000 ;
        RECT  3.525000 19.580000  3.725000 19.780000 ;
        RECT  3.525000 20.010000  3.725000 20.210000 ;
        RECT  3.525000 20.440000  3.725000 20.640000 ;
        RECT  3.525000 20.870000  3.725000 21.070000 ;
        RECT  3.525000 21.300000  3.725000 21.500000 ;
        RECT  3.525000 21.730000  3.725000 21.930000 ;
        RECT  3.525000 22.160000  3.725000 22.360000 ;
        RECT  3.605000 82.855000  3.805000 83.055000 ;
        RECT  3.605000 83.265000  3.805000 83.465000 ;
        RECT  3.605000 83.675000  3.805000 83.875000 ;
        RECT  3.605000 84.085000  3.805000 84.285000 ;
        RECT  3.605000 84.495000  3.805000 84.695000 ;
        RECT  3.605000 84.905000  3.805000 85.105000 ;
        RECT  3.605000 85.315000  3.805000 85.515000 ;
        RECT  3.605000 85.725000  3.805000 85.925000 ;
        RECT  3.605000 86.135000  3.805000 86.335000 ;
        RECT  3.605000 86.545000  3.805000 86.745000 ;
        RECT  3.605000 86.955000  3.805000 87.155000 ;
        RECT  3.605000 87.365000  3.805000 87.565000 ;
        RECT  3.605000 87.775000  3.805000 87.975000 ;
        RECT  3.605000 88.185000  3.805000 88.385000 ;
        RECT  3.605000 88.595000  3.805000 88.795000 ;
        RECT  3.605000 89.005000  3.805000 89.205000 ;
        RECT  3.605000 89.415000  3.805000 89.615000 ;
        RECT  3.605000 89.825000  3.805000 90.025000 ;
        RECT  3.605000 90.235000  3.805000 90.435000 ;
        RECT  3.605000 90.645000  3.805000 90.845000 ;
        RECT  3.605000 91.055000  3.805000 91.255000 ;
        RECT  3.605000 91.465000  3.805000 91.665000 ;
        RECT  3.605000 91.875000  3.805000 92.075000 ;
        RECT  3.605000 92.285000  3.805000 92.485000 ;
        RECT  3.605000 92.695000  3.805000 92.895000 ;
        RECT  3.645000 68.125000  3.845000 68.325000 ;
        RECT  3.645000 68.535000  3.845000 68.735000 ;
        RECT  3.645000 68.945000  3.845000 69.145000 ;
        RECT  3.645000 69.355000  3.845000 69.555000 ;
        RECT  3.645000 69.765000  3.845000 69.965000 ;
        RECT  3.645000 70.175000  3.845000 70.375000 ;
        RECT  3.645000 70.585000  3.845000 70.785000 ;
        RECT  3.645000 70.995000  3.845000 71.195000 ;
        RECT  3.645000 71.405000  3.845000 71.605000 ;
        RECT  3.645000 71.815000  3.845000 72.015000 ;
        RECT  3.645000 72.225000  3.845000 72.425000 ;
        RECT  3.645000 72.635000  3.845000 72.835000 ;
        RECT  3.645000 73.045000  3.845000 73.245000 ;
        RECT  3.645000 73.450000  3.845000 73.650000 ;
        RECT  3.645000 73.855000  3.845000 74.055000 ;
        RECT  3.645000 74.260000  3.845000 74.460000 ;
        RECT  3.645000 74.665000  3.845000 74.865000 ;
        RECT  3.645000 75.070000  3.845000 75.270000 ;
        RECT  3.645000 75.475000  3.845000 75.675000 ;
        RECT  3.645000 75.880000  3.845000 76.080000 ;
        RECT  3.645000 76.285000  3.845000 76.485000 ;
        RECT  3.645000 76.690000  3.845000 76.890000 ;
        RECT  3.645000 77.095000  3.845000 77.295000 ;
        RECT  3.645000 77.500000  3.845000 77.700000 ;
        RECT  3.645000 77.905000  3.845000 78.105000 ;
        RECT  3.645000 78.310000  3.845000 78.510000 ;
        RECT  3.645000 78.715000  3.845000 78.915000 ;
        RECT  3.645000 79.120000  3.845000 79.320000 ;
        RECT  3.645000 79.525000  3.845000 79.725000 ;
        RECT  3.645000 79.930000  3.845000 80.130000 ;
        RECT  3.645000 80.335000  3.845000 80.535000 ;
        RECT  3.645000 80.740000  3.845000 80.940000 ;
        RECT  3.645000 81.145000  3.845000 81.345000 ;
        RECT  3.645000 81.550000  3.845000 81.750000 ;
        RECT  3.645000 81.955000  3.845000 82.155000 ;
        RECT  3.645000 82.360000  3.845000 82.560000 ;
        RECT  3.930000 17.860000  4.130000 18.060000 ;
        RECT  3.930000 18.290000  4.130000 18.490000 ;
        RECT  3.930000 18.720000  4.130000 18.920000 ;
        RECT  3.930000 19.150000  4.130000 19.350000 ;
        RECT  3.930000 19.580000  4.130000 19.780000 ;
        RECT  3.930000 20.010000  4.130000 20.210000 ;
        RECT  3.930000 20.440000  4.130000 20.640000 ;
        RECT  3.930000 20.870000  4.130000 21.070000 ;
        RECT  3.930000 21.300000  4.130000 21.500000 ;
        RECT  3.930000 21.730000  4.130000 21.930000 ;
        RECT  3.930000 22.160000  4.130000 22.360000 ;
        RECT  4.015000 82.855000  4.215000 83.055000 ;
        RECT  4.015000 83.265000  4.215000 83.465000 ;
        RECT  4.015000 83.675000  4.215000 83.875000 ;
        RECT  4.015000 84.085000  4.215000 84.285000 ;
        RECT  4.015000 84.495000  4.215000 84.695000 ;
        RECT  4.015000 84.905000  4.215000 85.105000 ;
        RECT  4.015000 85.315000  4.215000 85.515000 ;
        RECT  4.015000 85.725000  4.215000 85.925000 ;
        RECT  4.015000 86.135000  4.215000 86.335000 ;
        RECT  4.015000 86.545000  4.215000 86.745000 ;
        RECT  4.015000 86.955000  4.215000 87.155000 ;
        RECT  4.015000 87.365000  4.215000 87.565000 ;
        RECT  4.015000 87.775000  4.215000 87.975000 ;
        RECT  4.015000 88.185000  4.215000 88.385000 ;
        RECT  4.015000 88.595000  4.215000 88.795000 ;
        RECT  4.015000 89.005000  4.215000 89.205000 ;
        RECT  4.015000 89.415000  4.215000 89.615000 ;
        RECT  4.015000 89.825000  4.215000 90.025000 ;
        RECT  4.015000 90.235000  4.215000 90.435000 ;
        RECT  4.015000 90.645000  4.215000 90.845000 ;
        RECT  4.015000 91.055000  4.215000 91.255000 ;
        RECT  4.015000 91.465000  4.215000 91.665000 ;
        RECT  4.015000 91.875000  4.215000 92.075000 ;
        RECT  4.015000 92.285000  4.215000 92.485000 ;
        RECT  4.015000 92.695000  4.215000 92.895000 ;
        RECT  4.045000 68.125000  4.245000 68.325000 ;
        RECT  4.045000 68.535000  4.245000 68.735000 ;
        RECT  4.045000 68.945000  4.245000 69.145000 ;
        RECT  4.045000 69.355000  4.245000 69.555000 ;
        RECT  4.045000 69.765000  4.245000 69.965000 ;
        RECT  4.045000 70.175000  4.245000 70.375000 ;
        RECT  4.045000 70.585000  4.245000 70.785000 ;
        RECT  4.045000 70.995000  4.245000 71.195000 ;
        RECT  4.045000 71.405000  4.245000 71.605000 ;
        RECT  4.045000 71.815000  4.245000 72.015000 ;
        RECT  4.045000 72.225000  4.245000 72.425000 ;
        RECT  4.045000 72.635000  4.245000 72.835000 ;
        RECT  4.045000 73.045000  4.245000 73.245000 ;
        RECT  4.045000 73.450000  4.245000 73.650000 ;
        RECT  4.045000 73.855000  4.245000 74.055000 ;
        RECT  4.045000 74.260000  4.245000 74.460000 ;
        RECT  4.045000 74.665000  4.245000 74.865000 ;
        RECT  4.045000 75.070000  4.245000 75.270000 ;
        RECT  4.045000 75.475000  4.245000 75.675000 ;
        RECT  4.045000 75.880000  4.245000 76.080000 ;
        RECT  4.045000 76.285000  4.245000 76.485000 ;
        RECT  4.045000 76.690000  4.245000 76.890000 ;
        RECT  4.045000 77.095000  4.245000 77.295000 ;
        RECT  4.045000 77.500000  4.245000 77.700000 ;
        RECT  4.045000 77.905000  4.245000 78.105000 ;
        RECT  4.045000 78.310000  4.245000 78.510000 ;
        RECT  4.045000 78.715000  4.245000 78.915000 ;
        RECT  4.045000 79.120000  4.245000 79.320000 ;
        RECT  4.045000 79.525000  4.245000 79.725000 ;
        RECT  4.045000 79.930000  4.245000 80.130000 ;
        RECT  4.045000 80.335000  4.245000 80.535000 ;
        RECT  4.045000 80.740000  4.245000 80.940000 ;
        RECT  4.045000 81.145000  4.245000 81.345000 ;
        RECT  4.045000 81.550000  4.245000 81.750000 ;
        RECT  4.045000 81.955000  4.245000 82.155000 ;
        RECT  4.045000 82.360000  4.245000 82.560000 ;
        RECT  4.335000 17.860000  4.535000 18.060000 ;
        RECT  4.335000 18.290000  4.535000 18.490000 ;
        RECT  4.335000 18.720000  4.535000 18.920000 ;
        RECT  4.335000 19.150000  4.535000 19.350000 ;
        RECT  4.335000 19.580000  4.535000 19.780000 ;
        RECT  4.335000 20.010000  4.535000 20.210000 ;
        RECT  4.335000 20.440000  4.535000 20.640000 ;
        RECT  4.335000 20.870000  4.535000 21.070000 ;
        RECT  4.335000 21.300000  4.535000 21.500000 ;
        RECT  4.335000 21.730000  4.535000 21.930000 ;
        RECT  4.335000 22.160000  4.535000 22.360000 ;
        RECT  4.425000 82.855000  4.625000 83.055000 ;
        RECT  4.425000 83.265000  4.625000 83.465000 ;
        RECT  4.425000 83.675000  4.625000 83.875000 ;
        RECT  4.425000 84.085000  4.625000 84.285000 ;
        RECT  4.425000 84.495000  4.625000 84.695000 ;
        RECT  4.425000 84.905000  4.625000 85.105000 ;
        RECT  4.425000 85.315000  4.625000 85.515000 ;
        RECT  4.425000 85.725000  4.625000 85.925000 ;
        RECT  4.425000 86.135000  4.625000 86.335000 ;
        RECT  4.425000 86.545000  4.625000 86.745000 ;
        RECT  4.425000 86.955000  4.625000 87.155000 ;
        RECT  4.425000 87.365000  4.625000 87.565000 ;
        RECT  4.425000 87.775000  4.625000 87.975000 ;
        RECT  4.425000 88.185000  4.625000 88.385000 ;
        RECT  4.425000 88.595000  4.625000 88.795000 ;
        RECT  4.425000 89.005000  4.625000 89.205000 ;
        RECT  4.425000 89.415000  4.625000 89.615000 ;
        RECT  4.425000 89.825000  4.625000 90.025000 ;
        RECT  4.425000 90.235000  4.625000 90.435000 ;
        RECT  4.425000 90.645000  4.625000 90.845000 ;
        RECT  4.425000 91.055000  4.625000 91.255000 ;
        RECT  4.425000 91.465000  4.625000 91.665000 ;
        RECT  4.425000 91.875000  4.625000 92.075000 ;
        RECT  4.425000 92.285000  4.625000 92.485000 ;
        RECT  4.425000 92.695000  4.625000 92.895000 ;
        RECT  4.445000 68.125000  4.645000 68.325000 ;
        RECT  4.445000 68.535000  4.645000 68.735000 ;
        RECT  4.445000 68.945000  4.645000 69.145000 ;
        RECT  4.445000 69.355000  4.645000 69.555000 ;
        RECT  4.445000 69.765000  4.645000 69.965000 ;
        RECT  4.445000 70.175000  4.645000 70.375000 ;
        RECT  4.445000 70.585000  4.645000 70.785000 ;
        RECT  4.445000 70.995000  4.645000 71.195000 ;
        RECT  4.445000 71.405000  4.645000 71.605000 ;
        RECT  4.445000 71.815000  4.645000 72.015000 ;
        RECT  4.445000 72.225000  4.645000 72.425000 ;
        RECT  4.445000 72.635000  4.645000 72.835000 ;
        RECT  4.445000 73.045000  4.645000 73.245000 ;
        RECT  4.445000 73.450000  4.645000 73.650000 ;
        RECT  4.445000 73.855000  4.645000 74.055000 ;
        RECT  4.445000 74.260000  4.645000 74.460000 ;
        RECT  4.445000 74.665000  4.645000 74.865000 ;
        RECT  4.445000 75.070000  4.645000 75.270000 ;
        RECT  4.445000 75.475000  4.645000 75.675000 ;
        RECT  4.445000 75.880000  4.645000 76.080000 ;
        RECT  4.445000 76.285000  4.645000 76.485000 ;
        RECT  4.445000 76.690000  4.645000 76.890000 ;
        RECT  4.445000 77.095000  4.645000 77.295000 ;
        RECT  4.445000 77.500000  4.645000 77.700000 ;
        RECT  4.445000 77.905000  4.645000 78.105000 ;
        RECT  4.445000 78.310000  4.645000 78.510000 ;
        RECT  4.445000 78.715000  4.645000 78.915000 ;
        RECT  4.445000 79.120000  4.645000 79.320000 ;
        RECT  4.445000 79.525000  4.645000 79.725000 ;
        RECT  4.445000 79.930000  4.645000 80.130000 ;
        RECT  4.445000 80.335000  4.645000 80.535000 ;
        RECT  4.445000 80.740000  4.645000 80.940000 ;
        RECT  4.445000 81.145000  4.645000 81.345000 ;
        RECT  4.445000 81.550000  4.645000 81.750000 ;
        RECT  4.445000 81.955000  4.645000 82.155000 ;
        RECT  4.445000 82.360000  4.645000 82.560000 ;
        RECT  4.740000 17.860000  4.940000 18.060000 ;
        RECT  4.740000 18.290000  4.940000 18.490000 ;
        RECT  4.740000 18.720000  4.940000 18.920000 ;
        RECT  4.740000 19.150000  4.940000 19.350000 ;
        RECT  4.740000 19.580000  4.940000 19.780000 ;
        RECT  4.740000 20.010000  4.940000 20.210000 ;
        RECT  4.740000 20.440000  4.940000 20.640000 ;
        RECT  4.740000 20.870000  4.940000 21.070000 ;
        RECT  4.740000 21.300000  4.940000 21.500000 ;
        RECT  4.740000 21.730000  4.940000 21.930000 ;
        RECT  4.740000 22.160000  4.940000 22.360000 ;
        RECT  4.835000 82.855000  5.035000 83.055000 ;
        RECT  4.835000 83.265000  5.035000 83.465000 ;
        RECT  4.835000 83.675000  5.035000 83.875000 ;
        RECT  4.835000 84.085000  5.035000 84.285000 ;
        RECT  4.835000 84.495000  5.035000 84.695000 ;
        RECT  4.835000 84.905000  5.035000 85.105000 ;
        RECT  4.835000 85.315000  5.035000 85.515000 ;
        RECT  4.835000 85.725000  5.035000 85.925000 ;
        RECT  4.835000 86.135000  5.035000 86.335000 ;
        RECT  4.835000 86.545000  5.035000 86.745000 ;
        RECT  4.835000 86.955000  5.035000 87.155000 ;
        RECT  4.835000 87.365000  5.035000 87.565000 ;
        RECT  4.835000 87.775000  5.035000 87.975000 ;
        RECT  4.835000 88.185000  5.035000 88.385000 ;
        RECT  4.835000 88.595000  5.035000 88.795000 ;
        RECT  4.835000 89.005000  5.035000 89.205000 ;
        RECT  4.835000 89.415000  5.035000 89.615000 ;
        RECT  4.835000 89.825000  5.035000 90.025000 ;
        RECT  4.835000 90.235000  5.035000 90.435000 ;
        RECT  4.835000 90.645000  5.035000 90.845000 ;
        RECT  4.835000 91.055000  5.035000 91.255000 ;
        RECT  4.835000 91.465000  5.035000 91.665000 ;
        RECT  4.835000 91.875000  5.035000 92.075000 ;
        RECT  4.835000 92.285000  5.035000 92.485000 ;
        RECT  4.835000 92.695000  5.035000 92.895000 ;
        RECT  4.845000 68.125000  5.045000 68.325000 ;
        RECT  4.845000 68.535000  5.045000 68.735000 ;
        RECT  4.845000 68.945000  5.045000 69.145000 ;
        RECT  4.845000 69.355000  5.045000 69.555000 ;
        RECT  4.845000 69.765000  5.045000 69.965000 ;
        RECT  4.845000 70.175000  5.045000 70.375000 ;
        RECT  4.845000 70.585000  5.045000 70.785000 ;
        RECT  4.845000 70.995000  5.045000 71.195000 ;
        RECT  4.845000 71.405000  5.045000 71.605000 ;
        RECT  4.845000 71.815000  5.045000 72.015000 ;
        RECT  4.845000 72.225000  5.045000 72.425000 ;
        RECT  4.845000 72.635000  5.045000 72.835000 ;
        RECT  4.845000 73.045000  5.045000 73.245000 ;
        RECT  4.845000 73.450000  5.045000 73.650000 ;
        RECT  4.845000 73.855000  5.045000 74.055000 ;
        RECT  4.845000 74.260000  5.045000 74.460000 ;
        RECT  4.845000 74.665000  5.045000 74.865000 ;
        RECT  4.845000 75.070000  5.045000 75.270000 ;
        RECT  4.845000 75.475000  5.045000 75.675000 ;
        RECT  4.845000 75.880000  5.045000 76.080000 ;
        RECT  4.845000 76.285000  5.045000 76.485000 ;
        RECT  4.845000 76.690000  5.045000 76.890000 ;
        RECT  4.845000 77.095000  5.045000 77.295000 ;
        RECT  4.845000 77.500000  5.045000 77.700000 ;
        RECT  4.845000 77.905000  5.045000 78.105000 ;
        RECT  4.845000 78.310000  5.045000 78.510000 ;
        RECT  4.845000 78.715000  5.045000 78.915000 ;
        RECT  4.845000 79.120000  5.045000 79.320000 ;
        RECT  4.845000 79.525000  5.045000 79.725000 ;
        RECT  4.845000 79.930000  5.045000 80.130000 ;
        RECT  4.845000 80.335000  5.045000 80.535000 ;
        RECT  4.845000 80.740000  5.045000 80.940000 ;
        RECT  4.845000 81.145000  5.045000 81.345000 ;
        RECT  4.845000 81.550000  5.045000 81.750000 ;
        RECT  4.845000 81.955000  5.045000 82.155000 ;
        RECT  4.845000 82.360000  5.045000 82.560000 ;
        RECT  5.145000 17.860000  5.345000 18.060000 ;
        RECT  5.145000 18.290000  5.345000 18.490000 ;
        RECT  5.145000 18.720000  5.345000 18.920000 ;
        RECT  5.145000 19.150000  5.345000 19.350000 ;
        RECT  5.145000 19.580000  5.345000 19.780000 ;
        RECT  5.145000 20.010000  5.345000 20.210000 ;
        RECT  5.145000 20.440000  5.345000 20.640000 ;
        RECT  5.145000 20.870000  5.345000 21.070000 ;
        RECT  5.145000 21.300000  5.345000 21.500000 ;
        RECT  5.145000 21.730000  5.345000 21.930000 ;
        RECT  5.145000 22.160000  5.345000 22.360000 ;
        RECT  5.245000 68.125000  5.445000 68.325000 ;
        RECT  5.245000 68.535000  5.445000 68.735000 ;
        RECT  5.245000 68.945000  5.445000 69.145000 ;
        RECT  5.245000 69.355000  5.445000 69.555000 ;
        RECT  5.245000 69.765000  5.445000 69.965000 ;
        RECT  5.245000 70.175000  5.445000 70.375000 ;
        RECT  5.245000 70.585000  5.445000 70.785000 ;
        RECT  5.245000 70.995000  5.445000 71.195000 ;
        RECT  5.245000 71.405000  5.445000 71.605000 ;
        RECT  5.245000 71.815000  5.445000 72.015000 ;
        RECT  5.245000 72.225000  5.445000 72.425000 ;
        RECT  5.245000 72.635000  5.445000 72.835000 ;
        RECT  5.245000 73.045000  5.445000 73.245000 ;
        RECT  5.245000 73.450000  5.445000 73.650000 ;
        RECT  5.245000 73.855000  5.445000 74.055000 ;
        RECT  5.245000 74.260000  5.445000 74.460000 ;
        RECT  5.245000 74.665000  5.445000 74.865000 ;
        RECT  5.245000 75.070000  5.445000 75.270000 ;
        RECT  5.245000 75.475000  5.445000 75.675000 ;
        RECT  5.245000 75.880000  5.445000 76.080000 ;
        RECT  5.245000 76.285000  5.445000 76.485000 ;
        RECT  5.245000 76.690000  5.445000 76.890000 ;
        RECT  5.245000 77.095000  5.445000 77.295000 ;
        RECT  5.245000 77.500000  5.445000 77.700000 ;
        RECT  5.245000 77.905000  5.445000 78.105000 ;
        RECT  5.245000 78.310000  5.445000 78.510000 ;
        RECT  5.245000 78.715000  5.445000 78.915000 ;
        RECT  5.245000 79.120000  5.445000 79.320000 ;
        RECT  5.245000 79.525000  5.445000 79.725000 ;
        RECT  5.245000 79.930000  5.445000 80.130000 ;
        RECT  5.245000 80.335000  5.445000 80.535000 ;
        RECT  5.245000 80.740000  5.445000 80.940000 ;
        RECT  5.245000 81.145000  5.445000 81.345000 ;
        RECT  5.245000 81.550000  5.445000 81.750000 ;
        RECT  5.245000 81.955000  5.445000 82.155000 ;
        RECT  5.245000 82.360000  5.445000 82.560000 ;
        RECT  5.245000 82.855000  5.445000 83.055000 ;
        RECT  5.245000 83.265000  5.445000 83.465000 ;
        RECT  5.245000 83.675000  5.445000 83.875000 ;
        RECT  5.245000 84.085000  5.445000 84.285000 ;
        RECT  5.245000 84.495000  5.445000 84.695000 ;
        RECT  5.245000 84.905000  5.445000 85.105000 ;
        RECT  5.245000 85.315000  5.445000 85.515000 ;
        RECT  5.245000 85.725000  5.445000 85.925000 ;
        RECT  5.245000 86.135000  5.445000 86.335000 ;
        RECT  5.245000 86.545000  5.445000 86.745000 ;
        RECT  5.245000 86.955000  5.445000 87.155000 ;
        RECT  5.245000 87.365000  5.445000 87.565000 ;
        RECT  5.245000 87.775000  5.445000 87.975000 ;
        RECT  5.245000 88.185000  5.445000 88.385000 ;
        RECT  5.245000 88.595000  5.445000 88.795000 ;
        RECT  5.245000 89.005000  5.445000 89.205000 ;
        RECT  5.245000 89.415000  5.445000 89.615000 ;
        RECT  5.245000 89.825000  5.445000 90.025000 ;
        RECT  5.245000 90.235000  5.445000 90.435000 ;
        RECT  5.245000 90.645000  5.445000 90.845000 ;
        RECT  5.245000 91.055000  5.445000 91.255000 ;
        RECT  5.245000 91.465000  5.445000 91.665000 ;
        RECT  5.245000 91.875000  5.445000 92.075000 ;
        RECT  5.245000 92.285000  5.445000 92.485000 ;
        RECT  5.245000 92.695000  5.445000 92.895000 ;
        RECT  5.550000 17.860000  5.750000 18.060000 ;
        RECT  5.550000 18.290000  5.750000 18.490000 ;
        RECT  5.550000 18.720000  5.750000 18.920000 ;
        RECT  5.550000 19.150000  5.750000 19.350000 ;
        RECT  5.550000 19.580000  5.750000 19.780000 ;
        RECT  5.550000 20.010000  5.750000 20.210000 ;
        RECT  5.550000 20.440000  5.750000 20.640000 ;
        RECT  5.550000 20.870000  5.750000 21.070000 ;
        RECT  5.550000 21.300000  5.750000 21.500000 ;
        RECT  5.550000 21.730000  5.750000 21.930000 ;
        RECT  5.550000 22.160000  5.750000 22.360000 ;
        RECT  5.645000 68.125000  5.845000 68.325000 ;
        RECT  5.645000 68.535000  5.845000 68.735000 ;
        RECT  5.645000 68.945000  5.845000 69.145000 ;
        RECT  5.645000 69.355000  5.845000 69.555000 ;
        RECT  5.645000 69.765000  5.845000 69.965000 ;
        RECT  5.645000 70.175000  5.845000 70.375000 ;
        RECT  5.645000 70.585000  5.845000 70.785000 ;
        RECT  5.645000 70.995000  5.845000 71.195000 ;
        RECT  5.645000 71.405000  5.845000 71.605000 ;
        RECT  5.645000 71.815000  5.845000 72.015000 ;
        RECT  5.645000 72.225000  5.845000 72.425000 ;
        RECT  5.645000 72.635000  5.845000 72.835000 ;
        RECT  5.645000 73.045000  5.845000 73.245000 ;
        RECT  5.645000 73.450000  5.845000 73.650000 ;
        RECT  5.645000 73.855000  5.845000 74.055000 ;
        RECT  5.645000 74.260000  5.845000 74.460000 ;
        RECT  5.645000 74.665000  5.845000 74.865000 ;
        RECT  5.645000 75.070000  5.845000 75.270000 ;
        RECT  5.645000 75.475000  5.845000 75.675000 ;
        RECT  5.645000 75.880000  5.845000 76.080000 ;
        RECT  5.645000 76.285000  5.845000 76.485000 ;
        RECT  5.645000 76.690000  5.845000 76.890000 ;
        RECT  5.645000 77.095000  5.845000 77.295000 ;
        RECT  5.645000 77.500000  5.845000 77.700000 ;
        RECT  5.645000 77.905000  5.845000 78.105000 ;
        RECT  5.645000 78.310000  5.845000 78.510000 ;
        RECT  5.645000 78.715000  5.845000 78.915000 ;
        RECT  5.645000 79.120000  5.845000 79.320000 ;
        RECT  5.645000 79.525000  5.845000 79.725000 ;
        RECT  5.645000 79.930000  5.845000 80.130000 ;
        RECT  5.645000 80.335000  5.845000 80.535000 ;
        RECT  5.645000 80.740000  5.845000 80.940000 ;
        RECT  5.645000 81.145000  5.845000 81.345000 ;
        RECT  5.645000 81.550000  5.845000 81.750000 ;
        RECT  5.645000 81.955000  5.845000 82.155000 ;
        RECT  5.645000 82.360000  5.845000 82.560000 ;
        RECT  5.655000 82.855000  5.855000 83.055000 ;
        RECT  5.655000 83.265000  5.855000 83.465000 ;
        RECT  5.655000 83.675000  5.855000 83.875000 ;
        RECT  5.655000 84.085000  5.855000 84.285000 ;
        RECT  5.655000 84.495000  5.855000 84.695000 ;
        RECT  5.655000 84.905000  5.855000 85.105000 ;
        RECT  5.655000 85.315000  5.855000 85.515000 ;
        RECT  5.655000 85.725000  5.855000 85.925000 ;
        RECT  5.655000 86.135000  5.855000 86.335000 ;
        RECT  5.655000 86.545000  5.855000 86.745000 ;
        RECT  5.655000 86.955000  5.855000 87.155000 ;
        RECT  5.655000 87.365000  5.855000 87.565000 ;
        RECT  5.655000 87.775000  5.855000 87.975000 ;
        RECT  5.655000 88.185000  5.855000 88.385000 ;
        RECT  5.655000 88.595000  5.855000 88.795000 ;
        RECT  5.655000 89.005000  5.855000 89.205000 ;
        RECT  5.655000 89.415000  5.855000 89.615000 ;
        RECT  5.655000 89.825000  5.855000 90.025000 ;
        RECT  5.655000 90.235000  5.855000 90.435000 ;
        RECT  5.655000 90.645000  5.855000 90.845000 ;
        RECT  5.655000 91.055000  5.855000 91.255000 ;
        RECT  5.655000 91.465000  5.855000 91.665000 ;
        RECT  5.655000 91.875000  5.855000 92.075000 ;
        RECT  5.655000 92.285000  5.855000 92.485000 ;
        RECT  5.655000 92.695000  5.855000 92.895000 ;
        RECT  5.955000 17.860000  6.155000 18.060000 ;
        RECT  5.955000 18.290000  6.155000 18.490000 ;
        RECT  5.955000 18.720000  6.155000 18.920000 ;
        RECT  5.955000 19.150000  6.155000 19.350000 ;
        RECT  5.955000 19.580000  6.155000 19.780000 ;
        RECT  5.955000 20.010000  6.155000 20.210000 ;
        RECT  5.955000 20.440000  6.155000 20.640000 ;
        RECT  5.955000 20.870000  6.155000 21.070000 ;
        RECT  5.955000 21.300000  6.155000 21.500000 ;
        RECT  5.955000 21.730000  6.155000 21.930000 ;
        RECT  5.955000 22.160000  6.155000 22.360000 ;
        RECT  6.045000 68.125000  6.245000 68.325000 ;
        RECT  6.045000 68.535000  6.245000 68.735000 ;
        RECT  6.045000 68.945000  6.245000 69.145000 ;
        RECT  6.045000 69.355000  6.245000 69.555000 ;
        RECT  6.045000 69.765000  6.245000 69.965000 ;
        RECT  6.045000 70.175000  6.245000 70.375000 ;
        RECT  6.045000 70.585000  6.245000 70.785000 ;
        RECT  6.045000 70.995000  6.245000 71.195000 ;
        RECT  6.045000 71.405000  6.245000 71.605000 ;
        RECT  6.045000 71.815000  6.245000 72.015000 ;
        RECT  6.045000 72.225000  6.245000 72.425000 ;
        RECT  6.045000 72.635000  6.245000 72.835000 ;
        RECT  6.045000 73.045000  6.245000 73.245000 ;
        RECT  6.045000 73.450000  6.245000 73.650000 ;
        RECT  6.045000 73.855000  6.245000 74.055000 ;
        RECT  6.045000 74.260000  6.245000 74.460000 ;
        RECT  6.045000 74.665000  6.245000 74.865000 ;
        RECT  6.045000 75.070000  6.245000 75.270000 ;
        RECT  6.045000 75.475000  6.245000 75.675000 ;
        RECT  6.045000 75.880000  6.245000 76.080000 ;
        RECT  6.045000 76.285000  6.245000 76.485000 ;
        RECT  6.045000 76.690000  6.245000 76.890000 ;
        RECT  6.045000 77.095000  6.245000 77.295000 ;
        RECT  6.045000 77.500000  6.245000 77.700000 ;
        RECT  6.045000 77.905000  6.245000 78.105000 ;
        RECT  6.045000 78.310000  6.245000 78.510000 ;
        RECT  6.045000 78.715000  6.245000 78.915000 ;
        RECT  6.045000 79.120000  6.245000 79.320000 ;
        RECT  6.045000 79.525000  6.245000 79.725000 ;
        RECT  6.045000 79.930000  6.245000 80.130000 ;
        RECT  6.045000 80.335000  6.245000 80.535000 ;
        RECT  6.045000 80.740000  6.245000 80.940000 ;
        RECT  6.045000 81.145000  6.245000 81.345000 ;
        RECT  6.045000 81.550000  6.245000 81.750000 ;
        RECT  6.045000 81.955000  6.245000 82.155000 ;
        RECT  6.045000 82.360000  6.245000 82.560000 ;
        RECT  6.065000 82.855000  6.265000 83.055000 ;
        RECT  6.065000 83.265000  6.265000 83.465000 ;
        RECT  6.065000 83.675000  6.265000 83.875000 ;
        RECT  6.065000 84.085000  6.265000 84.285000 ;
        RECT  6.065000 84.495000  6.265000 84.695000 ;
        RECT  6.065000 84.905000  6.265000 85.105000 ;
        RECT  6.065000 85.315000  6.265000 85.515000 ;
        RECT  6.065000 85.725000  6.265000 85.925000 ;
        RECT  6.065000 86.135000  6.265000 86.335000 ;
        RECT  6.065000 86.545000  6.265000 86.745000 ;
        RECT  6.065000 86.955000  6.265000 87.155000 ;
        RECT  6.065000 87.365000  6.265000 87.565000 ;
        RECT  6.065000 87.775000  6.265000 87.975000 ;
        RECT  6.065000 88.185000  6.265000 88.385000 ;
        RECT  6.065000 88.595000  6.265000 88.795000 ;
        RECT  6.065000 89.005000  6.265000 89.205000 ;
        RECT  6.065000 89.415000  6.265000 89.615000 ;
        RECT  6.065000 89.825000  6.265000 90.025000 ;
        RECT  6.065000 90.235000  6.265000 90.435000 ;
        RECT  6.065000 90.645000  6.265000 90.845000 ;
        RECT  6.065000 91.055000  6.265000 91.255000 ;
        RECT  6.065000 91.465000  6.265000 91.665000 ;
        RECT  6.065000 91.875000  6.265000 92.075000 ;
        RECT  6.065000 92.285000  6.265000 92.485000 ;
        RECT  6.065000 92.695000  6.265000 92.895000 ;
        RECT  6.360000 17.860000  6.560000 18.060000 ;
        RECT  6.360000 18.290000  6.560000 18.490000 ;
        RECT  6.360000 18.720000  6.560000 18.920000 ;
        RECT  6.360000 19.150000  6.560000 19.350000 ;
        RECT  6.360000 19.580000  6.560000 19.780000 ;
        RECT  6.360000 20.010000  6.560000 20.210000 ;
        RECT  6.360000 20.440000  6.560000 20.640000 ;
        RECT  6.360000 20.870000  6.560000 21.070000 ;
        RECT  6.360000 21.300000  6.560000 21.500000 ;
        RECT  6.360000 21.730000  6.560000 21.930000 ;
        RECT  6.360000 22.160000  6.560000 22.360000 ;
        RECT  6.445000 68.125000  6.645000 68.325000 ;
        RECT  6.445000 68.535000  6.645000 68.735000 ;
        RECT  6.445000 68.945000  6.645000 69.145000 ;
        RECT  6.445000 69.355000  6.645000 69.555000 ;
        RECT  6.445000 69.765000  6.645000 69.965000 ;
        RECT  6.445000 70.175000  6.645000 70.375000 ;
        RECT  6.445000 70.585000  6.645000 70.785000 ;
        RECT  6.445000 70.995000  6.645000 71.195000 ;
        RECT  6.445000 71.405000  6.645000 71.605000 ;
        RECT  6.445000 71.815000  6.645000 72.015000 ;
        RECT  6.445000 72.225000  6.645000 72.425000 ;
        RECT  6.445000 72.635000  6.645000 72.835000 ;
        RECT  6.445000 73.045000  6.645000 73.245000 ;
        RECT  6.445000 73.450000  6.645000 73.650000 ;
        RECT  6.445000 73.855000  6.645000 74.055000 ;
        RECT  6.445000 74.260000  6.645000 74.460000 ;
        RECT  6.445000 74.665000  6.645000 74.865000 ;
        RECT  6.445000 75.070000  6.645000 75.270000 ;
        RECT  6.445000 75.475000  6.645000 75.675000 ;
        RECT  6.445000 75.880000  6.645000 76.080000 ;
        RECT  6.445000 76.285000  6.645000 76.485000 ;
        RECT  6.445000 76.690000  6.645000 76.890000 ;
        RECT  6.445000 77.095000  6.645000 77.295000 ;
        RECT  6.445000 77.500000  6.645000 77.700000 ;
        RECT  6.445000 77.905000  6.645000 78.105000 ;
        RECT  6.445000 78.310000  6.645000 78.510000 ;
        RECT  6.445000 78.715000  6.645000 78.915000 ;
        RECT  6.445000 79.120000  6.645000 79.320000 ;
        RECT  6.445000 79.525000  6.645000 79.725000 ;
        RECT  6.445000 79.930000  6.645000 80.130000 ;
        RECT  6.445000 80.335000  6.645000 80.535000 ;
        RECT  6.445000 80.740000  6.645000 80.940000 ;
        RECT  6.445000 81.145000  6.645000 81.345000 ;
        RECT  6.445000 81.550000  6.645000 81.750000 ;
        RECT  6.445000 81.955000  6.645000 82.155000 ;
        RECT  6.445000 82.360000  6.645000 82.560000 ;
        RECT  6.475000 82.855000  6.675000 83.055000 ;
        RECT  6.475000 83.265000  6.675000 83.465000 ;
        RECT  6.475000 83.675000  6.675000 83.875000 ;
        RECT  6.475000 84.085000  6.675000 84.285000 ;
        RECT  6.475000 84.495000  6.675000 84.695000 ;
        RECT  6.475000 84.905000  6.675000 85.105000 ;
        RECT  6.475000 85.315000  6.675000 85.515000 ;
        RECT  6.475000 85.725000  6.675000 85.925000 ;
        RECT  6.475000 86.135000  6.675000 86.335000 ;
        RECT  6.475000 86.545000  6.675000 86.745000 ;
        RECT  6.475000 86.955000  6.675000 87.155000 ;
        RECT  6.475000 87.365000  6.675000 87.565000 ;
        RECT  6.475000 87.775000  6.675000 87.975000 ;
        RECT  6.475000 88.185000  6.675000 88.385000 ;
        RECT  6.475000 88.595000  6.675000 88.795000 ;
        RECT  6.475000 89.005000  6.675000 89.205000 ;
        RECT  6.475000 89.415000  6.675000 89.615000 ;
        RECT  6.475000 89.825000  6.675000 90.025000 ;
        RECT  6.475000 90.235000  6.675000 90.435000 ;
        RECT  6.475000 90.645000  6.675000 90.845000 ;
        RECT  6.475000 91.055000  6.675000 91.255000 ;
        RECT  6.475000 91.465000  6.675000 91.665000 ;
        RECT  6.475000 91.875000  6.675000 92.075000 ;
        RECT  6.475000 92.285000  6.675000 92.485000 ;
        RECT  6.475000 92.695000  6.675000 92.895000 ;
        RECT  6.765000 17.860000  6.965000 18.060000 ;
        RECT  6.765000 18.290000  6.965000 18.490000 ;
        RECT  6.765000 18.720000  6.965000 18.920000 ;
        RECT  6.765000 19.150000  6.965000 19.350000 ;
        RECT  6.765000 19.580000  6.965000 19.780000 ;
        RECT  6.765000 20.010000  6.965000 20.210000 ;
        RECT  6.765000 20.440000  6.965000 20.640000 ;
        RECT  6.765000 20.870000  6.965000 21.070000 ;
        RECT  6.765000 21.300000  6.965000 21.500000 ;
        RECT  6.765000 21.730000  6.965000 21.930000 ;
        RECT  6.765000 22.160000  6.965000 22.360000 ;
        RECT  6.845000 68.125000  7.045000 68.325000 ;
        RECT  6.845000 68.535000  7.045000 68.735000 ;
        RECT  6.845000 68.945000  7.045000 69.145000 ;
        RECT  6.845000 69.355000  7.045000 69.555000 ;
        RECT  6.845000 69.765000  7.045000 69.965000 ;
        RECT  6.845000 70.175000  7.045000 70.375000 ;
        RECT  6.845000 70.585000  7.045000 70.785000 ;
        RECT  6.845000 70.995000  7.045000 71.195000 ;
        RECT  6.845000 71.405000  7.045000 71.605000 ;
        RECT  6.845000 71.815000  7.045000 72.015000 ;
        RECT  6.845000 72.225000  7.045000 72.425000 ;
        RECT  6.845000 72.635000  7.045000 72.835000 ;
        RECT  6.845000 73.045000  7.045000 73.245000 ;
        RECT  6.845000 73.450000  7.045000 73.650000 ;
        RECT  6.845000 73.855000  7.045000 74.055000 ;
        RECT  6.845000 74.260000  7.045000 74.460000 ;
        RECT  6.845000 74.665000  7.045000 74.865000 ;
        RECT  6.845000 75.070000  7.045000 75.270000 ;
        RECT  6.845000 75.475000  7.045000 75.675000 ;
        RECT  6.845000 75.880000  7.045000 76.080000 ;
        RECT  6.845000 76.285000  7.045000 76.485000 ;
        RECT  6.845000 76.690000  7.045000 76.890000 ;
        RECT  6.845000 77.095000  7.045000 77.295000 ;
        RECT  6.845000 77.500000  7.045000 77.700000 ;
        RECT  6.845000 77.905000  7.045000 78.105000 ;
        RECT  6.845000 78.310000  7.045000 78.510000 ;
        RECT  6.845000 78.715000  7.045000 78.915000 ;
        RECT  6.845000 79.120000  7.045000 79.320000 ;
        RECT  6.845000 79.525000  7.045000 79.725000 ;
        RECT  6.845000 79.930000  7.045000 80.130000 ;
        RECT  6.845000 80.335000  7.045000 80.535000 ;
        RECT  6.845000 80.740000  7.045000 80.940000 ;
        RECT  6.845000 81.145000  7.045000 81.345000 ;
        RECT  6.845000 81.550000  7.045000 81.750000 ;
        RECT  6.845000 81.955000  7.045000 82.155000 ;
        RECT  6.845000 82.360000  7.045000 82.560000 ;
        RECT  6.885000 82.855000  7.085000 83.055000 ;
        RECT  6.885000 83.265000  7.085000 83.465000 ;
        RECT  6.885000 83.675000  7.085000 83.875000 ;
        RECT  6.885000 84.085000  7.085000 84.285000 ;
        RECT  6.885000 84.495000  7.085000 84.695000 ;
        RECT  6.885000 84.905000  7.085000 85.105000 ;
        RECT  6.885000 85.315000  7.085000 85.515000 ;
        RECT  6.885000 85.725000  7.085000 85.925000 ;
        RECT  6.885000 86.135000  7.085000 86.335000 ;
        RECT  6.885000 86.545000  7.085000 86.745000 ;
        RECT  6.885000 86.955000  7.085000 87.155000 ;
        RECT  6.885000 87.365000  7.085000 87.565000 ;
        RECT  6.885000 87.775000  7.085000 87.975000 ;
        RECT  6.885000 88.185000  7.085000 88.385000 ;
        RECT  6.885000 88.595000  7.085000 88.795000 ;
        RECT  6.885000 89.005000  7.085000 89.205000 ;
        RECT  6.885000 89.415000  7.085000 89.615000 ;
        RECT  6.885000 89.825000  7.085000 90.025000 ;
        RECT  6.885000 90.235000  7.085000 90.435000 ;
        RECT  6.885000 90.645000  7.085000 90.845000 ;
        RECT  6.885000 91.055000  7.085000 91.255000 ;
        RECT  6.885000 91.465000  7.085000 91.665000 ;
        RECT  6.885000 91.875000  7.085000 92.075000 ;
        RECT  6.885000 92.285000  7.085000 92.485000 ;
        RECT  6.885000 92.695000  7.085000 92.895000 ;
        RECT  7.170000 17.860000  7.370000 18.060000 ;
        RECT  7.170000 18.290000  7.370000 18.490000 ;
        RECT  7.170000 18.720000  7.370000 18.920000 ;
        RECT  7.170000 19.150000  7.370000 19.350000 ;
        RECT  7.170000 19.580000  7.370000 19.780000 ;
        RECT  7.170000 20.010000  7.370000 20.210000 ;
        RECT  7.170000 20.440000  7.370000 20.640000 ;
        RECT  7.170000 20.870000  7.370000 21.070000 ;
        RECT  7.170000 21.300000  7.370000 21.500000 ;
        RECT  7.170000 21.730000  7.370000 21.930000 ;
        RECT  7.170000 22.160000  7.370000 22.360000 ;
        RECT  7.245000 68.125000  7.445000 68.325000 ;
        RECT  7.245000 68.535000  7.445000 68.735000 ;
        RECT  7.245000 68.945000  7.445000 69.145000 ;
        RECT  7.245000 69.355000  7.445000 69.555000 ;
        RECT  7.245000 69.765000  7.445000 69.965000 ;
        RECT  7.245000 70.175000  7.445000 70.375000 ;
        RECT  7.245000 70.585000  7.445000 70.785000 ;
        RECT  7.245000 70.995000  7.445000 71.195000 ;
        RECT  7.245000 71.405000  7.445000 71.605000 ;
        RECT  7.245000 71.815000  7.445000 72.015000 ;
        RECT  7.245000 72.225000  7.445000 72.425000 ;
        RECT  7.245000 72.635000  7.445000 72.835000 ;
        RECT  7.245000 73.045000  7.445000 73.245000 ;
        RECT  7.245000 73.450000  7.445000 73.650000 ;
        RECT  7.245000 73.855000  7.445000 74.055000 ;
        RECT  7.245000 74.260000  7.445000 74.460000 ;
        RECT  7.245000 74.665000  7.445000 74.865000 ;
        RECT  7.245000 75.070000  7.445000 75.270000 ;
        RECT  7.245000 75.475000  7.445000 75.675000 ;
        RECT  7.245000 75.880000  7.445000 76.080000 ;
        RECT  7.245000 76.285000  7.445000 76.485000 ;
        RECT  7.245000 76.690000  7.445000 76.890000 ;
        RECT  7.245000 77.095000  7.445000 77.295000 ;
        RECT  7.245000 77.500000  7.445000 77.700000 ;
        RECT  7.245000 77.905000  7.445000 78.105000 ;
        RECT  7.245000 78.310000  7.445000 78.510000 ;
        RECT  7.245000 78.715000  7.445000 78.915000 ;
        RECT  7.245000 79.120000  7.445000 79.320000 ;
        RECT  7.245000 79.525000  7.445000 79.725000 ;
        RECT  7.245000 79.930000  7.445000 80.130000 ;
        RECT  7.245000 80.335000  7.445000 80.535000 ;
        RECT  7.245000 80.740000  7.445000 80.940000 ;
        RECT  7.245000 81.145000  7.445000 81.345000 ;
        RECT  7.245000 81.550000  7.445000 81.750000 ;
        RECT  7.245000 81.955000  7.445000 82.155000 ;
        RECT  7.245000 82.360000  7.445000 82.560000 ;
        RECT  7.295000 82.855000  7.495000 83.055000 ;
        RECT  7.295000 83.265000  7.495000 83.465000 ;
        RECT  7.295000 83.675000  7.495000 83.875000 ;
        RECT  7.295000 84.085000  7.495000 84.285000 ;
        RECT  7.295000 84.495000  7.495000 84.695000 ;
        RECT  7.295000 84.905000  7.495000 85.105000 ;
        RECT  7.295000 85.315000  7.495000 85.515000 ;
        RECT  7.295000 85.725000  7.495000 85.925000 ;
        RECT  7.295000 86.135000  7.495000 86.335000 ;
        RECT  7.295000 86.545000  7.495000 86.745000 ;
        RECT  7.295000 86.955000  7.495000 87.155000 ;
        RECT  7.295000 87.365000  7.495000 87.565000 ;
        RECT  7.295000 87.775000  7.495000 87.975000 ;
        RECT  7.295000 88.185000  7.495000 88.385000 ;
        RECT  7.295000 88.595000  7.495000 88.795000 ;
        RECT  7.295000 89.005000  7.495000 89.205000 ;
        RECT  7.295000 89.415000  7.495000 89.615000 ;
        RECT  7.295000 89.825000  7.495000 90.025000 ;
        RECT  7.295000 90.235000  7.495000 90.435000 ;
        RECT  7.295000 90.645000  7.495000 90.845000 ;
        RECT  7.295000 91.055000  7.495000 91.255000 ;
        RECT  7.295000 91.465000  7.495000 91.665000 ;
        RECT  7.295000 91.875000  7.495000 92.075000 ;
        RECT  7.295000 92.285000  7.495000 92.485000 ;
        RECT  7.295000 92.695000  7.495000 92.895000 ;
        RECT  7.575000 17.860000  7.775000 18.060000 ;
        RECT  7.575000 18.290000  7.775000 18.490000 ;
        RECT  7.575000 18.720000  7.775000 18.920000 ;
        RECT  7.575000 19.150000  7.775000 19.350000 ;
        RECT  7.575000 19.580000  7.775000 19.780000 ;
        RECT  7.575000 20.010000  7.775000 20.210000 ;
        RECT  7.575000 20.440000  7.775000 20.640000 ;
        RECT  7.575000 20.870000  7.775000 21.070000 ;
        RECT  7.575000 21.300000  7.775000 21.500000 ;
        RECT  7.575000 21.730000  7.775000 21.930000 ;
        RECT  7.575000 22.160000  7.775000 22.360000 ;
        RECT  7.645000 68.125000  7.845000 68.325000 ;
        RECT  7.645000 68.535000  7.845000 68.735000 ;
        RECT  7.645000 68.945000  7.845000 69.145000 ;
        RECT  7.645000 69.355000  7.845000 69.555000 ;
        RECT  7.645000 69.765000  7.845000 69.965000 ;
        RECT  7.645000 70.175000  7.845000 70.375000 ;
        RECT  7.645000 70.585000  7.845000 70.785000 ;
        RECT  7.645000 70.995000  7.845000 71.195000 ;
        RECT  7.645000 71.405000  7.845000 71.605000 ;
        RECT  7.645000 71.815000  7.845000 72.015000 ;
        RECT  7.645000 72.225000  7.845000 72.425000 ;
        RECT  7.645000 72.635000  7.845000 72.835000 ;
        RECT  7.645000 73.045000  7.845000 73.245000 ;
        RECT  7.645000 73.450000  7.845000 73.650000 ;
        RECT  7.645000 73.855000  7.845000 74.055000 ;
        RECT  7.645000 74.260000  7.845000 74.460000 ;
        RECT  7.645000 74.665000  7.845000 74.865000 ;
        RECT  7.645000 75.070000  7.845000 75.270000 ;
        RECT  7.645000 75.475000  7.845000 75.675000 ;
        RECT  7.645000 75.880000  7.845000 76.080000 ;
        RECT  7.645000 76.285000  7.845000 76.485000 ;
        RECT  7.645000 76.690000  7.845000 76.890000 ;
        RECT  7.645000 77.095000  7.845000 77.295000 ;
        RECT  7.645000 77.500000  7.845000 77.700000 ;
        RECT  7.645000 77.905000  7.845000 78.105000 ;
        RECT  7.645000 78.310000  7.845000 78.510000 ;
        RECT  7.645000 78.715000  7.845000 78.915000 ;
        RECT  7.645000 79.120000  7.845000 79.320000 ;
        RECT  7.645000 79.525000  7.845000 79.725000 ;
        RECT  7.645000 79.930000  7.845000 80.130000 ;
        RECT  7.645000 80.335000  7.845000 80.535000 ;
        RECT  7.645000 80.740000  7.845000 80.940000 ;
        RECT  7.645000 81.145000  7.845000 81.345000 ;
        RECT  7.645000 81.550000  7.845000 81.750000 ;
        RECT  7.645000 81.955000  7.845000 82.155000 ;
        RECT  7.645000 82.360000  7.845000 82.560000 ;
        RECT  7.705000 82.855000  7.905000 83.055000 ;
        RECT  7.705000 83.265000  7.905000 83.465000 ;
        RECT  7.705000 83.675000  7.905000 83.875000 ;
        RECT  7.705000 84.085000  7.905000 84.285000 ;
        RECT  7.705000 84.495000  7.905000 84.695000 ;
        RECT  7.705000 84.905000  7.905000 85.105000 ;
        RECT  7.705000 85.315000  7.905000 85.515000 ;
        RECT  7.705000 85.725000  7.905000 85.925000 ;
        RECT  7.705000 86.135000  7.905000 86.335000 ;
        RECT  7.705000 86.545000  7.905000 86.745000 ;
        RECT  7.705000 86.955000  7.905000 87.155000 ;
        RECT  7.705000 87.365000  7.905000 87.565000 ;
        RECT  7.705000 87.775000  7.905000 87.975000 ;
        RECT  7.705000 88.185000  7.905000 88.385000 ;
        RECT  7.705000 88.595000  7.905000 88.795000 ;
        RECT  7.705000 89.005000  7.905000 89.205000 ;
        RECT  7.705000 89.415000  7.905000 89.615000 ;
        RECT  7.705000 89.825000  7.905000 90.025000 ;
        RECT  7.705000 90.235000  7.905000 90.435000 ;
        RECT  7.705000 90.645000  7.905000 90.845000 ;
        RECT  7.705000 91.055000  7.905000 91.255000 ;
        RECT  7.705000 91.465000  7.905000 91.665000 ;
        RECT  7.705000 91.875000  7.905000 92.075000 ;
        RECT  7.705000 92.285000  7.905000 92.485000 ;
        RECT  7.705000 92.695000  7.905000 92.895000 ;
        RECT  7.980000 17.860000  8.180000 18.060000 ;
        RECT  7.980000 18.290000  8.180000 18.490000 ;
        RECT  7.980000 18.720000  8.180000 18.920000 ;
        RECT  7.980000 19.150000  8.180000 19.350000 ;
        RECT  7.980000 19.580000  8.180000 19.780000 ;
        RECT  7.980000 20.010000  8.180000 20.210000 ;
        RECT  7.980000 20.440000  8.180000 20.640000 ;
        RECT  7.980000 20.870000  8.180000 21.070000 ;
        RECT  7.980000 21.300000  8.180000 21.500000 ;
        RECT  7.980000 21.730000  8.180000 21.930000 ;
        RECT  7.980000 22.160000  8.180000 22.360000 ;
        RECT  8.045000 68.125000  8.245000 68.325000 ;
        RECT  8.045000 68.535000  8.245000 68.735000 ;
        RECT  8.045000 68.945000  8.245000 69.145000 ;
        RECT  8.045000 69.355000  8.245000 69.555000 ;
        RECT  8.045000 69.765000  8.245000 69.965000 ;
        RECT  8.045000 70.175000  8.245000 70.375000 ;
        RECT  8.045000 70.585000  8.245000 70.785000 ;
        RECT  8.045000 70.995000  8.245000 71.195000 ;
        RECT  8.045000 71.405000  8.245000 71.605000 ;
        RECT  8.045000 71.815000  8.245000 72.015000 ;
        RECT  8.045000 72.225000  8.245000 72.425000 ;
        RECT  8.045000 72.635000  8.245000 72.835000 ;
        RECT  8.045000 73.045000  8.245000 73.245000 ;
        RECT  8.045000 73.450000  8.245000 73.650000 ;
        RECT  8.045000 73.855000  8.245000 74.055000 ;
        RECT  8.045000 74.260000  8.245000 74.460000 ;
        RECT  8.045000 74.665000  8.245000 74.865000 ;
        RECT  8.045000 75.070000  8.245000 75.270000 ;
        RECT  8.045000 75.475000  8.245000 75.675000 ;
        RECT  8.045000 75.880000  8.245000 76.080000 ;
        RECT  8.045000 76.285000  8.245000 76.485000 ;
        RECT  8.045000 76.690000  8.245000 76.890000 ;
        RECT  8.045000 77.095000  8.245000 77.295000 ;
        RECT  8.045000 77.500000  8.245000 77.700000 ;
        RECT  8.045000 77.905000  8.245000 78.105000 ;
        RECT  8.045000 78.310000  8.245000 78.510000 ;
        RECT  8.045000 78.715000  8.245000 78.915000 ;
        RECT  8.045000 79.120000  8.245000 79.320000 ;
        RECT  8.045000 79.525000  8.245000 79.725000 ;
        RECT  8.045000 79.930000  8.245000 80.130000 ;
        RECT  8.045000 80.335000  8.245000 80.535000 ;
        RECT  8.045000 80.740000  8.245000 80.940000 ;
        RECT  8.045000 81.145000  8.245000 81.345000 ;
        RECT  8.045000 81.550000  8.245000 81.750000 ;
        RECT  8.045000 81.955000  8.245000 82.155000 ;
        RECT  8.045000 82.360000  8.245000 82.560000 ;
        RECT  8.115000 82.855000  8.315000 83.055000 ;
        RECT  8.115000 83.265000  8.315000 83.465000 ;
        RECT  8.115000 83.675000  8.315000 83.875000 ;
        RECT  8.115000 84.085000  8.315000 84.285000 ;
        RECT  8.115000 84.495000  8.315000 84.695000 ;
        RECT  8.115000 84.905000  8.315000 85.105000 ;
        RECT  8.115000 85.315000  8.315000 85.515000 ;
        RECT  8.115000 85.725000  8.315000 85.925000 ;
        RECT  8.115000 86.135000  8.315000 86.335000 ;
        RECT  8.115000 86.545000  8.315000 86.745000 ;
        RECT  8.115000 86.955000  8.315000 87.155000 ;
        RECT  8.115000 87.365000  8.315000 87.565000 ;
        RECT  8.115000 87.775000  8.315000 87.975000 ;
        RECT  8.115000 88.185000  8.315000 88.385000 ;
        RECT  8.115000 88.595000  8.315000 88.795000 ;
        RECT  8.115000 89.005000  8.315000 89.205000 ;
        RECT  8.115000 89.415000  8.315000 89.615000 ;
        RECT  8.115000 89.825000  8.315000 90.025000 ;
        RECT  8.115000 90.235000  8.315000 90.435000 ;
        RECT  8.115000 90.645000  8.315000 90.845000 ;
        RECT  8.115000 91.055000  8.315000 91.255000 ;
        RECT  8.115000 91.465000  8.315000 91.665000 ;
        RECT  8.115000 91.875000  8.315000 92.075000 ;
        RECT  8.115000 92.285000  8.315000 92.485000 ;
        RECT  8.115000 92.695000  8.315000 92.895000 ;
        RECT  8.385000 17.860000  8.585000 18.060000 ;
        RECT  8.385000 18.290000  8.585000 18.490000 ;
        RECT  8.385000 18.720000  8.585000 18.920000 ;
        RECT  8.385000 19.150000  8.585000 19.350000 ;
        RECT  8.385000 19.580000  8.585000 19.780000 ;
        RECT  8.385000 20.010000  8.585000 20.210000 ;
        RECT  8.385000 20.440000  8.585000 20.640000 ;
        RECT  8.385000 20.870000  8.585000 21.070000 ;
        RECT  8.385000 21.300000  8.585000 21.500000 ;
        RECT  8.385000 21.730000  8.585000 21.930000 ;
        RECT  8.385000 22.160000  8.585000 22.360000 ;
        RECT  8.445000 68.125000  8.645000 68.325000 ;
        RECT  8.445000 68.535000  8.645000 68.735000 ;
        RECT  8.445000 68.945000  8.645000 69.145000 ;
        RECT  8.445000 69.355000  8.645000 69.555000 ;
        RECT  8.445000 69.765000  8.645000 69.965000 ;
        RECT  8.445000 70.175000  8.645000 70.375000 ;
        RECT  8.445000 70.585000  8.645000 70.785000 ;
        RECT  8.445000 70.995000  8.645000 71.195000 ;
        RECT  8.445000 71.405000  8.645000 71.605000 ;
        RECT  8.445000 71.815000  8.645000 72.015000 ;
        RECT  8.445000 72.225000  8.645000 72.425000 ;
        RECT  8.445000 72.635000  8.645000 72.835000 ;
        RECT  8.445000 73.045000  8.645000 73.245000 ;
        RECT  8.445000 73.450000  8.645000 73.650000 ;
        RECT  8.445000 73.855000  8.645000 74.055000 ;
        RECT  8.445000 74.260000  8.645000 74.460000 ;
        RECT  8.445000 74.665000  8.645000 74.865000 ;
        RECT  8.445000 75.070000  8.645000 75.270000 ;
        RECT  8.445000 75.475000  8.645000 75.675000 ;
        RECT  8.445000 75.880000  8.645000 76.080000 ;
        RECT  8.445000 76.285000  8.645000 76.485000 ;
        RECT  8.445000 76.690000  8.645000 76.890000 ;
        RECT  8.445000 77.095000  8.645000 77.295000 ;
        RECT  8.445000 77.500000  8.645000 77.700000 ;
        RECT  8.445000 77.905000  8.645000 78.105000 ;
        RECT  8.445000 78.310000  8.645000 78.510000 ;
        RECT  8.445000 78.715000  8.645000 78.915000 ;
        RECT  8.445000 79.120000  8.645000 79.320000 ;
        RECT  8.445000 79.525000  8.645000 79.725000 ;
        RECT  8.445000 79.930000  8.645000 80.130000 ;
        RECT  8.445000 80.335000  8.645000 80.535000 ;
        RECT  8.445000 80.740000  8.645000 80.940000 ;
        RECT  8.445000 81.145000  8.645000 81.345000 ;
        RECT  8.445000 81.550000  8.645000 81.750000 ;
        RECT  8.445000 81.955000  8.645000 82.155000 ;
        RECT  8.445000 82.360000  8.645000 82.560000 ;
        RECT  8.525000 82.855000  8.725000 83.055000 ;
        RECT  8.525000 83.265000  8.725000 83.465000 ;
        RECT  8.525000 83.675000  8.725000 83.875000 ;
        RECT  8.525000 84.085000  8.725000 84.285000 ;
        RECT  8.525000 84.495000  8.725000 84.695000 ;
        RECT  8.525000 84.905000  8.725000 85.105000 ;
        RECT  8.525000 85.315000  8.725000 85.515000 ;
        RECT  8.525000 85.725000  8.725000 85.925000 ;
        RECT  8.525000 86.135000  8.725000 86.335000 ;
        RECT  8.525000 86.545000  8.725000 86.745000 ;
        RECT  8.525000 86.955000  8.725000 87.155000 ;
        RECT  8.525000 87.365000  8.725000 87.565000 ;
        RECT  8.525000 87.775000  8.725000 87.975000 ;
        RECT  8.525000 88.185000  8.725000 88.385000 ;
        RECT  8.525000 88.595000  8.725000 88.795000 ;
        RECT  8.525000 89.005000  8.725000 89.205000 ;
        RECT  8.525000 89.415000  8.725000 89.615000 ;
        RECT  8.525000 89.825000  8.725000 90.025000 ;
        RECT  8.525000 90.235000  8.725000 90.435000 ;
        RECT  8.525000 90.645000  8.725000 90.845000 ;
        RECT  8.525000 91.055000  8.725000 91.255000 ;
        RECT  8.525000 91.465000  8.725000 91.665000 ;
        RECT  8.525000 91.875000  8.725000 92.075000 ;
        RECT  8.525000 92.285000  8.725000 92.485000 ;
        RECT  8.525000 92.695000  8.725000 92.895000 ;
        RECT  8.790000 17.860000  8.990000 18.060000 ;
        RECT  8.790000 18.290000  8.990000 18.490000 ;
        RECT  8.790000 18.720000  8.990000 18.920000 ;
        RECT  8.790000 19.150000  8.990000 19.350000 ;
        RECT  8.790000 19.580000  8.990000 19.780000 ;
        RECT  8.790000 20.010000  8.990000 20.210000 ;
        RECT  8.790000 20.440000  8.990000 20.640000 ;
        RECT  8.790000 20.870000  8.990000 21.070000 ;
        RECT  8.790000 21.300000  8.990000 21.500000 ;
        RECT  8.790000 21.730000  8.990000 21.930000 ;
        RECT  8.790000 22.160000  8.990000 22.360000 ;
        RECT  8.845000 68.125000  9.045000 68.325000 ;
        RECT  8.845000 68.535000  9.045000 68.735000 ;
        RECT  8.845000 68.945000  9.045000 69.145000 ;
        RECT  8.845000 69.355000  9.045000 69.555000 ;
        RECT  8.845000 69.765000  9.045000 69.965000 ;
        RECT  8.845000 70.175000  9.045000 70.375000 ;
        RECT  8.845000 70.585000  9.045000 70.785000 ;
        RECT  8.845000 70.995000  9.045000 71.195000 ;
        RECT  8.845000 71.405000  9.045000 71.605000 ;
        RECT  8.845000 71.815000  9.045000 72.015000 ;
        RECT  8.845000 72.225000  9.045000 72.425000 ;
        RECT  8.845000 72.635000  9.045000 72.835000 ;
        RECT  8.845000 73.045000  9.045000 73.245000 ;
        RECT  8.845000 73.450000  9.045000 73.650000 ;
        RECT  8.845000 73.855000  9.045000 74.055000 ;
        RECT  8.845000 74.260000  9.045000 74.460000 ;
        RECT  8.845000 74.665000  9.045000 74.865000 ;
        RECT  8.845000 75.070000  9.045000 75.270000 ;
        RECT  8.845000 75.475000  9.045000 75.675000 ;
        RECT  8.845000 75.880000  9.045000 76.080000 ;
        RECT  8.845000 76.285000  9.045000 76.485000 ;
        RECT  8.845000 76.690000  9.045000 76.890000 ;
        RECT  8.845000 77.095000  9.045000 77.295000 ;
        RECT  8.845000 77.500000  9.045000 77.700000 ;
        RECT  8.845000 77.905000  9.045000 78.105000 ;
        RECT  8.845000 78.310000  9.045000 78.510000 ;
        RECT  8.845000 78.715000  9.045000 78.915000 ;
        RECT  8.845000 79.120000  9.045000 79.320000 ;
        RECT  8.845000 79.525000  9.045000 79.725000 ;
        RECT  8.845000 79.930000  9.045000 80.130000 ;
        RECT  8.845000 80.335000  9.045000 80.535000 ;
        RECT  8.845000 80.740000  9.045000 80.940000 ;
        RECT  8.845000 81.145000  9.045000 81.345000 ;
        RECT  8.845000 81.550000  9.045000 81.750000 ;
        RECT  8.845000 81.955000  9.045000 82.155000 ;
        RECT  8.845000 82.360000  9.045000 82.560000 ;
        RECT  8.935000 82.855000  9.135000 83.055000 ;
        RECT  8.935000 83.265000  9.135000 83.465000 ;
        RECT  8.935000 83.675000  9.135000 83.875000 ;
        RECT  8.935000 84.085000  9.135000 84.285000 ;
        RECT  8.935000 84.495000  9.135000 84.695000 ;
        RECT  8.935000 84.905000  9.135000 85.105000 ;
        RECT  8.935000 85.315000  9.135000 85.515000 ;
        RECT  8.935000 85.725000  9.135000 85.925000 ;
        RECT  8.935000 86.135000  9.135000 86.335000 ;
        RECT  8.935000 86.545000  9.135000 86.745000 ;
        RECT  8.935000 86.955000  9.135000 87.155000 ;
        RECT  8.935000 87.365000  9.135000 87.565000 ;
        RECT  8.935000 87.775000  9.135000 87.975000 ;
        RECT  8.935000 88.185000  9.135000 88.385000 ;
        RECT  8.935000 88.595000  9.135000 88.795000 ;
        RECT  8.935000 89.005000  9.135000 89.205000 ;
        RECT  8.935000 89.415000  9.135000 89.615000 ;
        RECT  8.935000 89.825000  9.135000 90.025000 ;
        RECT  8.935000 90.235000  9.135000 90.435000 ;
        RECT  8.935000 90.645000  9.135000 90.845000 ;
        RECT  8.935000 91.055000  9.135000 91.255000 ;
        RECT  8.935000 91.465000  9.135000 91.665000 ;
        RECT  8.935000 91.875000  9.135000 92.075000 ;
        RECT  8.935000 92.285000  9.135000 92.485000 ;
        RECT  8.935000 92.695000  9.135000 92.895000 ;
        RECT  9.195000 17.860000  9.395000 18.060000 ;
        RECT  9.195000 18.290000  9.395000 18.490000 ;
        RECT  9.195000 18.720000  9.395000 18.920000 ;
        RECT  9.195000 19.150000  9.395000 19.350000 ;
        RECT  9.195000 19.580000  9.395000 19.780000 ;
        RECT  9.195000 20.010000  9.395000 20.210000 ;
        RECT  9.195000 20.440000  9.395000 20.640000 ;
        RECT  9.195000 20.870000  9.395000 21.070000 ;
        RECT  9.195000 21.300000  9.395000 21.500000 ;
        RECT  9.195000 21.730000  9.395000 21.930000 ;
        RECT  9.195000 22.160000  9.395000 22.360000 ;
        RECT  9.245000 68.125000  9.445000 68.325000 ;
        RECT  9.245000 68.535000  9.445000 68.735000 ;
        RECT  9.245000 68.945000  9.445000 69.145000 ;
        RECT  9.245000 69.355000  9.445000 69.555000 ;
        RECT  9.245000 69.765000  9.445000 69.965000 ;
        RECT  9.245000 70.175000  9.445000 70.375000 ;
        RECT  9.245000 70.585000  9.445000 70.785000 ;
        RECT  9.245000 70.995000  9.445000 71.195000 ;
        RECT  9.245000 71.405000  9.445000 71.605000 ;
        RECT  9.245000 71.815000  9.445000 72.015000 ;
        RECT  9.245000 72.225000  9.445000 72.425000 ;
        RECT  9.245000 72.635000  9.445000 72.835000 ;
        RECT  9.245000 73.045000  9.445000 73.245000 ;
        RECT  9.245000 73.450000  9.445000 73.650000 ;
        RECT  9.245000 73.855000  9.445000 74.055000 ;
        RECT  9.245000 74.260000  9.445000 74.460000 ;
        RECT  9.245000 74.665000  9.445000 74.865000 ;
        RECT  9.245000 75.070000  9.445000 75.270000 ;
        RECT  9.245000 75.475000  9.445000 75.675000 ;
        RECT  9.245000 75.880000  9.445000 76.080000 ;
        RECT  9.245000 76.285000  9.445000 76.485000 ;
        RECT  9.245000 76.690000  9.445000 76.890000 ;
        RECT  9.245000 77.095000  9.445000 77.295000 ;
        RECT  9.245000 77.500000  9.445000 77.700000 ;
        RECT  9.245000 77.905000  9.445000 78.105000 ;
        RECT  9.245000 78.310000  9.445000 78.510000 ;
        RECT  9.245000 78.715000  9.445000 78.915000 ;
        RECT  9.245000 79.120000  9.445000 79.320000 ;
        RECT  9.245000 79.525000  9.445000 79.725000 ;
        RECT  9.245000 79.930000  9.445000 80.130000 ;
        RECT  9.245000 80.335000  9.445000 80.535000 ;
        RECT  9.245000 80.740000  9.445000 80.940000 ;
        RECT  9.245000 81.145000  9.445000 81.345000 ;
        RECT  9.245000 81.550000  9.445000 81.750000 ;
        RECT  9.245000 81.955000  9.445000 82.155000 ;
        RECT  9.245000 82.360000  9.445000 82.560000 ;
        RECT  9.345000 82.855000  9.545000 83.055000 ;
        RECT  9.345000 83.265000  9.545000 83.465000 ;
        RECT  9.345000 83.675000  9.545000 83.875000 ;
        RECT  9.345000 84.085000  9.545000 84.285000 ;
        RECT  9.345000 84.495000  9.545000 84.695000 ;
        RECT  9.345000 84.905000  9.545000 85.105000 ;
        RECT  9.345000 85.315000  9.545000 85.515000 ;
        RECT  9.345000 85.725000  9.545000 85.925000 ;
        RECT  9.345000 86.135000  9.545000 86.335000 ;
        RECT  9.345000 86.545000  9.545000 86.745000 ;
        RECT  9.345000 86.955000  9.545000 87.155000 ;
        RECT  9.345000 87.365000  9.545000 87.565000 ;
        RECT  9.345000 87.775000  9.545000 87.975000 ;
        RECT  9.345000 88.185000  9.545000 88.385000 ;
        RECT  9.345000 88.595000  9.545000 88.795000 ;
        RECT  9.345000 89.005000  9.545000 89.205000 ;
        RECT  9.345000 89.415000  9.545000 89.615000 ;
        RECT  9.345000 89.825000  9.545000 90.025000 ;
        RECT  9.345000 90.235000  9.545000 90.435000 ;
        RECT  9.345000 90.645000  9.545000 90.845000 ;
        RECT  9.345000 91.055000  9.545000 91.255000 ;
        RECT  9.345000 91.465000  9.545000 91.665000 ;
        RECT  9.345000 91.875000  9.545000 92.075000 ;
        RECT  9.345000 92.285000  9.545000 92.485000 ;
        RECT  9.345000 92.695000  9.545000 92.895000 ;
        RECT  9.600000 17.860000  9.800000 18.060000 ;
        RECT  9.600000 18.290000  9.800000 18.490000 ;
        RECT  9.600000 18.720000  9.800000 18.920000 ;
        RECT  9.600000 19.150000  9.800000 19.350000 ;
        RECT  9.600000 19.580000  9.800000 19.780000 ;
        RECT  9.600000 20.010000  9.800000 20.210000 ;
        RECT  9.600000 20.440000  9.800000 20.640000 ;
        RECT  9.600000 20.870000  9.800000 21.070000 ;
        RECT  9.600000 21.300000  9.800000 21.500000 ;
        RECT  9.600000 21.730000  9.800000 21.930000 ;
        RECT  9.600000 22.160000  9.800000 22.360000 ;
        RECT  9.645000 68.125000  9.845000 68.325000 ;
        RECT  9.645000 68.535000  9.845000 68.735000 ;
        RECT  9.645000 68.945000  9.845000 69.145000 ;
        RECT  9.645000 69.355000  9.845000 69.555000 ;
        RECT  9.645000 69.765000  9.845000 69.965000 ;
        RECT  9.645000 70.175000  9.845000 70.375000 ;
        RECT  9.645000 70.585000  9.845000 70.785000 ;
        RECT  9.645000 70.995000  9.845000 71.195000 ;
        RECT  9.645000 71.405000  9.845000 71.605000 ;
        RECT  9.645000 71.815000  9.845000 72.015000 ;
        RECT  9.645000 72.225000  9.845000 72.425000 ;
        RECT  9.645000 72.635000  9.845000 72.835000 ;
        RECT  9.645000 73.045000  9.845000 73.245000 ;
        RECT  9.645000 73.450000  9.845000 73.650000 ;
        RECT  9.645000 73.855000  9.845000 74.055000 ;
        RECT  9.645000 74.260000  9.845000 74.460000 ;
        RECT  9.645000 74.665000  9.845000 74.865000 ;
        RECT  9.645000 75.070000  9.845000 75.270000 ;
        RECT  9.645000 75.475000  9.845000 75.675000 ;
        RECT  9.645000 75.880000  9.845000 76.080000 ;
        RECT  9.645000 76.285000  9.845000 76.485000 ;
        RECT  9.645000 76.690000  9.845000 76.890000 ;
        RECT  9.645000 77.095000  9.845000 77.295000 ;
        RECT  9.645000 77.500000  9.845000 77.700000 ;
        RECT  9.645000 77.905000  9.845000 78.105000 ;
        RECT  9.645000 78.310000  9.845000 78.510000 ;
        RECT  9.645000 78.715000  9.845000 78.915000 ;
        RECT  9.645000 79.120000  9.845000 79.320000 ;
        RECT  9.645000 79.525000  9.845000 79.725000 ;
        RECT  9.645000 79.930000  9.845000 80.130000 ;
        RECT  9.645000 80.335000  9.845000 80.535000 ;
        RECT  9.645000 80.740000  9.845000 80.940000 ;
        RECT  9.645000 81.145000  9.845000 81.345000 ;
        RECT  9.645000 81.550000  9.845000 81.750000 ;
        RECT  9.645000 81.955000  9.845000 82.155000 ;
        RECT  9.645000 82.360000  9.845000 82.560000 ;
        RECT  9.755000 82.855000  9.955000 83.055000 ;
        RECT  9.755000 83.265000  9.955000 83.465000 ;
        RECT  9.755000 83.675000  9.955000 83.875000 ;
        RECT  9.755000 84.085000  9.955000 84.285000 ;
        RECT  9.755000 84.495000  9.955000 84.695000 ;
        RECT  9.755000 84.905000  9.955000 85.105000 ;
        RECT  9.755000 85.315000  9.955000 85.515000 ;
        RECT  9.755000 85.725000  9.955000 85.925000 ;
        RECT  9.755000 86.135000  9.955000 86.335000 ;
        RECT  9.755000 86.545000  9.955000 86.745000 ;
        RECT  9.755000 86.955000  9.955000 87.155000 ;
        RECT  9.755000 87.365000  9.955000 87.565000 ;
        RECT  9.755000 87.775000  9.955000 87.975000 ;
        RECT  9.755000 88.185000  9.955000 88.385000 ;
        RECT  9.755000 88.595000  9.955000 88.795000 ;
        RECT  9.755000 89.005000  9.955000 89.205000 ;
        RECT  9.755000 89.415000  9.955000 89.615000 ;
        RECT  9.755000 89.825000  9.955000 90.025000 ;
        RECT  9.755000 90.235000  9.955000 90.435000 ;
        RECT  9.755000 90.645000  9.955000 90.845000 ;
        RECT  9.755000 91.055000  9.955000 91.255000 ;
        RECT  9.755000 91.465000  9.955000 91.665000 ;
        RECT  9.755000 91.875000  9.955000 92.075000 ;
        RECT  9.755000 92.285000  9.955000 92.485000 ;
        RECT  9.755000 92.695000  9.955000 92.895000 ;
        RECT 10.005000 17.860000 10.205000 18.060000 ;
        RECT 10.005000 18.290000 10.205000 18.490000 ;
        RECT 10.005000 18.720000 10.205000 18.920000 ;
        RECT 10.005000 19.150000 10.205000 19.350000 ;
        RECT 10.005000 19.580000 10.205000 19.780000 ;
        RECT 10.005000 20.010000 10.205000 20.210000 ;
        RECT 10.005000 20.440000 10.205000 20.640000 ;
        RECT 10.005000 20.870000 10.205000 21.070000 ;
        RECT 10.005000 21.300000 10.205000 21.500000 ;
        RECT 10.005000 21.730000 10.205000 21.930000 ;
        RECT 10.005000 22.160000 10.205000 22.360000 ;
        RECT 10.045000 68.125000 10.245000 68.325000 ;
        RECT 10.045000 68.535000 10.245000 68.735000 ;
        RECT 10.045000 68.945000 10.245000 69.145000 ;
        RECT 10.045000 69.355000 10.245000 69.555000 ;
        RECT 10.045000 69.765000 10.245000 69.965000 ;
        RECT 10.045000 70.175000 10.245000 70.375000 ;
        RECT 10.045000 70.585000 10.245000 70.785000 ;
        RECT 10.045000 70.995000 10.245000 71.195000 ;
        RECT 10.045000 71.405000 10.245000 71.605000 ;
        RECT 10.045000 71.815000 10.245000 72.015000 ;
        RECT 10.045000 72.225000 10.245000 72.425000 ;
        RECT 10.045000 72.635000 10.245000 72.835000 ;
        RECT 10.045000 73.045000 10.245000 73.245000 ;
        RECT 10.045000 73.450000 10.245000 73.650000 ;
        RECT 10.045000 73.855000 10.245000 74.055000 ;
        RECT 10.045000 74.260000 10.245000 74.460000 ;
        RECT 10.045000 74.665000 10.245000 74.865000 ;
        RECT 10.045000 75.070000 10.245000 75.270000 ;
        RECT 10.045000 75.475000 10.245000 75.675000 ;
        RECT 10.045000 75.880000 10.245000 76.080000 ;
        RECT 10.045000 76.285000 10.245000 76.485000 ;
        RECT 10.045000 76.690000 10.245000 76.890000 ;
        RECT 10.045000 77.095000 10.245000 77.295000 ;
        RECT 10.045000 77.500000 10.245000 77.700000 ;
        RECT 10.045000 77.905000 10.245000 78.105000 ;
        RECT 10.045000 78.310000 10.245000 78.510000 ;
        RECT 10.045000 78.715000 10.245000 78.915000 ;
        RECT 10.045000 79.120000 10.245000 79.320000 ;
        RECT 10.045000 79.525000 10.245000 79.725000 ;
        RECT 10.045000 79.930000 10.245000 80.130000 ;
        RECT 10.045000 80.335000 10.245000 80.535000 ;
        RECT 10.045000 80.740000 10.245000 80.940000 ;
        RECT 10.045000 81.145000 10.245000 81.345000 ;
        RECT 10.045000 81.550000 10.245000 81.750000 ;
        RECT 10.045000 81.955000 10.245000 82.155000 ;
        RECT 10.045000 82.360000 10.245000 82.560000 ;
        RECT 10.165000 82.855000 10.365000 83.055000 ;
        RECT 10.165000 83.265000 10.365000 83.465000 ;
        RECT 10.165000 83.675000 10.365000 83.875000 ;
        RECT 10.165000 84.085000 10.365000 84.285000 ;
        RECT 10.165000 84.495000 10.365000 84.695000 ;
        RECT 10.165000 84.905000 10.365000 85.105000 ;
        RECT 10.165000 85.315000 10.365000 85.515000 ;
        RECT 10.165000 85.725000 10.365000 85.925000 ;
        RECT 10.165000 86.135000 10.365000 86.335000 ;
        RECT 10.165000 86.545000 10.365000 86.745000 ;
        RECT 10.165000 86.955000 10.365000 87.155000 ;
        RECT 10.165000 87.365000 10.365000 87.565000 ;
        RECT 10.165000 87.775000 10.365000 87.975000 ;
        RECT 10.165000 88.185000 10.365000 88.385000 ;
        RECT 10.165000 88.595000 10.365000 88.795000 ;
        RECT 10.165000 89.005000 10.365000 89.205000 ;
        RECT 10.165000 89.415000 10.365000 89.615000 ;
        RECT 10.165000 89.825000 10.365000 90.025000 ;
        RECT 10.165000 90.235000 10.365000 90.435000 ;
        RECT 10.165000 90.645000 10.365000 90.845000 ;
        RECT 10.165000 91.055000 10.365000 91.255000 ;
        RECT 10.165000 91.465000 10.365000 91.665000 ;
        RECT 10.165000 91.875000 10.365000 92.075000 ;
        RECT 10.165000 92.285000 10.365000 92.485000 ;
        RECT 10.165000 92.695000 10.365000 92.895000 ;
        RECT 10.410000 17.860000 10.610000 18.060000 ;
        RECT 10.410000 18.290000 10.610000 18.490000 ;
        RECT 10.410000 18.720000 10.610000 18.920000 ;
        RECT 10.410000 19.150000 10.610000 19.350000 ;
        RECT 10.410000 19.580000 10.610000 19.780000 ;
        RECT 10.410000 20.010000 10.610000 20.210000 ;
        RECT 10.410000 20.440000 10.610000 20.640000 ;
        RECT 10.410000 20.870000 10.610000 21.070000 ;
        RECT 10.410000 21.300000 10.610000 21.500000 ;
        RECT 10.410000 21.730000 10.610000 21.930000 ;
        RECT 10.410000 22.160000 10.610000 22.360000 ;
        RECT 10.445000 68.125000 10.645000 68.325000 ;
        RECT 10.445000 68.535000 10.645000 68.735000 ;
        RECT 10.445000 68.945000 10.645000 69.145000 ;
        RECT 10.445000 69.355000 10.645000 69.555000 ;
        RECT 10.445000 69.765000 10.645000 69.965000 ;
        RECT 10.445000 70.175000 10.645000 70.375000 ;
        RECT 10.445000 70.585000 10.645000 70.785000 ;
        RECT 10.445000 70.995000 10.645000 71.195000 ;
        RECT 10.445000 71.405000 10.645000 71.605000 ;
        RECT 10.445000 71.815000 10.645000 72.015000 ;
        RECT 10.445000 72.225000 10.645000 72.425000 ;
        RECT 10.445000 72.635000 10.645000 72.835000 ;
        RECT 10.445000 73.045000 10.645000 73.245000 ;
        RECT 10.445000 73.450000 10.645000 73.650000 ;
        RECT 10.445000 73.855000 10.645000 74.055000 ;
        RECT 10.445000 74.260000 10.645000 74.460000 ;
        RECT 10.445000 74.665000 10.645000 74.865000 ;
        RECT 10.445000 75.070000 10.645000 75.270000 ;
        RECT 10.445000 75.475000 10.645000 75.675000 ;
        RECT 10.445000 75.880000 10.645000 76.080000 ;
        RECT 10.445000 76.285000 10.645000 76.485000 ;
        RECT 10.445000 76.690000 10.645000 76.890000 ;
        RECT 10.445000 77.095000 10.645000 77.295000 ;
        RECT 10.445000 77.500000 10.645000 77.700000 ;
        RECT 10.445000 77.905000 10.645000 78.105000 ;
        RECT 10.445000 78.310000 10.645000 78.510000 ;
        RECT 10.445000 78.715000 10.645000 78.915000 ;
        RECT 10.445000 79.120000 10.645000 79.320000 ;
        RECT 10.445000 79.525000 10.645000 79.725000 ;
        RECT 10.445000 79.930000 10.645000 80.130000 ;
        RECT 10.445000 80.335000 10.645000 80.535000 ;
        RECT 10.445000 80.740000 10.645000 80.940000 ;
        RECT 10.445000 81.145000 10.645000 81.345000 ;
        RECT 10.445000 81.550000 10.645000 81.750000 ;
        RECT 10.445000 81.955000 10.645000 82.155000 ;
        RECT 10.445000 82.360000 10.645000 82.560000 ;
        RECT 10.575000 82.855000 10.775000 83.055000 ;
        RECT 10.575000 83.265000 10.775000 83.465000 ;
        RECT 10.575000 83.675000 10.775000 83.875000 ;
        RECT 10.575000 84.085000 10.775000 84.285000 ;
        RECT 10.575000 84.495000 10.775000 84.695000 ;
        RECT 10.575000 84.905000 10.775000 85.105000 ;
        RECT 10.575000 85.315000 10.775000 85.515000 ;
        RECT 10.575000 85.725000 10.775000 85.925000 ;
        RECT 10.575000 86.135000 10.775000 86.335000 ;
        RECT 10.575000 86.545000 10.775000 86.745000 ;
        RECT 10.575000 86.955000 10.775000 87.155000 ;
        RECT 10.575000 87.365000 10.775000 87.565000 ;
        RECT 10.575000 87.775000 10.775000 87.975000 ;
        RECT 10.575000 88.185000 10.775000 88.385000 ;
        RECT 10.575000 88.595000 10.775000 88.795000 ;
        RECT 10.575000 89.005000 10.775000 89.205000 ;
        RECT 10.575000 89.415000 10.775000 89.615000 ;
        RECT 10.575000 89.825000 10.775000 90.025000 ;
        RECT 10.575000 90.235000 10.775000 90.435000 ;
        RECT 10.575000 90.645000 10.775000 90.845000 ;
        RECT 10.575000 91.055000 10.775000 91.255000 ;
        RECT 10.575000 91.465000 10.775000 91.665000 ;
        RECT 10.575000 91.875000 10.775000 92.075000 ;
        RECT 10.575000 92.285000 10.775000 92.485000 ;
        RECT 10.575000 92.695000 10.775000 92.895000 ;
        RECT 10.815000 17.860000 11.015000 18.060000 ;
        RECT 10.815000 18.290000 11.015000 18.490000 ;
        RECT 10.815000 18.720000 11.015000 18.920000 ;
        RECT 10.815000 19.150000 11.015000 19.350000 ;
        RECT 10.815000 19.580000 11.015000 19.780000 ;
        RECT 10.815000 20.010000 11.015000 20.210000 ;
        RECT 10.815000 20.440000 11.015000 20.640000 ;
        RECT 10.815000 20.870000 11.015000 21.070000 ;
        RECT 10.815000 21.300000 11.015000 21.500000 ;
        RECT 10.815000 21.730000 11.015000 21.930000 ;
        RECT 10.815000 22.160000 11.015000 22.360000 ;
        RECT 10.845000 68.125000 11.045000 68.325000 ;
        RECT 10.845000 68.535000 11.045000 68.735000 ;
        RECT 10.845000 68.945000 11.045000 69.145000 ;
        RECT 10.845000 69.355000 11.045000 69.555000 ;
        RECT 10.845000 69.765000 11.045000 69.965000 ;
        RECT 10.845000 70.175000 11.045000 70.375000 ;
        RECT 10.845000 70.585000 11.045000 70.785000 ;
        RECT 10.845000 70.995000 11.045000 71.195000 ;
        RECT 10.845000 71.405000 11.045000 71.605000 ;
        RECT 10.845000 71.815000 11.045000 72.015000 ;
        RECT 10.845000 72.225000 11.045000 72.425000 ;
        RECT 10.845000 72.635000 11.045000 72.835000 ;
        RECT 10.845000 73.045000 11.045000 73.245000 ;
        RECT 10.845000 73.450000 11.045000 73.650000 ;
        RECT 10.845000 73.855000 11.045000 74.055000 ;
        RECT 10.845000 74.260000 11.045000 74.460000 ;
        RECT 10.845000 74.665000 11.045000 74.865000 ;
        RECT 10.845000 75.070000 11.045000 75.270000 ;
        RECT 10.845000 75.475000 11.045000 75.675000 ;
        RECT 10.845000 75.880000 11.045000 76.080000 ;
        RECT 10.845000 76.285000 11.045000 76.485000 ;
        RECT 10.845000 76.690000 11.045000 76.890000 ;
        RECT 10.845000 77.095000 11.045000 77.295000 ;
        RECT 10.845000 77.500000 11.045000 77.700000 ;
        RECT 10.845000 77.905000 11.045000 78.105000 ;
        RECT 10.845000 78.310000 11.045000 78.510000 ;
        RECT 10.845000 78.715000 11.045000 78.915000 ;
        RECT 10.845000 79.120000 11.045000 79.320000 ;
        RECT 10.845000 79.525000 11.045000 79.725000 ;
        RECT 10.845000 79.930000 11.045000 80.130000 ;
        RECT 10.845000 80.335000 11.045000 80.535000 ;
        RECT 10.845000 80.740000 11.045000 80.940000 ;
        RECT 10.845000 81.145000 11.045000 81.345000 ;
        RECT 10.845000 81.550000 11.045000 81.750000 ;
        RECT 10.845000 81.955000 11.045000 82.155000 ;
        RECT 10.845000 82.360000 11.045000 82.560000 ;
        RECT 10.985000 82.855000 11.185000 83.055000 ;
        RECT 10.985000 83.265000 11.185000 83.465000 ;
        RECT 10.985000 83.675000 11.185000 83.875000 ;
        RECT 10.985000 84.085000 11.185000 84.285000 ;
        RECT 10.985000 84.495000 11.185000 84.695000 ;
        RECT 10.985000 84.905000 11.185000 85.105000 ;
        RECT 10.985000 85.315000 11.185000 85.515000 ;
        RECT 10.985000 85.725000 11.185000 85.925000 ;
        RECT 10.985000 86.135000 11.185000 86.335000 ;
        RECT 10.985000 86.545000 11.185000 86.745000 ;
        RECT 10.985000 86.955000 11.185000 87.155000 ;
        RECT 10.985000 87.365000 11.185000 87.565000 ;
        RECT 10.985000 87.775000 11.185000 87.975000 ;
        RECT 10.985000 88.185000 11.185000 88.385000 ;
        RECT 10.985000 88.595000 11.185000 88.795000 ;
        RECT 10.985000 89.005000 11.185000 89.205000 ;
        RECT 10.985000 89.415000 11.185000 89.615000 ;
        RECT 10.985000 89.825000 11.185000 90.025000 ;
        RECT 10.985000 90.235000 11.185000 90.435000 ;
        RECT 10.985000 90.645000 11.185000 90.845000 ;
        RECT 10.985000 91.055000 11.185000 91.255000 ;
        RECT 10.985000 91.465000 11.185000 91.665000 ;
        RECT 10.985000 91.875000 11.185000 92.075000 ;
        RECT 10.985000 92.285000 11.185000 92.485000 ;
        RECT 10.985000 92.695000 11.185000 92.895000 ;
        RECT 11.220000 17.860000 11.420000 18.060000 ;
        RECT 11.220000 18.290000 11.420000 18.490000 ;
        RECT 11.220000 18.720000 11.420000 18.920000 ;
        RECT 11.220000 19.150000 11.420000 19.350000 ;
        RECT 11.220000 19.580000 11.420000 19.780000 ;
        RECT 11.220000 20.010000 11.420000 20.210000 ;
        RECT 11.220000 20.440000 11.420000 20.640000 ;
        RECT 11.220000 20.870000 11.420000 21.070000 ;
        RECT 11.220000 21.300000 11.420000 21.500000 ;
        RECT 11.220000 21.730000 11.420000 21.930000 ;
        RECT 11.220000 22.160000 11.420000 22.360000 ;
        RECT 11.245000 68.125000 11.445000 68.325000 ;
        RECT 11.245000 68.535000 11.445000 68.735000 ;
        RECT 11.245000 68.945000 11.445000 69.145000 ;
        RECT 11.245000 69.355000 11.445000 69.555000 ;
        RECT 11.245000 69.765000 11.445000 69.965000 ;
        RECT 11.245000 70.175000 11.445000 70.375000 ;
        RECT 11.245000 70.585000 11.445000 70.785000 ;
        RECT 11.245000 70.995000 11.445000 71.195000 ;
        RECT 11.245000 71.405000 11.445000 71.605000 ;
        RECT 11.245000 71.815000 11.445000 72.015000 ;
        RECT 11.245000 72.225000 11.445000 72.425000 ;
        RECT 11.245000 72.635000 11.445000 72.835000 ;
        RECT 11.245000 73.045000 11.445000 73.245000 ;
        RECT 11.245000 73.450000 11.445000 73.650000 ;
        RECT 11.245000 73.855000 11.445000 74.055000 ;
        RECT 11.245000 74.260000 11.445000 74.460000 ;
        RECT 11.245000 74.665000 11.445000 74.865000 ;
        RECT 11.245000 75.070000 11.445000 75.270000 ;
        RECT 11.245000 75.475000 11.445000 75.675000 ;
        RECT 11.245000 75.880000 11.445000 76.080000 ;
        RECT 11.245000 76.285000 11.445000 76.485000 ;
        RECT 11.245000 76.690000 11.445000 76.890000 ;
        RECT 11.245000 77.095000 11.445000 77.295000 ;
        RECT 11.245000 77.500000 11.445000 77.700000 ;
        RECT 11.245000 77.905000 11.445000 78.105000 ;
        RECT 11.245000 78.310000 11.445000 78.510000 ;
        RECT 11.245000 78.715000 11.445000 78.915000 ;
        RECT 11.245000 79.120000 11.445000 79.320000 ;
        RECT 11.245000 79.525000 11.445000 79.725000 ;
        RECT 11.245000 79.930000 11.445000 80.130000 ;
        RECT 11.245000 80.335000 11.445000 80.535000 ;
        RECT 11.245000 80.740000 11.445000 80.940000 ;
        RECT 11.245000 81.145000 11.445000 81.345000 ;
        RECT 11.245000 81.550000 11.445000 81.750000 ;
        RECT 11.245000 81.955000 11.445000 82.155000 ;
        RECT 11.245000 82.360000 11.445000 82.560000 ;
        RECT 11.395000 82.855000 11.595000 83.055000 ;
        RECT 11.395000 83.265000 11.595000 83.465000 ;
        RECT 11.395000 83.675000 11.595000 83.875000 ;
        RECT 11.395000 84.085000 11.595000 84.285000 ;
        RECT 11.395000 84.495000 11.595000 84.695000 ;
        RECT 11.395000 84.905000 11.595000 85.105000 ;
        RECT 11.395000 85.315000 11.595000 85.515000 ;
        RECT 11.395000 85.725000 11.595000 85.925000 ;
        RECT 11.395000 86.135000 11.595000 86.335000 ;
        RECT 11.395000 86.545000 11.595000 86.745000 ;
        RECT 11.395000 86.955000 11.595000 87.155000 ;
        RECT 11.395000 87.365000 11.595000 87.565000 ;
        RECT 11.395000 87.775000 11.595000 87.975000 ;
        RECT 11.395000 88.185000 11.595000 88.385000 ;
        RECT 11.395000 88.595000 11.595000 88.795000 ;
        RECT 11.395000 89.005000 11.595000 89.205000 ;
        RECT 11.395000 89.415000 11.595000 89.615000 ;
        RECT 11.395000 89.825000 11.595000 90.025000 ;
        RECT 11.395000 90.235000 11.595000 90.435000 ;
        RECT 11.395000 90.645000 11.595000 90.845000 ;
        RECT 11.395000 91.055000 11.595000 91.255000 ;
        RECT 11.395000 91.465000 11.595000 91.665000 ;
        RECT 11.395000 91.875000 11.595000 92.075000 ;
        RECT 11.395000 92.285000 11.595000 92.485000 ;
        RECT 11.395000 92.695000 11.595000 92.895000 ;
        RECT 11.625000 17.860000 11.825000 18.060000 ;
        RECT 11.625000 18.290000 11.825000 18.490000 ;
        RECT 11.625000 18.720000 11.825000 18.920000 ;
        RECT 11.625000 19.150000 11.825000 19.350000 ;
        RECT 11.625000 19.580000 11.825000 19.780000 ;
        RECT 11.625000 20.010000 11.825000 20.210000 ;
        RECT 11.625000 20.440000 11.825000 20.640000 ;
        RECT 11.625000 20.870000 11.825000 21.070000 ;
        RECT 11.625000 21.300000 11.825000 21.500000 ;
        RECT 11.625000 21.730000 11.825000 21.930000 ;
        RECT 11.625000 22.160000 11.825000 22.360000 ;
        RECT 11.645000 68.125000 11.845000 68.325000 ;
        RECT 11.645000 68.535000 11.845000 68.735000 ;
        RECT 11.645000 68.945000 11.845000 69.145000 ;
        RECT 11.645000 69.355000 11.845000 69.555000 ;
        RECT 11.645000 69.765000 11.845000 69.965000 ;
        RECT 11.645000 70.175000 11.845000 70.375000 ;
        RECT 11.645000 70.585000 11.845000 70.785000 ;
        RECT 11.645000 70.995000 11.845000 71.195000 ;
        RECT 11.645000 71.405000 11.845000 71.605000 ;
        RECT 11.645000 71.815000 11.845000 72.015000 ;
        RECT 11.645000 72.225000 11.845000 72.425000 ;
        RECT 11.645000 72.635000 11.845000 72.835000 ;
        RECT 11.645000 73.045000 11.845000 73.245000 ;
        RECT 11.645000 73.450000 11.845000 73.650000 ;
        RECT 11.645000 73.855000 11.845000 74.055000 ;
        RECT 11.645000 74.260000 11.845000 74.460000 ;
        RECT 11.645000 74.665000 11.845000 74.865000 ;
        RECT 11.645000 75.070000 11.845000 75.270000 ;
        RECT 11.645000 75.475000 11.845000 75.675000 ;
        RECT 11.645000 75.880000 11.845000 76.080000 ;
        RECT 11.645000 76.285000 11.845000 76.485000 ;
        RECT 11.645000 76.690000 11.845000 76.890000 ;
        RECT 11.645000 77.095000 11.845000 77.295000 ;
        RECT 11.645000 77.500000 11.845000 77.700000 ;
        RECT 11.645000 77.905000 11.845000 78.105000 ;
        RECT 11.645000 78.310000 11.845000 78.510000 ;
        RECT 11.645000 78.715000 11.845000 78.915000 ;
        RECT 11.645000 79.120000 11.845000 79.320000 ;
        RECT 11.645000 79.525000 11.845000 79.725000 ;
        RECT 11.645000 79.930000 11.845000 80.130000 ;
        RECT 11.645000 80.335000 11.845000 80.535000 ;
        RECT 11.645000 80.740000 11.845000 80.940000 ;
        RECT 11.645000 81.145000 11.845000 81.345000 ;
        RECT 11.645000 81.550000 11.845000 81.750000 ;
        RECT 11.645000 81.955000 11.845000 82.155000 ;
        RECT 11.645000 82.360000 11.845000 82.560000 ;
        RECT 11.805000 82.855000 12.005000 83.055000 ;
        RECT 11.805000 83.265000 12.005000 83.465000 ;
        RECT 11.805000 83.675000 12.005000 83.875000 ;
        RECT 11.805000 84.085000 12.005000 84.285000 ;
        RECT 11.805000 84.495000 12.005000 84.695000 ;
        RECT 11.805000 84.905000 12.005000 85.105000 ;
        RECT 11.805000 85.315000 12.005000 85.515000 ;
        RECT 11.805000 85.725000 12.005000 85.925000 ;
        RECT 11.805000 86.135000 12.005000 86.335000 ;
        RECT 11.805000 86.545000 12.005000 86.745000 ;
        RECT 11.805000 86.955000 12.005000 87.155000 ;
        RECT 11.805000 87.365000 12.005000 87.565000 ;
        RECT 11.805000 87.775000 12.005000 87.975000 ;
        RECT 11.805000 88.185000 12.005000 88.385000 ;
        RECT 11.805000 88.595000 12.005000 88.795000 ;
        RECT 11.805000 89.005000 12.005000 89.205000 ;
        RECT 11.805000 89.415000 12.005000 89.615000 ;
        RECT 11.805000 89.825000 12.005000 90.025000 ;
        RECT 11.805000 90.235000 12.005000 90.435000 ;
        RECT 11.805000 90.645000 12.005000 90.845000 ;
        RECT 11.805000 91.055000 12.005000 91.255000 ;
        RECT 11.805000 91.465000 12.005000 91.665000 ;
        RECT 11.805000 91.875000 12.005000 92.075000 ;
        RECT 11.805000 92.285000 12.005000 92.485000 ;
        RECT 11.805000 92.695000 12.005000 92.895000 ;
        RECT 12.030000 17.860000 12.230000 18.060000 ;
        RECT 12.030000 18.290000 12.230000 18.490000 ;
        RECT 12.030000 18.720000 12.230000 18.920000 ;
        RECT 12.030000 19.150000 12.230000 19.350000 ;
        RECT 12.030000 19.580000 12.230000 19.780000 ;
        RECT 12.030000 20.010000 12.230000 20.210000 ;
        RECT 12.030000 20.440000 12.230000 20.640000 ;
        RECT 12.030000 20.870000 12.230000 21.070000 ;
        RECT 12.030000 21.300000 12.230000 21.500000 ;
        RECT 12.030000 21.730000 12.230000 21.930000 ;
        RECT 12.030000 22.160000 12.230000 22.360000 ;
        RECT 12.045000 68.125000 12.245000 68.325000 ;
        RECT 12.045000 68.535000 12.245000 68.735000 ;
        RECT 12.045000 68.945000 12.245000 69.145000 ;
        RECT 12.045000 69.355000 12.245000 69.555000 ;
        RECT 12.045000 69.765000 12.245000 69.965000 ;
        RECT 12.045000 70.175000 12.245000 70.375000 ;
        RECT 12.045000 70.585000 12.245000 70.785000 ;
        RECT 12.045000 70.995000 12.245000 71.195000 ;
        RECT 12.045000 71.405000 12.245000 71.605000 ;
        RECT 12.045000 71.815000 12.245000 72.015000 ;
        RECT 12.045000 72.225000 12.245000 72.425000 ;
        RECT 12.045000 72.635000 12.245000 72.835000 ;
        RECT 12.045000 73.045000 12.245000 73.245000 ;
        RECT 12.045000 73.450000 12.245000 73.650000 ;
        RECT 12.045000 73.855000 12.245000 74.055000 ;
        RECT 12.045000 74.260000 12.245000 74.460000 ;
        RECT 12.045000 74.665000 12.245000 74.865000 ;
        RECT 12.045000 75.070000 12.245000 75.270000 ;
        RECT 12.045000 75.475000 12.245000 75.675000 ;
        RECT 12.045000 75.880000 12.245000 76.080000 ;
        RECT 12.045000 76.285000 12.245000 76.485000 ;
        RECT 12.045000 76.690000 12.245000 76.890000 ;
        RECT 12.045000 77.095000 12.245000 77.295000 ;
        RECT 12.045000 77.500000 12.245000 77.700000 ;
        RECT 12.045000 77.905000 12.245000 78.105000 ;
        RECT 12.045000 78.310000 12.245000 78.510000 ;
        RECT 12.045000 78.715000 12.245000 78.915000 ;
        RECT 12.045000 79.120000 12.245000 79.320000 ;
        RECT 12.045000 79.525000 12.245000 79.725000 ;
        RECT 12.045000 79.930000 12.245000 80.130000 ;
        RECT 12.045000 80.335000 12.245000 80.535000 ;
        RECT 12.045000 80.740000 12.245000 80.940000 ;
        RECT 12.045000 81.145000 12.245000 81.345000 ;
        RECT 12.045000 81.550000 12.245000 81.750000 ;
        RECT 12.045000 81.955000 12.245000 82.155000 ;
        RECT 12.045000 82.360000 12.245000 82.560000 ;
        RECT 12.215000 82.855000 12.415000 83.055000 ;
        RECT 12.215000 83.265000 12.415000 83.465000 ;
        RECT 12.215000 83.675000 12.415000 83.875000 ;
        RECT 12.215000 84.085000 12.415000 84.285000 ;
        RECT 12.215000 84.495000 12.415000 84.695000 ;
        RECT 12.215000 84.905000 12.415000 85.105000 ;
        RECT 12.215000 85.315000 12.415000 85.515000 ;
        RECT 12.215000 85.725000 12.415000 85.925000 ;
        RECT 12.215000 86.135000 12.415000 86.335000 ;
        RECT 12.215000 86.545000 12.415000 86.745000 ;
        RECT 12.215000 86.955000 12.415000 87.155000 ;
        RECT 12.215000 87.365000 12.415000 87.565000 ;
        RECT 12.215000 87.775000 12.415000 87.975000 ;
        RECT 12.215000 88.185000 12.415000 88.385000 ;
        RECT 12.215000 88.595000 12.415000 88.795000 ;
        RECT 12.215000 89.005000 12.415000 89.205000 ;
        RECT 12.215000 89.415000 12.415000 89.615000 ;
        RECT 12.215000 89.825000 12.415000 90.025000 ;
        RECT 12.215000 90.235000 12.415000 90.435000 ;
        RECT 12.215000 90.645000 12.415000 90.845000 ;
        RECT 12.215000 91.055000 12.415000 91.255000 ;
        RECT 12.215000 91.465000 12.415000 91.665000 ;
        RECT 12.215000 91.875000 12.415000 92.075000 ;
        RECT 12.215000 92.285000 12.415000 92.485000 ;
        RECT 12.215000 92.695000 12.415000 92.895000 ;
        RECT 12.435000 17.860000 12.635000 18.060000 ;
        RECT 12.435000 18.290000 12.635000 18.490000 ;
        RECT 12.435000 18.720000 12.635000 18.920000 ;
        RECT 12.435000 19.150000 12.635000 19.350000 ;
        RECT 12.435000 19.580000 12.635000 19.780000 ;
        RECT 12.435000 20.010000 12.635000 20.210000 ;
        RECT 12.435000 20.440000 12.635000 20.640000 ;
        RECT 12.435000 20.870000 12.635000 21.070000 ;
        RECT 12.435000 21.300000 12.635000 21.500000 ;
        RECT 12.435000 21.730000 12.635000 21.930000 ;
        RECT 12.435000 22.160000 12.635000 22.360000 ;
        RECT 12.445000 68.125000 12.645000 68.325000 ;
        RECT 12.445000 68.535000 12.645000 68.735000 ;
        RECT 12.445000 68.945000 12.645000 69.145000 ;
        RECT 12.445000 69.355000 12.645000 69.555000 ;
        RECT 12.445000 69.765000 12.645000 69.965000 ;
        RECT 12.445000 70.175000 12.645000 70.375000 ;
        RECT 12.445000 70.585000 12.645000 70.785000 ;
        RECT 12.445000 70.995000 12.645000 71.195000 ;
        RECT 12.445000 71.405000 12.645000 71.605000 ;
        RECT 12.445000 71.815000 12.645000 72.015000 ;
        RECT 12.445000 72.225000 12.645000 72.425000 ;
        RECT 12.445000 72.635000 12.645000 72.835000 ;
        RECT 12.445000 73.045000 12.645000 73.245000 ;
        RECT 12.445000 73.450000 12.645000 73.650000 ;
        RECT 12.445000 73.855000 12.645000 74.055000 ;
        RECT 12.445000 74.260000 12.645000 74.460000 ;
        RECT 12.445000 74.665000 12.645000 74.865000 ;
        RECT 12.445000 75.070000 12.645000 75.270000 ;
        RECT 12.445000 75.475000 12.645000 75.675000 ;
        RECT 12.445000 75.880000 12.645000 76.080000 ;
        RECT 12.445000 76.285000 12.645000 76.485000 ;
        RECT 12.445000 76.690000 12.645000 76.890000 ;
        RECT 12.445000 77.095000 12.645000 77.295000 ;
        RECT 12.445000 77.500000 12.645000 77.700000 ;
        RECT 12.445000 77.905000 12.645000 78.105000 ;
        RECT 12.445000 78.310000 12.645000 78.510000 ;
        RECT 12.445000 78.715000 12.645000 78.915000 ;
        RECT 12.445000 79.120000 12.645000 79.320000 ;
        RECT 12.445000 79.525000 12.645000 79.725000 ;
        RECT 12.445000 79.930000 12.645000 80.130000 ;
        RECT 12.445000 80.335000 12.645000 80.535000 ;
        RECT 12.445000 80.740000 12.645000 80.940000 ;
        RECT 12.445000 81.145000 12.645000 81.345000 ;
        RECT 12.445000 81.550000 12.645000 81.750000 ;
        RECT 12.445000 81.955000 12.645000 82.155000 ;
        RECT 12.445000 82.360000 12.645000 82.560000 ;
        RECT 12.625000 82.855000 12.825000 83.055000 ;
        RECT 12.625000 83.265000 12.825000 83.465000 ;
        RECT 12.625000 83.675000 12.825000 83.875000 ;
        RECT 12.625000 84.085000 12.825000 84.285000 ;
        RECT 12.625000 84.495000 12.825000 84.695000 ;
        RECT 12.625000 84.905000 12.825000 85.105000 ;
        RECT 12.625000 85.315000 12.825000 85.515000 ;
        RECT 12.625000 85.725000 12.825000 85.925000 ;
        RECT 12.625000 86.135000 12.825000 86.335000 ;
        RECT 12.625000 86.545000 12.825000 86.745000 ;
        RECT 12.625000 86.955000 12.825000 87.155000 ;
        RECT 12.625000 87.365000 12.825000 87.565000 ;
        RECT 12.625000 87.775000 12.825000 87.975000 ;
        RECT 12.625000 88.185000 12.825000 88.385000 ;
        RECT 12.625000 88.595000 12.825000 88.795000 ;
        RECT 12.625000 89.005000 12.825000 89.205000 ;
        RECT 12.625000 89.415000 12.825000 89.615000 ;
        RECT 12.625000 89.825000 12.825000 90.025000 ;
        RECT 12.625000 90.235000 12.825000 90.435000 ;
        RECT 12.625000 90.645000 12.825000 90.845000 ;
        RECT 12.625000 91.055000 12.825000 91.255000 ;
        RECT 12.625000 91.465000 12.825000 91.665000 ;
        RECT 12.625000 91.875000 12.825000 92.075000 ;
        RECT 12.625000 92.285000 12.825000 92.485000 ;
        RECT 12.625000 92.695000 12.825000 92.895000 ;
        RECT 12.840000 17.860000 13.040000 18.060000 ;
        RECT 12.840000 18.290000 13.040000 18.490000 ;
        RECT 12.840000 18.720000 13.040000 18.920000 ;
        RECT 12.840000 19.150000 13.040000 19.350000 ;
        RECT 12.840000 19.580000 13.040000 19.780000 ;
        RECT 12.840000 20.010000 13.040000 20.210000 ;
        RECT 12.840000 20.440000 13.040000 20.640000 ;
        RECT 12.840000 20.870000 13.040000 21.070000 ;
        RECT 12.840000 21.300000 13.040000 21.500000 ;
        RECT 12.840000 21.730000 13.040000 21.930000 ;
        RECT 12.840000 22.160000 13.040000 22.360000 ;
        RECT 12.845000 68.125000 13.045000 68.325000 ;
        RECT 12.845000 68.535000 13.045000 68.735000 ;
        RECT 12.845000 68.945000 13.045000 69.145000 ;
        RECT 12.845000 69.355000 13.045000 69.555000 ;
        RECT 12.845000 69.765000 13.045000 69.965000 ;
        RECT 12.845000 70.175000 13.045000 70.375000 ;
        RECT 12.845000 70.585000 13.045000 70.785000 ;
        RECT 12.845000 70.995000 13.045000 71.195000 ;
        RECT 12.845000 71.405000 13.045000 71.605000 ;
        RECT 12.845000 71.815000 13.045000 72.015000 ;
        RECT 12.845000 72.225000 13.045000 72.425000 ;
        RECT 12.845000 72.635000 13.045000 72.835000 ;
        RECT 12.845000 73.045000 13.045000 73.245000 ;
        RECT 12.845000 73.450000 13.045000 73.650000 ;
        RECT 12.845000 73.855000 13.045000 74.055000 ;
        RECT 12.845000 74.260000 13.045000 74.460000 ;
        RECT 12.845000 74.665000 13.045000 74.865000 ;
        RECT 12.845000 75.070000 13.045000 75.270000 ;
        RECT 12.845000 75.475000 13.045000 75.675000 ;
        RECT 12.845000 75.880000 13.045000 76.080000 ;
        RECT 12.845000 76.285000 13.045000 76.485000 ;
        RECT 12.845000 76.690000 13.045000 76.890000 ;
        RECT 12.845000 77.095000 13.045000 77.295000 ;
        RECT 12.845000 77.500000 13.045000 77.700000 ;
        RECT 12.845000 77.905000 13.045000 78.105000 ;
        RECT 12.845000 78.310000 13.045000 78.510000 ;
        RECT 12.845000 78.715000 13.045000 78.915000 ;
        RECT 12.845000 79.120000 13.045000 79.320000 ;
        RECT 12.845000 79.525000 13.045000 79.725000 ;
        RECT 12.845000 79.930000 13.045000 80.130000 ;
        RECT 12.845000 80.335000 13.045000 80.535000 ;
        RECT 12.845000 80.740000 13.045000 80.940000 ;
        RECT 12.845000 81.145000 13.045000 81.345000 ;
        RECT 12.845000 81.550000 13.045000 81.750000 ;
        RECT 12.845000 81.955000 13.045000 82.155000 ;
        RECT 12.845000 82.360000 13.045000 82.560000 ;
        RECT 13.030000 82.855000 13.230000 83.055000 ;
        RECT 13.030000 83.265000 13.230000 83.465000 ;
        RECT 13.030000 83.675000 13.230000 83.875000 ;
        RECT 13.030000 84.085000 13.230000 84.285000 ;
        RECT 13.030000 84.495000 13.230000 84.695000 ;
        RECT 13.030000 84.905000 13.230000 85.105000 ;
        RECT 13.030000 85.315000 13.230000 85.515000 ;
        RECT 13.030000 85.725000 13.230000 85.925000 ;
        RECT 13.030000 86.135000 13.230000 86.335000 ;
        RECT 13.030000 86.545000 13.230000 86.745000 ;
        RECT 13.030000 86.955000 13.230000 87.155000 ;
        RECT 13.030000 87.365000 13.230000 87.565000 ;
        RECT 13.030000 87.775000 13.230000 87.975000 ;
        RECT 13.030000 88.185000 13.230000 88.385000 ;
        RECT 13.030000 88.595000 13.230000 88.795000 ;
        RECT 13.030000 89.005000 13.230000 89.205000 ;
        RECT 13.030000 89.415000 13.230000 89.615000 ;
        RECT 13.030000 89.825000 13.230000 90.025000 ;
        RECT 13.030000 90.235000 13.230000 90.435000 ;
        RECT 13.030000 90.645000 13.230000 90.845000 ;
        RECT 13.030000 91.055000 13.230000 91.255000 ;
        RECT 13.030000 91.465000 13.230000 91.665000 ;
        RECT 13.030000 91.875000 13.230000 92.075000 ;
        RECT 13.030000 92.285000 13.230000 92.485000 ;
        RECT 13.030000 92.695000 13.230000 92.895000 ;
        RECT 13.245000 17.860000 13.445000 18.060000 ;
        RECT 13.245000 18.290000 13.445000 18.490000 ;
        RECT 13.245000 18.720000 13.445000 18.920000 ;
        RECT 13.245000 19.150000 13.445000 19.350000 ;
        RECT 13.245000 19.580000 13.445000 19.780000 ;
        RECT 13.245000 20.010000 13.445000 20.210000 ;
        RECT 13.245000 20.440000 13.445000 20.640000 ;
        RECT 13.245000 20.870000 13.445000 21.070000 ;
        RECT 13.245000 21.300000 13.445000 21.500000 ;
        RECT 13.245000 21.730000 13.445000 21.930000 ;
        RECT 13.245000 22.160000 13.445000 22.360000 ;
        RECT 13.245000 68.125000 13.445000 68.325000 ;
        RECT 13.245000 68.535000 13.445000 68.735000 ;
        RECT 13.245000 68.945000 13.445000 69.145000 ;
        RECT 13.245000 69.355000 13.445000 69.555000 ;
        RECT 13.245000 69.765000 13.445000 69.965000 ;
        RECT 13.245000 70.175000 13.445000 70.375000 ;
        RECT 13.245000 70.585000 13.445000 70.785000 ;
        RECT 13.245000 70.995000 13.445000 71.195000 ;
        RECT 13.245000 71.405000 13.445000 71.605000 ;
        RECT 13.245000 71.815000 13.445000 72.015000 ;
        RECT 13.245000 72.225000 13.445000 72.425000 ;
        RECT 13.245000 72.635000 13.445000 72.835000 ;
        RECT 13.245000 73.045000 13.445000 73.245000 ;
        RECT 13.245000 73.450000 13.445000 73.650000 ;
        RECT 13.245000 73.855000 13.445000 74.055000 ;
        RECT 13.245000 74.260000 13.445000 74.460000 ;
        RECT 13.245000 74.665000 13.445000 74.865000 ;
        RECT 13.245000 75.070000 13.445000 75.270000 ;
        RECT 13.245000 75.475000 13.445000 75.675000 ;
        RECT 13.245000 75.880000 13.445000 76.080000 ;
        RECT 13.245000 76.285000 13.445000 76.485000 ;
        RECT 13.245000 76.690000 13.445000 76.890000 ;
        RECT 13.245000 77.095000 13.445000 77.295000 ;
        RECT 13.245000 77.500000 13.445000 77.700000 ;
        RECT 13.245000 77.905000 13.445000 78.105000 ;
        RECT 13.245000 78.310000 13.445000 78.510000 ;
        RECT 13.245000 78.715000 13.445000 78.915000 ;
        RECT 13.245000 79.120000 13.445000 79.320000 ;
        RECT 13.245000 79.525000 13.445000 79.725000 ;
        RECT 13.245000 79.930000 13.445000 80.130000 ;
        RECT 13.245000 80.335000 13.445000 80.535000 ;
        RECT 13.245000 80.740000 13.445000 80.940000 ;
        RECT 13.245000 81.145000 13.445000 81.345000 ;
        RECT 13.245000 81.550000 13.445000 81.750000 ;
        RECT 13.245000 81.955000 13.445000 82.155000 ;
        RECT 13.245000 82.360000 13.445000 82.560000 ;
        RECT 13.435000 82.855000 13.635000 83.055000 ;
        RECT 13.435000 83.265000 13.635000 83.465000 ;
        RECT 13.435000 83.675000 13.635000 83.875000 ;
        RECT 13.435000 84.085000 13.635000 84.285000 ;
        RECT 13.435000 84.495000 13.635000 84.695000 ;
        RECT 13.435000 84.905000 13.635000 85.105000 ;
        RECT 13.435000 85.315000 13.635000 85.515000 ;
        RECT 13.435000 85.725000 13.635000 85.925000 ;
        RECT 13.435000 86.135000 13.635000 86.335000 ;
        RECT 13.435000 86.545000 13.635000 86.745000 ;
        RECT 13.435000 86.955000 13.635000 87.155000 ;
        RECT 13.435000 87.365000 13.635000 87.565000 ;
        RECT 13.435000 87.775000 13.635000 87.975000 ;
        RECT 13.435000 88.185000 13.635000 88.385000 ;
        RECT 13.435000 88.595000 13.635000 88.795000 ;
        RECT 13.435000 89.005000 13.635000 89.205000 ;
        RECT 13.435000 89.415000 13.635000 89.615000 ;
        RECT 13.435000 89.825000 13.635000 90.025000 ;
        RECT 13.435000 90.235000 13.635000 90.435000 ;
        RECT 13.435000 90.645000 13.635000 90.845000 ;
        RECT 13.435000 91.055000 13.635000 91.255000 ;
        RECT 13.435000 91.465000 13.635000 91.665000 ;
        RECT 13.435000 91.875000 13.635000 92.075000 ;
        RECT 13.435000 92.285000 13.635000 92.485000 ;
        RECT 13.435000 92.695000 13.635000 92.895000 ;
        RECT 13.645000 68.125000 13.845000 68.325000 ;
        RECT 13.645000 68.535000 13.845000 68.735000 ;
        RECT 13.645000 68.945000 13.845000 69.145000 ;
        RECT 13.645000 69.355000 13.845000 69.555000 ;
        RECT 13.645000 69.765000 13.845000 69.965000 ;
        RECT 13.645000 70.175000 13.845000 70.375000 ;
        RECT 13.645000 70.585000 13.845000 70.785000 ;
        RECT 13.645000 70.995000 13.845000 71.195000 ;
        RECT 13.645000 71.405000 13.845000 71.605000 ;
        RECT 13.645000 71.815000 13.845000 72.015000 ;
        RECT 13.645000 72.225000 13.845000 72.425000 ;
        RECT 13.645000 72.635000 13.845000 72.835000 ;
        RECT 13.645000 73.045000 13.845000 73.245000 ;
        RECT 13.645000 73.450000 13.845000 73.650000 ;
        RECT 13.645000 73.855000 13.845000 74.055000 ;
        RECT 13.645000 74.260000 13.845000 74.460000 ;
        RECT 13.645000 74.665000 13.845000 74.865000 ;
        RECT 13.645000 75.070000 13.845000 75.270000 ;
        RECT 13.645000 75.475000 13.845000 75.675000 ;
        RECT 13.645000 75.880000 13.845000 76.080000 ;
        RECT 13.645000 76.285000 13.845000 76.485000 ;
        RECT 13.645000 76.690000 13.845000 76.890000 ;
        RECT 13.645000 77.095000 13.845000 77.295000 ;
        RECT 13.645000 77.500000 13.845000 77.700000 ;
        RECT 13.645000 77.905000 13.845000 78.105000 ;
        RECT 13.645000 78.310000 13.845000 78.510000 ;
        RECT 13.645000 78.715000 13.845000 78.915000 ;
        RECT 13.645000 79.120000 13.845000 79.320000 ;
        RECT 13.645000 79.525000 13.845000 79.725000 ;
        RECT 13.645000 79.930000 13.845000 80.130000 ;
        RECT 13.645000 80.335000 13.845000 80.535000 ;
        RECT 13.645000 80.740000 13.845000 80.940000 ;
        RECT 13.645000 81.145000 13.845000 81.345000 ;
        RECT 13.645000 81.550000 13.845000 81.750000 ;
        RECT 13.645000 81.955000 13.845000 82.155000 ;
        RECT 13.645000 82.360000 13.845000 82.560000 ;
        RECT 13.650000 17.860000 13.850000 18.060000 ;
        RECT 13.650000 18.290000 13.850000 18.490000 ;
        RECT 13.650000 18.720000 13.850000 18.920000 ;
        RECT 13.650000 19.150000 13.850000 19.350000 ;
        RECT 13.650000 19.580000 13.850000 19.780000 ;
        RECT 13.650000 20.010000 13.850000 20.210000 ;
        RECT 13.650000 20.440000 13.850000 20.640000 ;
        RECT 13.650000 20.870000 13.850000 21.070000 ;
        RECT 13.650000 21.300000 13.850000 21.500000 ;
        RECT 13.650000 21.730000 13.850000 21.930000 ;
        RECT 13.650000 22.160000 13.850000 22.360000 ;
        RECT 13.840000 82.855000 14.040000 83.055000 ;
        RECT 13.840000 83.265000 14.040000 83.465000 ;
        RECT 13.840000 83.675000 14.040000 83.875000 ;
        RECT 13.840000 84.085000 14.040000 84.285000 ;
        RECT 13.840000 84.495000 14.040000 84.695000 ;
        RECT 13.840000 84.905000 14.040000 85.105000 ;
        RECT 13.840000 85.315000 14.040000 85.515000 ;
        RECT 13.840000 85.725000 14.040000 85.925000 ;
        RECT 13.840000 86.135000 14.040000 86.335000 ;
        RECT 13.840000 86.545000 14.040000 86.745000 ;
        RECT 13.840000 86.955000 14.040000 87.155000 ;
        RECT 13.840000 87.365000 14.040000 87.565000 ;
        RECT 13.840000 87.775000 14.040000 87.975000 ;
        RECT 13.840000 88.185000 14.040000 88.385000 ;
        RECT 13.840000 88.595000 14.040000 88.795000 ;
        RECT 13.840000 89.005000 14.040000 89.205000 ;
        RECT 13.840000 89.415000 14.040000 89.615000 ;
        RECT 13.840000 89.825000 14.040000 90.025000 ;
        RECT 13.840000 90.235000 14.040000 90.435000 ;
        RECT 13.840000 90.645000 14.040000 90.845000 ;
        RECT 13.840000 91.055000 14.040000 91.255000 ;
        RECT 13.840000 91.465000 14.040000 91.665000 ;
        RECT 13.840000 91.875000 14.040000 92.075000 ;
        RECT 13.840000 92.285000 14.040000 92.485000 ;
        RECT 13.840000 92.695000 14.040000 92.895000 ;
        RECT 14.045000 68.125000 14.245000 68.325000 ;
        RECT 14.045000 68.535000 14.245000 68.735000 ;
        RECT 14.045000 68.945000 14.245000 69.145000 ;
        RECT 14.045000 69.355000 14.245000 69.555000 ;
        RECT 14.045000 69.765000 14.245000 69.965000 ;
        RECT 14.045000 70.175000 14.245000 70.375000 ;
        RECT 14.045000 70.585000 14.245000 70.785000 ;
        RECT 14.045000 70.995000 14.245000 71.195000 ;
        RECT 14.045000 71.405000 14.245000 71.605000 ;
        RECT 14.045000 71.815000 14.245000 72.015000 ;
        RECT 14.045000 72.225000 14.245000 72.425000 ;
        RECT 14.045000 72.635000 14.245000 72.835000 ;
        RECT 14.045000 73.045000 14.245000 73.245000 ;
        RECT 14.045000 73.450000 14.245000 73.650000 ;
        RECT 14.045000 73.855000 14.245000 74.055000 ;
        RECT 14.045000 74.260000 14.245000 74.460000 ;
        RECT 14.045000 74.665000 14.245000 74.865000 ;
        RECT 14.045000 75.070000 14.245000 75.270000 ;
        RECT 14.045000 75.475000 14.245000 75.675000 ;
        RECT 14.045000 75.880000 14.245000 76.080000 ;
        RECT 14.045000 76.285000 14.245000 76.485000 ;
        RECT 14.045000 76.690000 14.245000 76.890000 ;
        RECT 14.045000 77.095000 14.245000 77.295000 ;
        RECT 14.045000 77.500000 14.245000 77.700000 ;
        RECT 14.045000 77.905000 14.245000 78.105000 ;
        RECT 14.045000 78.310000 14.245000 78.510000 ;
        RECT 14.045000 78.715000 14.245000 78.915000 ;
        RECT 14.045000 79.120000 14.245000 79.320000 ;
        RECT 14.045000 79.525000 14.245000 79.725000 ;
        RECT 14.045000 79.930000 14.245000 80.130000 ;
        RECT 14.045000 80.335000 14.245000 80.535000 ;
        RECT 14.045000 80.740000 14.245000 80.940000 ;
        RECT 14.045000 81.145000 14.245000 81.345000 ;
        RECT 14.045000 81.550000 14.245000 81.750000 ;
        RECT 14.045000 81.955000 14.245000 82.155000 ;
        RECT 14.045000 82.360000 14.245000 82.560000 ;
        RECT 14.055000 17.860000 14.255000 18.060000 ;
        RECT 14.055000 18.290000 14.255000 18.490000 ;
        RECT 14.055000 18.720000 14.255000 18.920000 ;
        RECT 14.055000 19.150000 14.255000 19.350000 ;
        RECT 14.055000 19.580000 14.255000 19.780000 ;
        RECT 14.055000 20.010000 14.255000 20.210000 ;
        RECT 14.055000 20.440000 14.255000 20.640000 ;
        RECT 14.055000 20.870000 14.255000 21.070000 ;
        RECT 14.055000 21.300000 14.255000 21.500000 ;
        RECT 14.055000 21.730000 14.255000 21.930000 ;
        RECT 14.055000 22.160000 14.255000 22.360000 ;
        RECT 14.320000 91.015000 14.520000 91.215000 ;
        RECT 14.320000 91.445000 14.520000 91.645000 ;
        RECT 14.340000 88.410000 14.540000 88.610000 ;
        RECT 14.340000 88.835000 14.540000 89.035000 ;
        RECT 14.340000 89.265000 14.540000 89.465000 ;
        RECT 14.340000 89.695000 14.540000 89.895000 ;
        RECT 14.340000 90.125000 14.540000 90.325000 ;
        RECT 14.340000 90.555000 14.540000 90.755000 ;
        RECT 14.445000 68.125000 14.645000 68.325000 ;
        RECT 14.445000 68.535000 14.645000 68.735000 ;
        RECT 14.445000 68.945000 14.645000 69.145000 ;
        RECT 14.445000 69.355000 14.645000 69.555000 ;
        RECT 14.445000 69.765000 14.645000 69.965000 ;
        RECT 14.445000 70.175000 14.645000 70.375000 ;
        RECT 14.445000 70.585000 14.645000 70.785000 ;
        RECT 14.445000 70.995000 14.645000 71.195000 ;
        RECT 14.445000 71.405000 14.645000 71.605000 ;
        RECT 14.445000 71.815000 14.645000 72.015000 ;
        RECT 14.445000 72.225000 14.645000 72.425000 ;
        RECT 14.445000 72.635000 14.645000 72.835000 ;
        RECT 14.445000 73.045000 14.645000 73.245000 ;
        RECT 14.445000 73.450000 14.645000 73.650000 ;
        RECT 14.445000 73.855000 14.645000 74.055000 ;
        RECT 14.445000 74.260000 14.645000 74.460000 ;
        RECT 14.445000 74.665000 14.645000 74.865000 ;
        RECT 14.445000 75.070000 14.645000 75.270000 ;
        RECT 14.445000 75.475000 14.645000 75.675000 ;
        RECT 14.445000 75.880000 14.645000 76.080000 ;
        RECT 14.445000 76.285000 14.645000 76.485000 ;
        RECT 14.445000 76.690000 14.645000 76.890000 ;
        RECT 14.445000 77.095000 14.645000 77.295000 ;
        RECT 14.445000 77.500000 14.645000 77.700000 ;
        RECT 14.445000 77.905000 14.645000 78.105000 ;
        RECT 14.445000 78.310000 14.645000 78.510000 ;
        RECT 14.445000 78.715000 14.645000 78.915000 ;
        RECT 14.445000 79.120000 14.645000 79.320000 ;
        RECT 14.445000 79.525000 14.645000 79.725000 ;
        RECT 14.445000 79.930000 14.645000 80.130000 ;
        RECT 14.445000 80.335000 14.645000 80.535000 ;
        RECT 14.445000 80.740000 14.645000 80.940000 ;
        RECT 14.445000 81.145000 14.645000 81.345000 ;
        RECT 14.445000 81.550000 14.645000 81.750000 ;
        RECT 14.445000 81.955000 14.645000 82.155000 ;
        RECT 14.445000 82.360000 14.645000 82.560000 ;
        RECT 14.460000 17.860000 14.660000 18.060000 ;
        RECT 14.460000 18.290000 14.660000 18.490000 ;
        RECT 14.460000 18.720000 14.660000 18.920000 ;
        RECT 14.460000 19.150000 14.660000 19.350000 ;
        RECT 14.460000 19.580000 14.660000 19.780000 ;
        RECT 14.460000 20.010000 14.660000 20.210000 ;
        RECT 14.460000 20.440000 14.660000 20.640000 ;
        RECT 14.460000 20.870000 14.660000 21.070000 ;
        RECT 14.460000 21.300000 14.660000 21.500000 ;
        RECT 14.460000 21.730000 14.660000 21.930000 ;
        RECT 14.460000 22.160000 14.660000 22.360000 ;
        RECT 14.465000 83.055000 14.665000 83.255000 ;
        RECT 14.465000 83.455000 14.665000 83.655000 ;
        RECT 14.465000 83.855000 14.665000 84.055000 ;
        RECT 14.465000 84.255000 14.665000 84.455000 ;
        RECT 14.465000 84.655000 14.665000 84.855000 ;
        RECT 14.465000 85.055000 14.665000 85.255000 ;
        RECT 14.465000 85.455000 14.665000 85.655000 ;
        RECT 14.465000 85.855000 14.665000 86.055000 ;
        RECT 14.465000 86.255000 14.665000 86.455000 ;
        RECT 14.465000 86.660000 14.665000 86.860000 ;
        RECT 14.465000 87.065000 14.665000 87.265000 ;
        RECT 14.465000 87.470000 14.665000 87.670000 ;
        RECT 14.465000 87.875000 14.665000 88.075000 ;
        RECT 14.750000 88.410000 14.950000 88.610000 ;
        RECT 14.750000 88.835000 14.950000 89.035000 ;
        RECT 14.750000 89.265000 14.950000 89.465000 ;
        RECT 14.750000 89.695000 14.950000 89.895000 ;
        RECT 14.750000 90.125000 14.950000 90.325000 ;
        RECT 14.750000 90.555000 14.950000 90.755000 ;
        RECT 14.845000 68.125000 15.045000 68.325000 ;
        RECT 14.845000 68.535000 15.045000 68.735000 ;
        RECT 14.845000 68.945000 15.045000 69.145000 ;
        RECT 14.845000 69.355000 15.045000 69.555000 ;
        RECT 14.845000 69.765000 15.045000 69.965000 ;
        RECT 14.845000 70.175000 15.045000 70.375000 ;
        RECT 14.845000 70.585000 15.045000 70.785000 ;
        RECT 14.845000 70.995000 15.045000 71.195000 ;
        RECT 14.845000 71.405000 15.045000 71.605000 ;
        RECT 14.845000 71.815000 15.045000 72.015000 ;
        RECT 14.845000 72.225000 15.045000 72.425000 ;
        RECT 14.845000 72.635000 15.045000 72.835000 ;
        RECT 14.845000 73.045000 15.045000 73.245000 ;
        RECT 14.845000 73.450000 15.045000 73.650000 ;
        RECT 14.845000 73.855000 15.045000 74.055000 ;
        RECT 14.845000 74.260000 15.045000 74.460000 ;
        RECT 14.845000 74.665000 15.045000 74.865000 ;
        RECT 14.845000 75.070000 15.045000 75.270000 ;
        RECT 14.845000 75.475000 15.045000 75.675000 ;
        RECT 14.845000 75.880000 15.045000 76.080000 ;
        RECT 14.845000 76.285000 15.045000 76.485000 ;
        RECT 14.845000 76.690000 15.045000 76.890000 ;
        RECT 14.845000 77.095000 15.045000 77.295000 ;
        RECT 14.845000 77.500000 15.045000 77.700000 ;
        RECT 14.845000 77.905000 15.045000 78.105000 ;
        RECT 14.845000 78.310000 15.045000 78.510000 ;
        RECT 14.845000 78.715000 15.045000 78.915000 ;
        RECT 14.845000 79.120000 15.045000 79.320000 ;
        RECT 14.845000 79.525000 15.045000 79.725000 ;
        RECT 14.845000 79.930000 15.045000 80.130000 ;
        RECT 14.845000 80.335000 15.045000 80.535000 ;
        RECT 14.845000 80.740000 15.045000 80.940000 ;
        RECT 14.845000 81.145000 15.045000 81.345000 ;
        RECT 14.845000 81.550000 15.045000 81.750000 ;
        RECT 14.845000 81.955000 15.045000 82.155000 ;
        RECT 14.845000 82.360000 15.045000 82.560000 ;
        RECT 14.865000 17.860000 15.065000 18.060000 ;
        RECT 14.865000 18.290000 15.065000 18.490000 ;
        RECT 14.865000 18.720000 15.065000 18.920000 ;
        RECT 14.865000 19.150000 15.065000 19.350000 ;
        RECT 14.865000 19.580000 15.065000 19.780000 ;
        RECT 14.865000 20.010000 15.065000 20.210000 ;
        RECT 14.865000 20.440000 15.065000 20.640000 ;
        RECT 14.865000 20.870000 15.065000 21.070000 ;
        RECT 14.865000 21.300000 15.065000 21.500000 ;
        RECT 14.865000 21.730000 15.065000 21.930000 ;
        RECT 14.865000 22.160000 15.065000 22.360000 ;
        RECT 14.875000 83.055000 15.075000 83.255000 ;
        RECT 14.875000 83.455000 15.075000 83.655000 ;
        RECT 14.875000 83.855000 15.075000 84.055000 ;
        RECT 14.875000 84.255000 15.075000 84.455000 ;
        RECT 14.875000 84.655000 15.075000 84.855000 ;
        RECT 14.875000 85.055000 15.075000 85.255000 ;
        RECT 14.875000 85.455000 15.075000 85.655000 ;
        RECT 14.875000 85.855000 15.075000 86.055000 ;
        RECT 14.875000 86.255000 15.075000 86.455000 ;
        RECT 14.875000 86.660000 15.075000 86.860000 ;
        RECT 14.875000 87.065000 15.075000 87.265000 ;
        RECT 14.875000 87.470000 15.075000 87.670000 ;
        RECT 14.875000 87.875000 15.075000 88.075000 ;
        RECT 15.100000 91.015000 15.300000 91.215000 ;
        RECT 15.100000 91.445000 15.300000 91.645000 ;
        RECT 15.160000 88.410000 15.360000 88.610000 ;
        RECT 15.160000 88.835000 15.360000 89.035000 ;
        RECT 15.160000 89.265000 15.360000 89.465000 ;
        RECT 15.160000 89.695000 15.360000 89.895000 ;
        RECT 15.160000 90.125000 15.360000 90.325000 ;
        RECT 15.160000 90.555000 15.360000 90.755000 ;
        RECT 15.245000 68.125000 15.445000 68.325000 ;
        RECT 15.245000 68.535000 15.445000 68.735000 ;
        RECT 15.245000 68.945000 15.445000 69.145000 ;
        RECT 15.245000 69.355000 15.445000 69.555000 ;
        RECT 15.245000 69.765000 15.445000 69.965000 ;
        RECT 15.245000 70.175000 15.445000 70.375000 ;
        RECT 15.245000 70.585000 15.445000 70.785000 ;
        RECT 15.245000 70.995000 15.445000 71.195000 ;
        RECT 15.245000 71.405000 15.445000 71.605000 ;
        RECT 15.245000 71.815000 15.445000 72.015000 ;
        RECT 15.245000 72.225000 15.445000 72.425000 ;
        RECT 15.245000 72.635000 15.445000 72.835000 ;
        RECT 15.245000 73.045000 15.445000 73.245000 ;
        RECT 15.245000 73.450000 15.445000 73.650000 ;
        RECT 15.245000 73.855000 15.445000 74.055000 ;
        RECT 15.245000 74.260000 15.445000 74.460000 ;
        RECT 15.245000 74.665000 15.445000 74.865000 ;
        RECT 15.245000 75.070000 15.445000 75.270000 ;
        RECT 15.245000 75.475000 15.445000 75.675000 ;
        RECT 15.245000 75.880000 15.445000 76.080000 ;
        RECT 15.245000 76.285000 15.445000 76.485000 ;
        RECT 15.245000 76.690000 15.445000 76.890000 ;
        RECT 15.245000 77.095000 15.445000 77.295000 ;
        RECT 15.245000 77.500000 15.445000 77.700000 ;
        RECT 15.245000 77.905000 15.445000 78.105000 ;
        RECT 15.245000 78.310000 15.445000 78.510000 ;
        RECT 15.245000 78.715000 15.445000 78.915000 ;
        RECT 15.245000 79.120000 15.445000 79.320000 ;
        RECT 15.245000 79.525000 15.445000 79.725000 ;
        RECT 15.245000 79.930000 15.445000 80.130000 ;
        RECT 15.245000 80.335000 15.445000 80.535000 ;
        RECT 15.245000 80.740000 15.445000 80.940000 ;
        RECT 15.245000 81.145000 15.445000 81.345000 ;
        RECT 15.245000 81.550000 15.445000 81.750000 ;
        RECT 15.245000 81.955000 15.445000 82.155000 ;
        RECT 15.245000 82.360000 15.445000 82.560000 ;
        RECT 15.270000 17.860000 15.470000 18.060000 ;
        RECT 15.270000 18.290000 15.470000 18.490000 ;
        RECT 15.270000 18.720000 15.470000 18.920000 ;
        RECT 15.270000 19.150000 15.470000 19.350000 ;
        RECT 15.270000 19.580000 15.470000 19.780000 ;
        RECT 15.270000 20.010000 15.470000 20.210000 ;
        RECT 15.270000 20.440000 15.470000 20.640000 ;
        RECT 15.270000 20.870000 15.470000 21.070000 ;
        RECT 15.270000 21.300000 15.470000 21.500000 ;
        RECT 15.270000 21.730000 15.470000 21.930000 ;
        RECT 15.270000 22.160000 15.470000 22.360000 ;
        RECT 15.285000 83.055000 15.485000 83.255000 ;
        RECT 15.285000 83.455000 15.485000 83.655000 ;
        RECT 15.285000 83.855000 15.485000 84.055000 ;
        RECT 15.285000 84.255000 15.485000 84.455000 ;
        RECT 15.285000 84.655000 15.485000 84.855000 ;
        RECT 15.285000 85.055000 15.485000 85.255000 ;
        RECT 15.285000 85.455000 15.485000 85.655000 ;
        RECT 15.285000 85.855000 15.485000 86.055000 ;
        RECT 15.285000 86.255000 15.485000 86.455000 ;
        RECT 15.285000 86.660000 15.485000 86.860000 ;
        RECT 15.285000 87.065000 15.485000 87.265000 ;
        RECT 15.285000 87.470000 15.485000 87.670000 ;
        RECT 15.285000 87.875000 15.485000 88.075000 ;
        RECT 15.570000 88.410000 15.770000 88.610000 ;
        RECT 15.570000 88.835000 15.770000 89.035000 ;
        RECT 15.570000 89.265000 15.770000 89.465000 ;
        RECT 15.570000 89.695000 15.770000 89.895000 ;
        RECT 15.570000 90.125000 15.770000 90.325000 ;
        RECT 15.570000 90.555000 15.770000 90.755000 ;
        RECT 15.645000 68.125000 15.845000 68.325000 ;
        RECT 15.645000 68.535000 15.845000 68.735000 ;
        RECT 15.645000 68.945000 15.845000 69.145000 ;
        RECT 15.645000 69.355000 15.845000 69.555000 ;
        RECT 15.645000 69.765000 15.845000 69.965000 ;
        RECT 15.645000 70.175000 15.845000 70.375000 ;
        RECT 15.645000 70.585000 15.845000 70.785000 ;
        RECT 15.645000 70.995000 15.845000 71.195000 ;
        RECT 15.645000 71.405000 15.845000 71.605000 ;
        RECT 15.645000 71.815000 15.845000 72.015000 ;
        RECT 15.645000 72.225000 15.845000 72.425000 ;
        RECT 15.645000 72.635000 15.845000 72.835000 ;
        RECT 15.645000 73.045000 15.845000 73.245000 ;
        RECT 15.645000 73.450000 15.845000 73.650000 ;
        RECT 15.645000 73.855000 15.845000 74.055000 ;
        RECT 15.645000 74.260000 15.845000 74.460000 ;
        RECT 15.645000 74.665000 15.845000 74.865000 ;
        RECT 15.645000 75.070000 15.845000 75.270000 ;
        RECT 15.645000 75.475000 15.845000 75.675000 ;
        RECT 15.645000 75.880000 15.845000 76.080000 ;
        RECT 15.645000 76.285000 15.845000 76.485000 ;
        RECT 15.645000 76.690000 15.845000 76.890000 ;
        RECT 15.645000 77.095000 15.845000 77.295000 ;
        RECT 15.645000 77.500000 15.845000 77.700000 ;
        RECT 15.645000 77.905000 15.845000 78.105000 ;
        RECT 15.645000 78.310000 15.845000 78.510000 ;
        RECT 15.645000 78.715000 15.845000 78.915000 ;
        RECT 15.645000 79.120000 15.845000 79.320000 ;
        RECT 15.645000 79.525000 15.845000 79.725000 ;
        RECT 15.645000 79.930000 15.845000 80.130000 ;
        RECT 15.645000 80.335000 15.845000 80.535000 ;
        RECT 15.645000 80.740000 15.845000 80.940000 ;
        RECT 15.645000 81.145000 15.845000 81.345000 ;
        RECT 15.645000 81.550000 15.845000 81.750000 ;
        RECT 15.645000 81.955000 15.845000 82.155000 ;
        RECT 15.645000 82.360000 15.845000 82.560000 ;
        RECT 15.675000 17.860000 15.875000 18.060000 ;
        RECT 15.675000 18.290000 15.875000 18.490000 ;
        RECT 15.675000 18.720000 15.875000 18.920000 ;
        RECT 15.675000 19.150000 15.875000 19.350000 ;
        RECT 15.675000 19.580000 15.875000 19.780000 ;
        RECT 15.675000 20.010000 15.875000 20.210000 ;
        RECT 15.675000 20.440000 15.875000 20.640000 ;
        RECT 15.675000 20.870000 15.875000 21.070000 ;
        RECT 15.675000 21.300000 15.875000 21.500000 ;
        RECT 15.675000 21.730000 15.875000 21.930000 ;
        RECT 15.675000 22.160000 15.875000 22.360000 ;
        RECT 15.695000 83.055000 15.895000 83.255000 ;
        RECT 15.695000 83.455000 15.895000 83.655000 ;
        RECT 15.695000 83.855000 15.895000 84.055000 ;
        RECT 15.695000 84.255000 15.895000 84.455000 ;
        RECT 15.695000 84.655000 15.895000 84.855000 ;
        RECT 15.695000 85.055000 15.895000 85.255000 ;
        RECT 15.695000 85.455000 15.895000 85.655000 ;
        RECT 15.695000 85.855000 15.895000 86.055000 ;
        RECT 15.695000 86.255000 15.895000 86.455000 ;
        RECT 15.695000 86.660000 15.895000 86.860000 ;
        RECT 15.695000 87.065000 15.895000 87.265000 ;
        RECT 15.695000 87.470000 15.895000 87.670000 ;
        RECT 15.695000 87.875000 15.895000 88.075000 ;
        RECT 15.980000 88.410000 16.180000 88.610000 ;
        RECT 15.980000 88.835000 16.180000 89.035000 ;
        RECT 15.980000 89.265000 16.180000 89.465000 ;
        RECT 15.980000 89.695000 16.180000 89.895000 ;
        RECT 15.980000 90.125000 16.180000 90.325000 ;
        RECT 15.980000 90.555000 16.180000 90.755000 ;
        RECT 16.045000 68.125000 16.245000 68.325000 ;
        RECT 16.045000 68.535000 16.245000 68.735000 ;
        RECT 16.045000 68.945000 16.245000 69.145000 ;
        RECT 16.045000 69.355000 16.245000 69.555000 ;
        RECT 16.045000 69.765000 16.245000 69.965000 ;
        RECT 16.045000 70.175000 16.245000 70.375000 ;
        RECT 16.045000 70.585000 16.245000 70.785000 ;
        RECT 16.045000 70.995000 16.245000 71.195000 ;
        RECT 16.045000 71.405000 16.245000 71.605000 ;
        RECT 16.045000 71.815000 16.245000 72.015000 ;
        RECT 16.045000 72.225000 16.245000 72.425000 ;
        RECT 16.045000 72.635000 16.245000 72.835000 ;
        RECT 16.045000 73.045000 16.245000 73.245000 ;
        RECT 16.045000 73.450000 16.245000 73.650000 ;
        RECT 16.045000 73.855000 16.245000 74.055000 ;
        RECT 16.045000 74.260000 16.245000 74.460000 ;
        RECT 16.045000 74.665000 16.245000 74.865000 ;
        RECT 16.045000 75.070000 16.245000 75.270000 ;
        RECT 16.045000 75.475000 16.245000 75.675000 ;
        RECT 16.045000 75.880000 16.245000 76.080000 ;
        RECT 16.045000 76.285000 16.245000 76.485000 ;
        RECT 16.045000 76.690000 16.245000 76.890000 ;
        RECT 16.045000 77.095000 16.245000 77.295000 ;
        RECT 16.045000 77.500000 16.245000 77.700000 ;
        RECT 16.045000 77.905000 16.245000 78.105000 ;
        RECT 16.045000 78.310000 16.245000 78.510000 ;
        RECT 16.045000 78.715000 16.245000 78.915000 ;
        RECT 16.045000 79.120000 16.245000 79.320000 ;
        RECT 16.045000 79.525000 16.245000 79.725000 ;
        RECT 16.045000 79.930000 16.245000 80.130000 ;
        RECT 16.045000 80.335000 16.245000 80.535000 ;
        RECT 16.045000 80.740000 16.245000 80.940000 ;
        RECT 16.045000 81.145000 16.245000 81.345000 ;
        RECT 16.045000 81.550000 16.245000 81.750000 ;
        RECT 16.045000 81.955000 16.245000 82.155000 ;
        RECT 16.045000 82.360000 16.245000 82.560000 ;
        RECT 16.080000 17.860000 16.280000 18.060000 ;
        RECT 16.080000 18.290000 16.280000 18.490000 ;
        RECT 16.080000 18.720000 16.280000 18.920000 ;
        RECT 16.080000 19.150000 16.280000 19.350000 ;
        RECT 16.080000 19.580000 16.280000 19.780000 ;
        RECT 16.080000 20.010000 16.280000 20.210000 ;
        RECT 16.080000 20.440000 16.280000 20.640000 ;
        RECT 16.080000 20.870000 16.280000 21.070000 ;
        RECT 16.080000 21.300000 16.280000 21.500000 ;
        RECT 16.080000 21.730000 16.280000 21.930000 ;
        RECT 16.080000 22.160000 16.280000 22.360000 ;
        RECT 16.105000 83.055000 16.305000 83.255000 ;
        RECT 16.105000 83.455000 16.305000 83.655000 ;
        RECT 16.105000 83.855000 16.305000 84.055000 ;
        RECT 16.105000 84.255000 16.305000 84.455000 ;
        RECT 16.105000 84.655000 16.305000 84.855000 ;
        RECT 16.105000 85.055000 16.305000 85.255000 ;
        RECT 16.105000 85.455000 16.305000 85.655000 ;
        RECT 16.105000 85.855000 16.305000 86.055000 ;
        RECT 16.105000 86.255000 16.305000 86.455000 ;
        RECT 16.105000 86.660000 16.305000 86.860000 ;
        RECT 16.105000 87.065000 16.305000 87.265000 ;
        RECT 16.105000 87.470000 16.305000 87.670000 ;
        RECT 16.105000 87.875000 16.305000 88.075000 ;
        RECT 16.445000 68.125000 16.645000 68.325000 ;
        RECT 16.445000 68.535000 16.645000 68.735000 ;
        RECT 16.445000 68.945000 16.645000 69.145000 ;
        RECT 16.445000 69.355000 16.645000 69.555000 ;
        RECT 16.445000 69.765000 16.645000 69.965000 ;
        RECT 16.445000 70.175000 16.645000 70.375000 ;
        RECT 16.445000 70.585000 16.645000 70.785000 ;
        RECT 16.445000 70.995000 16.645000 71.195000 ;
        RECT 16.445000 71.405000 16.645000 71.605000 ;
        RECT 16.445000 71.815000 16.645000 72.015000 ;
        RECT 16.445000 72.225000 16.645000 72.425000 ;
        RECT 16.445000 72.635000 16.645000 72.835000 ;
        RECT 16.445000 73.045000 16.645000 73.245000 ;
        RECT 16.445000 73.450000 16.645000 73.650000 ;
        RECT 16.445000 73.855000 16.645000 74.055000 ;
        RECT 16.445000 74.260000 16.645000 74.460000 ;
        RECT 16.445000 74.665000 16.645000 74.865000 ;
        RECT 16.445000 75.070000 16.645000 75.270000 ;
        RECT 16.445000 75.475000 16.645000 75.675000 ;
        RECT 16.445000 75.880000 16.645000 76.080000 ;
        RECT 16.445000 76.285000 16.645000 76.485000 ;
        RECT 16.445000 76.690000 16.645000 76.890000 ;
        RECT 16.445000 77.095000 16.645000 77.295000 ;
        RECT 16.445000 77.500000 16.645000 77.700000 ;
        RECT 16.445000 77.905000 16.645000 78.105000 ;
        RECT 16.445000 78.310000 16.645000 78.510000 ;
        RECT 16.445000 78.715000 16.645000 78.915000 ;
        RECT 16.445000 79.120000 16.645000 79.320000 ;
        RECT 16.445000 79.525000 16.645000 79.725000 ;
        RECT 16.445000 79.930000 16.645000 80.130000 ;
        RECT 16.445000 80.335000 16.645000 80.535000 ;
        RECT 16.445000 80.740000 16.645000 80.940000 ;
        RECT 16.445000 81.145000 16.645000 81.345000 ;
        RECT 16.445000 81.550000 16.645000 81.750000 ;
        RECT 16.445000 81.955000 16.645000 82.155000 ;
        RECT 16.445000 82.360000 16.645000 82.560000 ;
        RECT 16.480000 88.430000 16.680000 88.630000 ;
        RECT 16.480000 88.845000 16.680000 89.045000 ;
        RECT 16.480000 89.265000 16.680000 89.465000 ;
        RECT 16.485000 17.860000 16.685000 18.060000 ;
        RECT 16.485000 18.290000 16.685000 18.490000 ;
        RECT 16.485000 18.720000 16.685000 18.920000 ;
        RECT 16.485000 19.150000 16.685000 19.350000 ;
        RECT 16.485000 19.580000 16.685000 19.780000 ;
        RECT 16.485000 20.010000 16.685000 20.210000 ;
        RECT 16.485000 20.440000 16.685000 20.640000 ;
        RECT 16.485000 20.870000 16.685000 21.070000 ;
        RECT 16.485000 21.300000 16.685000 21.500000 ;
        RECT 16.485000 21.730000 16.685000 21.930000 ;
        RECT 16.485000 22.160000 16.685000 22.360000 ;
        RECT 16.515000 83.055000 16.715000 83.255000 ;
        RECT 16.515000 83.455000 16.715000 83.655000 ;
        RECT 16.515000 83.855000 16.715000 84.055000 ;
        RECT 16.515000 84.255000 16.715000 84.455000 ;
        RECT 16.515000 84.655000 16.715000 84.855000 ;
        RECT 16.515000 85.055000 16.715000 85.255000 ;
        RECT 16.515000 85.455000 16.715000 85.655000 ;
        RECT 16.515000 85.855000 16.715000 86.055000 ;
        RECT 16.515000 86.255000 16.715000 86.455000 ;
        RECT 16.515000 86.660000 16.715000 86.860000 ;
        RECT 16.515000 87.065000 16.715000 87.265000 ;
        RECT 16.515000 87.470000 16.715000 87.670000 ;
        RECT 16.515000 87.875000 16.715000 88.075000 ;
        RECT 16.845000 68.125000 17.045000 68.325000 ;
        RECT 16.845000 68.535000 17.045000 68.735000 ;
        RECT 16.845000 68.945000 17.045000 69.145000 ;
        RECT 16.845000 69.355000 17.045000 69.555000 ;
        RECT 16.845000 69.765000 17.045000 69.965000 ;
        RECT 16.845000 70.175000 17.045000 70.375000 ;
        RECT 16.845000 70.585000 17.045000 70.785000 ;
        RECT 16.845000 70.995000 17.045000 71.195000 ;
        RECT 16.845000 71.405000 17.045000 71.605000 ;
        RECT 16.845000 71.815000 17.045000 72.015000 ;
        RECT 16.845000 72.225000 17.045000 72.425000 ;
        RECT 16.845000 72.635000 17.045000 72.835000 ;
        RECT 16.845000 73.045000 17.045000 73.245000 ;
        RECT 16.845000 73.450000 17.045000 73.650000 ;
        RECT 16.845000 73.855000 17.045000 74.055000 ;
        RECT 16.845000 74.260000 17.045000 74.460000 ;
        RECT 16.845000 74.665000 17.045000 74.865000 ;
        RECT 16.845000 75.070000 17.045000 75.270000 ;
        RECT 16.845000 75.475000 17.045000 75.675000 ;
        RECT 16.845000 75.880000 17.045000 76.080000 ;
        RECT 16.845000 76.285000 17.045000 76.485000 ;
        RECT 16.845000 76.690000 17.045000 76.890000 ;
        RECT 16.845000 77.095000 17.045000 77.295000 ;
        RECT 16.845000 77.500000 17.045000 77.700000 ;
        RECT 16.845000 77.905000 17.045000 78.105000 ;
        RECT 16.845000 78.310000 17.045000 78.510000 ;
        RECT 16.845000 78.715000 17.045000 78.915000 ;
        RECT 16.845000 79.120000 17.045000 79.320000 ;
        RECT 16.845000 79.525000 17.045000 79.725000 ;
        RECT 16.845000 79.930000 17.045000 80.130000 ;
        RECT 16.845000 80.335000 17.045000 80.535000 ;
        RECT 16.845000 80.740000 17.045000 80.940000 ;
        RECT 16.845000 81.145000 17.045000 81.345000 ;
        RECT 16.845000 81.550000 17.045000 81.750000 ;
        RECT 16.845000 81.955000 17.045000 82.155000 ;
        RECT 16.845000 82.360000 17.045000 82.560000 ;
        RECT 16.890000 17.860000 17.090000 18.060000 ;
        RECT 16.890000 18.290000 17.090000 18.490000 ;
        RECT 16.890000 18.720000 17.090000 18.920000 ;
        RECT 16.890000 19.150000 17.090000 19.350000 ;
        RECT 16.890000 19.580000 17.090000 19.780000 ;
        RECT 16.890000 20.010000 17.090000 20.210000 ;
        RECT 16.890000 20.440000 17.090000 20.640000 ;
        RECT 16.890000 20.870000 17.090000 21.070000 ;
        RECT 16.890000 21.300000 17.090000 21.500000 ;
        RECT 16.890000 21.730000 17.090000 21.930000 ;
        RECT 16.890000 22.160000 17.090000 22.360000 ;
        RECT 16.925000 83.055000 17.125000 83.255000 ;
        RECT 16.925000 83.455000 17.125000 83.655000 ;
        RECT 16.925000 83.855000 17.125000 84.055000 ;
        RECT 16.925000 84.255000 17.125000 84.455000 ;
        RECT 16.925000 84.655000 17.125000 84.855000 ;
        RECT 16.925000 85.055000 17.125000 85.255000 ;
        RECT 16.925000 85.455000 17.125000 85.655000 ;
        RECT 16.925000 85.855000 17.125000 86.055000 ;
        RECT 16.925000 86.255000 17.125000 86.455000 ;
        RECT 16.925000 86.660000 17.125000 86.860000 ;
        RECT 16.925000 87.065000 17.125000 87.265000 ;
        RECT 16.925000 87.470000 17.125000 87.670000 ;
        RECT 16.925000 87.875000 17.125000 88.075000 ;
        RECT 17.245000 68.125000 17.445000 68.325000 ;
        RECT 17.245000 68.535000 17.445000 68.735000 ;
        RECT 17.245000 68.945000 17.445000 69.145000 ;
        RECT 17.245000 69.355000 17.445000 69.555000 ;
        RECT 17.245000 69.765000 17.445000 69.965000 ;
        RECT 17.245000 70.175000 17.445000 70.375000 ;
        RECT 17.245000 70.585000 17.445000 70.785000 ;
        RECT 17.245000 70.995000 17.445000 71.195000 ;
        RECT 17.245000 71.405000 17.445000 71.605000 ;
        RECT 17.245000 71.815000 17.445000 72.015000 ;
        RECT 17.245000 72.225000 17.445000 72.425000 ;
        RECT 17.245000 72.635000 17.445000 72.835000 ;
        RECT 17.245000 73.045000 17.445000 73.245000 ;
        RECT 17.245000 73.450000 17.445000 73.650000 ;
        RECT 17.245000 73.855000 17.445000 74.055000 ;
        RECT 17.245000 74.260000 17.445000 74.460000 ;
        RECT 17.245000 74.665000 17.445000 74.865000 ;
        RECT 17.245000 75.070000 17.445000 75.270000 ;
        RECT 17.245000 75.475000 17.445000 75.675000 ;
        RECT 17.245000 75.880000 17.445000 76.080000 ;
        RECT 17.245000 76.285000 17.445000 76.485000 ;
        RECT 17.245000 76.690000 17.445000 76.890000 ;
        RECT 17.245000 77.095000 17.445000 77.295000 ;
        RECT 17.245000 77.500000 17.445000 77.700000 ;
        RECT 17.245000 77.905000 17.445000 78.105000 ;
        RECT 17.245000 78.310000 17.445000 78.510000 ;
        RECT 17.245000 78.715000 17.445000 78.915000 ;
        RECT 17.245000 79.120000 17.445000 79.320000 ;
        RECT 17.245000 79.525000 17.445000 79.725000 ;
        RECT 17.245000 79.930000 17.445000 80.130000 ;
        RECT 17.245000 80.335000 17.445000 80.535000 ;
        RECT 17.245000 80.740000 17.445000 80.940000 ;
        RECT 17.245000 81.145000 17.445000 81.345000 ;
        RECT 17.245000 81.550000 17.445000 81.750000 ;
        RECT 17.245000 81.955000 17.445000 82.155000 ;
        RECT 17.245000 82.360000 17.445000 82.560000 ;
        RECT 17.260000 88.430000 17.460000 88.630000 ;
        RECT 17.260000 88.845000 17.460000 89.045000 ;
        RECT 17.260000 89.265000 17.460000 89.465000 ;
        RECT 17.295000 17.860000 17.495000 18.060000 ;
        RECT 17.295000 18.290000 17.495000 18.490000 ;
        RECT 17.295000 18.720000 17.495000 18.920000 ;
        RECT 17.295000 19.150000 17.495000 19.350000 ;
        RECT 17.295000 19.580000 17.495000 19.780000 ;
        RECT 17.295000 20.010000 17.495000 20.210000 ;
        RECT 17.295000 20.440000 17.495000 20.640000 ;
        RECT 17.295000 20.870000 17.495000 21.070000 ;
        RECT 17.295000 21.300000 17.495000 21.500000 ;
        RECT 17.295000 21.730000 17.495000 21.930000 ;
        RECT 17.295000 22.160000 17.495000 22.360000 ;
        RECT 17.335000 83.055000 17.535000 83.255000 ;
        RECT 17.335000 83.455000 17.535000 83.655000 ;
        RECT 17.335000 83.855000 17.535000 84.055000 ;
        RECT 17.335000 84.255000 17.535000 84.455000 ;
        RECT 17.335000 84.655000 17.535000 84.855000 ;
        RECT 17.335000 85.055000 17.535000 85.255000 ;
        RECT 17.335000 85.455000 17.535000 85.655000 ;
        RECT 17.335000 85.855000 17.535000 86.055000 ;
        RECT 17.335000 86.255000 17.535000 86.455000 ;
        RECT 17.335000 86.660000 17.535000 86.860000 ;
        RECT 17.335000 87.065000 17.535000 87.265000 ;
        RECT 17.335000 87.470000 17.535000 87.670000 ;
        RECT 17.335000 87.875000 17.535000 88.075000 ;
        RECT 17.645000 68.125000 17.845000 68.325000 ;
        RECT 17.645000 68.535000 17.845000 68.735000 ;
        RECT 17.645000 68.945000 17.845000 69.145000 ;
        RECT 17.645000 69.355000 17.845000 69.555000 ;
        RECT 17.645000 69.765000 17.845000 69.965000 ;
        RECT 17.645000 70.175000 17.845000 70.375000 ;
        RECT 17.645000 70.585000 17.845000 70.785000 ;
        RECT 17.645000 70.995000 17.845000 71.195000 ;
        RECT 17.645000 71.405000 17.845000 71.605000 ;
        RECT 17.645000 71.815000 17.845000 72.015000 ;
        RECT 17.645000 72.225000 17.845000 72.425000 ;
        RECT 17.645000 72.635000 17.845000 72.835000 ;
        RECT 17.645000 73.045000 17.845000 73.245000 ;
        RECT 17.645000 73.450000 17.845000 73.650000 ;
        RECT 17.645000 73.855000 17.845000 74.055000 ;
        RECT 17.645000 74.260000 17.845000 74.460000 ;
        RECT 17.645000 74.665000 17.845000 74.865000 ;
        RECT 17.645000 75.070000 17.845000 75.270000 ;
        RECT 17.645000 75.475000 17.845000 75.675000 ;
        RECT 17.645000 75.880000 17.845000 76.080000 ;
        RECT 17.645000 76.285000 17.845000 76.485000 ;
        RECT 17.645000 76.690000 17.845000 76.890000 ;
        RECT 17.645000 77.095000 17.845000 77.295000 ;
        RECT 17.645000 77.500000 17.845000 77.700000 ;
        RECT 17.645000 77.905000 17.845000 78.105000 ;
        RECT 17.645000 78.310000 17.845000 78.510000 ;
        RECT 17.645000 78.715000 17.845000 78.915000 ;
        RECT 17.645000 79.120000 17.845000 79.320000 ;
        RECT 17.645000 79.525000 17.845000 79.725000 ;
        RECT 17.645000 79.930000 17.845000 80.130000 ;
        RECT 17.645000 80.335000 17.845000 80.535000 ;
        RECT 17.645000 80.740000 17.845000 80.940000 ;
        RECT 17.645000 81.145000 17.845000 81.345000 ;
        RECT 17.645000 81.550000 17.845000 81.750000 ;
        RECT 17.645000 81.955000 17.845000 82.155000 ;
        RECT 17.645000 82.360000 17.845000 82.560000 ;
        RECT 17.700000 17.860000 17.900000 18.060000 ;
        RECT 17.700000 18.290000 17.900000 18.490000 ;
        RECT 17.700000 18.720000 17.900000 18.920000 ;
        RECT 17.700000 19.150000 17.900000 19.350000 ;
        RECT 17.700000 19.580000 17.900000 19.780000 ;
        RECT 17.700000 20.010000 17.900000 20.210000 ;
        RECT 17.700000 20.440000 17.900000 20.640000 ;
        RECT 17.700000 20.870000 17.900000 21.070000 ;
        RECT 17.700000 21.300000 17.900000 21.500000 ;
        RECT 17.700000 21.730000 17.900000 21.930000 ;
        RECT 17.700000 22.160000 17.900000 22.360000 ;
        RECT 17.745000 83.055000 17.945000 83.255000 ;
        RECT 17.745000 83.455000 17.945000 83.655000 ;
        RECT 17.745000 83.855000 17.945000 84.055000 ;
        RECT 17.745000 84.255000 17.945000 84.455000 ;
        RECT 17.745000 84.655000 17.945000 84.855000 ;
        RECT 17.745000 85.055000 17.945000 85.255000 ;
        RECT 17.745000 85.455000 17.945000 85.655000 ;
        RECT 17.745000 85.855000 17.945000 86.055000 ;
        RECT 17.745000 86.255000 17.945000 86.455000 ;
        RECT 17.745000 86.660000 17.945000 86.860000 ;
        RECT 17.745000 87.065000 17.945000 87.265000 ;
        RECT 17.745000 87.470000 17.945000 87.670000 ;
        RECT 17.745000 87.875000 17.945000 88.075000 ;
        RECT 18.045000 68.125000 18.245000 68.325000 ;
        RECT 18.045000 68.535000 18.245000 68.735000 ;
        RECT 18.045000 68.945000 18.245000 69.145000 ;
        RECT 18.045000 69.355000 18.245000 69.555000 ;
        RECT 18.045000 69.765000 18.245000 69.965000 ;
        RECT 18.045000 70.175000 18.245000 70.375000 ;
        RECT 18.045000 70.585000 18.245000 70.785000 ;
        RECT 18.045000 70.995000 18.245000 71.195000 ;
        RECT 18.045000 71.405000 18.245000 71.605000 ;
        RECT 18.045000 71.815000 18.245000 72.015000 ;
        RECT 18.045000 72.225000 18.245000 72.425000 ;
        RECT 18.045000 72.635000 18.245000 72.835000 ;
        RECT 18.045000 73.045000 18.245000 73.245000 ;
        RECT 18.045000 73.450000 18.245000 73.650000 ;
        RECT 18.045000 73.855000 18.245000 74.055000 ;
        RECT 18.045000 74.260000 18.245000 74.460000 ;
        RECT 18.045000 74.665000 18.245000 74.865000 ;
        RECT 18.045000 75.070000 18.245000 75.270000 ;
        RECT 18.045000 75.475000 18.245000 75.675000 ;
        RECT 18.045000 75.880000 18.245000 76.080000 ;
        RECT 18.045000 76.285000 18.245000 76.485000 ;
        RECT 18.045000 76.690000 18.245000 76.890000 ;
        RECT 18.045000 77.095000 18.245000 77.295000 ;
        RECT 18.045000 77.500000 18.245000 77.700000 ;
        RECT 18.045000 77.905000 18.245000 78.105000 ;
        RECT 18.045000 78.310000 18.245000 78.510000 ;
        RECT 18.045000 78.715000 18.245000 78.915000 ;
        RECT 18.045000 79.120000 18.245000 79.320000 ;
        RECT 18.045000 79.525000 18.245000 79.725000 ;
        RECT 18.045000 79.930000 18.245000 80.130000 ;
        RECT 18.045000 80.335000 18.245000 80.535000 ;
        RECT 18.045000 80.740000 18.245000 80.940000 ;
        RECT 18.045000 81.145000 18.245000 81.345000 ;
        RECT 18.045000 81.550000 18.245000 81.750000 ;
        RECT 18.045000 81.955000 18.245000 82.155000 ;
        RECT 18.045000 82.360000 18.245000 82.560000 ;
        RECT 18.105000 17.860000 18.305000 18.060000 ;
        RECT 18.105000 18.290000 18.305000 18.490000 ;
        RECT 18.105000 18.720000 18.305000 18.920000 ;
        RECT 18.105000 19.150000 18.305000 19.350000 ;
        RECT 18.105000 19.580000 18.305000 19.780000 ;
        RECT 18.105000 20.010000 18.305000 20.210000 ;
        RECT 18.105000 20.440000 18.305000 20.640000 ;
        RECT 18.105000 20.870000 18.305000 21.070000 ;
        RECT 18.105000 21.300000 18.305000 21.500000 ;
        RECT 18.105000 21.730000 18.305000 21.930000 ;
        RECT 18.105000 22.160000 18.305000 22.360000 ;
        RECT 18.155000 83.055000 18.355000 83.255000 ;
        RECT 18.155000 83.455000 18.355000 83.655000 ;
        RECT 18.155000 83.855000 18.355000 84.055000 ;
        RECT 18.155000 84.255000 18.355000 84.455000 ;
        RECT 18.155000 84.655000 18.355000 84.855000 ;
        RECT 18.155000 85.055000 18.355000 85.255000 ;
        RECT 18.155000 85.455000 18.355000 85.655000 ;
        RECT 18.155000 85.855000 18.355000 86.055000 ;
        RECT 18.155000 86.255000 18.355000 86.455000 ;
        RECT 18.155000 86.660000 18.355000 86.860000 ;
        RECT 18.155000 87.065000 18.355000 87.265000 ;
        RECT 18.155000 87.470000 18.355000 87.670000 ;
        RECT 18.155000 87.875000 18.355000 88.075000 ;
        RECT 18.445000 68.125000 18.645000 68.325000 ;
        RECT 18.445000 68.535000 18.645000 68.735000 ;
        RECT 18.445000 68.945000 18.645000 69.145000 ;
        RECT 18.445000 69.355000 18.645000 69.555000 ;
        RECT 18.445000 69.765000 18.645000 69.965000 ;
        RECT 18.445000 70.175000 18.645000 70.375000 ;
        RECT 18.445000 70.585000 18.645000 70.785000 ;
        RECT 18.445000 70.995000 18.645000 71.195000 ;
        RECT 18.445000 71.405000 18.645000 71.605000 ;
        RECT 18.445000 71.815000 18.645000 72.015000 ;
        RECT 18.445000 72.225000 18.645000 72.425000 ;
        RECT 18.445000 72.635000 18.645000 72.835000 ;
        RECT 18.445000 73.045000 18.645000 73.245000 ;
        RECT 18.445000 73.450000 18.645000 73.650000 ;
        RECT 18.445000 73.855000 18.645000 74.055000 ;
        RECT 18.445000 74.260000 18.645000 74.460000 ;
        RECT 18.445000 74.665000 18.645000 74.865000 ;
        RECT 18.445000 75.070000 18.645000 75.270000 ;
        RECT 18.445000 75.475000 18.645000 75.675000 ;
        RECT 18.445000 75.880000 18.645000 76.080000 ;
        RECT 18.445000 76.285000 18.645000 76.485000 ;
        RECT 18.445000 76.690000 18.645000 76.890000 ;
        RECT 18.445000 77.095000 18.645000 77.295000 ;
        RECT 18.445000 77.500000 18.645000 77.700000 ;
        RECT 18.445000 77.905000 18.645000 78.105000 ;
        RECT 18.445000 78.310000 18.645000 78.510000 ;
        RECT 18.445000 78.715000 18.645000 78.915000 ;
        RECT 18.445000 79.120000 18.645000 79.320000 ;
        RECT 18.445000 79.525000 18.645000 79.725000 ;
        RECT 18.445000 79.930000 18.645000 80.130000 ;
        RECT 18.445000 80.335000 18.645000 80.535000 ;
        RECT 18.445000 80.740000 18.645000 80.940000 ;
        RECT 18.445000 81.145000 18.645000 81.345000 ;
        RECT 18.445000 81.550000 18.645000 81.750000 ;
        RECT 18.445000 81.955000 18.645000 82.155000 ;
        RECT 18.445000 82.360000 18.645000 82.560000 ;
        RECT 18.510000 17.860000 18.710000 18.060000 ;
        RECT 18.510000 18.290000 18.710000 18.490000 ;
        RECT 18.510000 18.720000 18.710000 18.920000 ;
        RECT 18.510000 19.150000 18.710000 19.350000 ;
        RECT 18.510000 19.580000 18.710000 19.780000 ;
        RECT 18.510000 20.010000 18.710000 20.210000 ;
        RECT 18.510000 20.440000 18.710000 20.640000 ;
        RECT 18.510000 20.870000 18.710000 21.070000 ;
        RECT 18.510000 21.300000 18.710000 21.500000 ;
        RECT 18.510000 21.730000 18.710000 21.930000 ;
        RECT 18.510000 22.160000 18.710000 22.360000 ;
        RECT 18.565000 83.055000 18.765000 83.255000 ;
        RECT 18.565000 83.455000 18.765000 83.655000 ;
        RECT 18.565000 83.855000 18.765000 84.055000 ;
        RECT 18.565000 84.255000 18.765000 84.455000 ;
        RECT 18.565000 84.655000 18.765000 84.855000 ;
        RECT 18.565000 85.055000 18.765000 85.255000 ;
        RECT 18.565000 85.455000 18.765000 85.655000 ;
        RECT 18.565000 85.855000 18.765000 86.055000 ;
        RECT 18.565000 86.255000 18.765000 86.455000 ;
        RECT 18.565000 86.660000 18.765000 86.860000 ;
        RECT 18.565000 87.065000 18.765000 87.265000 ;
        RECT 18.565000 87.470000 18.765000 87.670000 ;
        RECT 18.565000 87.875000 18.765000 88.075000 ;
        RECT 18.845000 68.125000 19.045000 68.325000 ;
        RECT 18.845000 68.535000 19.045000 68.735000 ;
        RECT 18.845000 68.945000 19.045000 69.145000 ;
        RECT 18.845000 69.355000 19.045000 69.555000 ;
        RECT 18.845000 69.765000 19.045000 69.965000 ;
        RECT 18.845000 70.175000 19.045000 70.375000 ;
        RECT 18.845000 70.585000 19.045000 70.785000 ;
        RECT 18.845000 70.995000 19.045000 71.195000 ;
        RECT 18.845000 71.405000 19.045000 71.605000 ;
        RECT 18.845000 71.815000 19.045000 72.015000 ;
        RECT 18.845000 72.225000 19.045000 72.425000 ;
        RECT 18.845000 72.635000 19.045000 72.835000 ;
        RECT 18.845000 73.045000 19.045000 73.245000 ;
        RECT 18.845000 73.450000 19.045000 73.650000 ;
        RECT 18.845000 73.855000 19.045000 74.055000 ;
        RECT 18.845000 74.260000 19.045000 74.460000 ;
        RECT 18.845000 74.665000 19.045000 74.865000 ;
        RECT 18.845000 75.070000 19.045000 75.270000 ;
        RECT 18.845000 75.475000 19.045000 75.675000 ;
        RECT 18.845000 75.880000 19.045000 76.080000 ;
        RECT 18.845000 76.285000 19.045000 76.485000 ;
        RECT 18.845000 76.690000 19.045000 76.890000 ;
        RECT 18.845000 77.095000 19.045000 77.295000 ;
        RECT 18.845000 77.500000 19.045000 77.700000 ;
        RECT 18.845000 77.905000 19.045000 78.105000 ;
        RECT 18.845000 78.310000 19.045000 78.510000 ;
        RECT 18.845000 78.715000 19.045000 78.915000 ;
        RECT 18.845000 79.120000 19.045000 79.320000 ;
        RECT 18.845000 79.525000 19.045000 79.725000 ;
        RECT 18.845000 79.930000 19.045000 80.130000 ;
        RECT 18.845000 80.335000 19.045000 80.535000 ;
        RECT 18.845000 80.740000 19.045000 80.940000 ;
        RECT 18.845000 81.145000 19.045000 81.345000 ;
        RECT 18.845000 81.550000 19.045000 81.750000 ;
        RECT 18.845000 81.955000 19.045000 82.155000 ;
        RECT 18.845000 82.360000 19.045000 82.560000 ;
        RECT 18.915000 17.860000 19.115000 18.060000 ;
        RECT 18.915000 18.290000 19.115000 18.490000 ;
        RECT 18.915000 18.720000 19.115000 18.920000 ;
        RECT 18.915000 19.150000 19.115000 19.350000 ;
        RECT 18.915000 19.580000 19.115000 19.780000 ;
        RECT 18.915000 20.010000 19.115000 20.210000 ;
        RECT 18.915000 20.440000 19.115000 20.640000 ;
        RECT 18.915000 20.870000 19.115000 21.070000 ;
        RECT 18.915000 21.300000 19.115000 21.500000 ;
        RECT 18.915000 21.730000 19.115000 21.930000 ;
        RECT 18.915000 22.160000 19.115000 22.360000 ;
        RECT 19.060000 85.875000 19.260000 86.075000 ;
        RECT 19.060000 86.310000 19.260000 86.510000 ;
        RECT 19.060000 86.750000 19.260000 86.950000 ;
        RECT 19.245000 68.125000 19.445000 68.325000 ;
        RECT 19.245000 68.535000 19.445000 68.735000 ;
        RECT 19.245000 68.945000 19.445000 69.145000 ;
        RECT 19.245000 69.355000 19.445000 69.555000 ;
        RECT 19.245000 69.765000 19.445000 69.965000 ;
        RECT 19.245000 70.175000 19.445000 70.375000 ;
        RECT 19.245000 70.585000 19.445000 70.785000 ;
        RECT 19.245000 70.995000 19.445000 71.195000 ;
        RECT 19.245000 71.405000 19.445000 71.605000 ;
        RECT 19.245000 71.815000 19.445000 72.015000 ;
        RECT 19.245000 72.225000 19.445000 72.425000 ;
        RECT 19.245000 72.635000 19.445000 72.835000 ;
        RECT 19.245000 73.045000 19.445000 73.245000 ;
        RECT 19.245000 73.450000 19.445000 73.650000 ;
        RECT 19.245000 73.855000 19.445000 74.055000 ;
        RECT 19.245000 74.260000 19.445000 74.460000 ;
        RECT 19.245000 74.665000 19.445000 74.865000 ;
        RECT 19.245000 75.070000 19.445000 75.270000 ;
        RECT 19.245000 75.475000 19.445000 75.675000 ;
        RECT 19.245000 75.880000 19.445000 76.080000 ;
        RECT 19.245000 76.285000 19.445000 76.485000 ;
        RECT 19.245000 76.690000 19.445000 76.890000 ;
        RECT 19.245000 77.095000 19.445000 77.295000 ;
        RECT 19.245000 77.500000 19.445000 77.700000 ;
        RECT 19.245000 77.905000 19.445000 78.105000 ;
        RECT 19.245000 78.310000 19.445000 78.510000 ;
        RECT 19.245000 78.715000 19.445000 78.915000 ;
        RECT 19.245000 79.120000 19.445000 79.320000 ;
        RECT 19.245000 79.525000 19.445000 79.725000 ;
        RECT 19.245000 79.930000 19.445000 80.130000 ;
        RECT 19.245000 80.335000 19.445000 80.535000 ;
        RECT 19.245000 80.740000 19.445000 80.940000 ;
        RECT 19.245000 81.145000 19.445000 81.345000 ;
        RECT 19.245000 81.550000 19.445000 81.750000 ;
        RECT 19.245000 81.955000 19.445000 82.155000 ;
        RECT 19.245000 82.360000 19.445000 82.560000 ;
        RECT 19.250000 83.010000 19.450000 83.210000 ;
        RECT 19.250000 83.470000 19.450000 83.670000 ;
        RECT 19.250000 83.930000 19.450000 84.130000 ;
        RECT 19.250000 84.395000 19.450000 84.595000 ;
        RECT 19.250000 84.860000 19.450000 85.060000 ;
        RECT 19.250000 85.325000 19.450000 85.525000 ;
        RECT 19.320000 17.860000 19.520000 18.060000 ;
        RECT 19.320000 18.290000 19.520000 18.490000 ;
        RECT 19.320000 18.720000 19.520000 18.920000 ;
        RECT 19.320000 19.150000 19.520000 19.350000 ;
        RECT 19.320000 19.580000 19.520000 19.780000 ;
        RECT 19.320000 20.010000 19.520000 20.210000 ;
        RECT 19.320000 20.440000 19.520000 20.640000 ;
        RECT 19.320000 20.870000 19.520000 21.070000 ;
        RECT 19.320000 21.300000 19.520000 21.500000 ;
        RECT 19.320000 21.730000 19.520000 21.930000 ;
        RECT 19.320000 22.160000 19.520000 22.360000 ;
        RECT 19.645000 68.125000 19.845000 68.325000 ;
        RECT 19.645000 68.535000 19.845000 68.735000 ;
        RECT 19.645000 68.945000 19.845000 69.145000 ;
        RECT 19.645000 69.355000 19.845000 69.555000 ;
        RECT 19.645000 69.765000 19.845000 69.965000 ;
        RECT 19.645000 70.175000 19.845000 70.375000 ;
        RECT 19.645000 70.585000 19.845000 70.785000 ;
        RECT 19.645000 70.995000 19.845000 71.195000 ;
        RECT 19.645000 71.405000 19.845000 71.605000 ;
        RECT 19.645000 71.815000 19.845000 72.015000 ;
        RECT 19.645000 72.225000 19.845000 72.425000 ;
        RECT 19.645000 72.635000 19.845000 72.835000 ;
        RECT 19.645000 73.045000 19.845000 73.245000 ;
        RECT 19.645000 73.450000 19.845000 73.650000 ;
        RECT 19.645000 73.855000 19.845000 74.055000 ;
        RECT 19.645000 74.260000 19.845000 74.460000 ;
        RECT 19.645000 74.665000 19.845000 74.865000 ;
        RECT 19.645000 75.070000 19.845000 75.270000 ;
        RECT 19.645000 75.475000 19.845000 75.675000 ;
        RECT 19.645000 75.880000 19.845000 76.080000 ;
        RECT 19.645000 76.285000 19.845000 76.485000 ;
        RECT 19.645000 76.690000 19.845000 76.890000 ;
        RECT 19.645000 77.095000 19.845000 77.295000 ;
        RECT 19.645000 77.500000 19.845000 77.700000 ;
        RECT 19.645000 77.905000 19.845000 78.105000 ;
        RECT 19.645000 78.310000 19.845000 78.510000 ;
        RECT 19.645000 78.715000 19.845000 78.915000 ;
        RECT 19.645000 79.120000 19.845000 79.320000 ;
        RECT 19.645000 79.525000 19.845000 79.725000 ;
        RECT 19.645000 79.930000 19.845000 80.130000 ;
        RECT 19.645000 80.335000 19.845000 80.535000 ;
        RECT 19.645000 80.740000 19.845000 80.940000 ;
        RECT 19.645000 81.145000 19.845000 81.345000 ;
        RECT 19.645000 81.550000 19.845000 81.750000 ;
        RECT 19.645000 81.955000 19.845000 82.155000 ;
        RECT 19.645000 82.360000 19.845000 82.560000 ;
        RECT 19.725000 17.860000 19.925000 18.060000 ;
        RECT 19.725000 18.290000 19.925000 18.490000 ;
        RECT 19.725000 18.720000 19.925000 18.920000 ;
        RECT 19.725000 19.150000 19.925000 19.350000 ;
        RECT 19.725000 19.580000 19.925000 19.780000 ;
        RECT 19.725000 20.010000 19.925000 20.210000 ;
        RECT 19.725000 20.440000 19.925000 20.640000 ;
        RECT 19.725000 20.870000 19.925000 21.070000 ;
        RECT 19.725000 21.300000 19.925000 21.500000 ;
        RECT 19.725000 21.730000 19.925000 21.930000 ;
        RECT 19.725000 22.160000 19.925000 22.360000 ;
        RECT 19.730000 83.010000 19.930000 83.210000 ;
        RECT 19.730000 83.470000 19.930000 83.670000 ;
        RECT 19.730000 83.930000 19.930000 84.130000 ;
        RECT 19.730000 84.395000 19.930000 84.595000 ;
        RECT 19.730000 84.860000 19.930000 85.060000 ;
        RECT 19.730000 85.325000 19.930000 85.525000 ;
        RECT 19.800000 85.875000 20.000000 86.075000 ;
        RECT 19.800000 86.310000 20.000000 86.510000 ;
        RECT 19.800000 86.750000 20.000000 86.950000 ;
        RECT 20.045000 68.125000 20.245000 68.325000 ;
        RECT 20.045000 68.535000 20.245000 68.735000 ;
        RECT 20.045000 68.945000 20.245000 69.145000 ;
        RECT 20.045000 69.355000 20.245000 69.555000 ;
        RECT 20.045000 69.765000 20.245000 69.965000 ;
        RECT 20.045000 70.175000 20.245000 70.375000 ;
        RECT 20.045000 70.585000 20.245000 70.785000 ;
        RECT 20.045000 70.995000 20.245000 71.195000 ;
        RECT 20.045000 71.405000 20.245000 71.605000 ;
        RECT 20.045000 71.815000 20.245000 72.015000 ;
        RECT 20.045000 72.225000 20.245000 72.425000 ;
        RECT 20.045000 72.635000 20.245000 72.835000 ;
        RECT 20.045000 73.045000 20.245000 73.245000 ;
        RECT 20.045000 73.450000 20.245000 73.650000 ;
        RECT 20.045000 73.855000 20.245000 74.055000 ;
        RECT 20.045000 74.260000 20.245000 74.460000 ;
        RECT 20.045000 74.665000 20.245000 74.865000 ;
        RECT 20.045000 75.070000 20.245000 75.270000 ;
        RECT 20.045000 75.475000 20.245000 75.675000 ;
        RECT 20.045000 75.880000 20.245000 76.080000 ;
        RECT 20.045000 76.285000 20.245000 76.485000 ;
        RECT 20.045000 76.690000 20.245000 76.890000 ;
        RECT 20.045000 77.095000 20.245000 77.295000 ;
        RECT 20.045000 77.500000 20.245000 77.700000 ;
        RECT 20.045000 77.905000 20.245000 78.105000 ;
        RECT 20.045000 78.310000 20.245000 78.510000 ;
        RECT 20.045000 78.715000 20.245000 78.915000 ;
        RECT 20.045000 79.120000 20.245000 79.320000 ;
        RECT 20.045000 79.525000 20.245000 79.725000 ;
        RECT 20.045000 79.930000 20.245000 80.130000 ;
        RECT 20.045000 80.335000 20.245000 80.535000 ;
        RECT 20.045000 80.740000 20.245000 80.940000 ;
        RECT 20.045000 81.145000 20.245000 81.345000 ;
        RECT 20.045000 81.550000 20.245000 81.750000 ;
        RECT 20.045000 81.955000 20.245000 82.155000 ;
        RECT 20.045000 82.360000 20.245000 82.560000 ;
        RECT 20.130000 17.860000 20.330000 18.060000 ;
        RECT 20.130000 18.290000 20.330000 18.490000 ;
        RECT 20.130000 18.720000 20.330000 18.920000 ;
        RECT 20.130000 19.150000 20.330000 19.350000 ;
        RECT 20.130000 19.580000 20.330000 19.780000 ;
        RECT 20.130000 20.010000 20.330000 20.210000 ;
        RECT 20.130000 20.440000 20.330000 20.640000 ;
        RECT 20.130000 20.870000 20.330000 21.070000 ;
        RECT 20.130000 21.300000 20.330000 21.500000 ;
        RECT 20.130000 21.730000 20.330000 21.930000 ;
        RECT 20.130000 22.160000 20.330000 22.360000 ;
        RECT 20.210000 83.010000 20.410000 83.210000 ;
        RECT 20.210000 83.470000 20.410000 83.670000 ;
        RECT 20.210000 83.930000 20.410000 84.130000 ;
        RECT 20.210000 84.395000 20.410000 84.595000 ;
        RECT 20.210000 84.860000 20.410000 85.060000 ;
        RECT 20.210000 85.325000 20.410000 85.525000 ;
        RECT 20.445000 68.125000 20.645000 68.325000 ;
        RECT 20.445000 68.535000 20.645000 68.735000 ;
        RECT 20.445000 68.945000 20.645000 69.145000 ;
        RECT 20.445000 69.355000 20.645000 69.555000 ;
        RECT 20.445000 69.765000 20.645000 69.965000 ;
        RECT 20.445000 70.175000 20.645000 70.375000 ;
        RECT 20.445000 70.585000 20.645000 70.785000 ;
        RECT 20.445000 70.995000 20.645000 71.195000 ;
        RECT 20.445000 71.405000 20.645000 71.605000 ;
        RECT 20.445000 71.815000 20.645000 72.015000 ;
        RECT 20.445000 72.225000 20.645000 72.425000 ;
        RECT 20.445000 72.635000 20.645000 72.835000 ;
        RECT 20.445000 73.045000 20.645000 73.245000 ;
        RECT 20.445000 73.450000 20.645000 73.650000 ;
        RECT 20.445000 73.855000 20.645000 74.055000 ;
        RECT 20.445000 74.260000 20.645000 74.460000 ;
        RECT 20.445000 74.665000 20.645000 74.865000 ;
        RECT 20.445000 75.070000 20.645000 75.270000 ;
        RECT 20.445000 75.475000 20.645000 75.675000 ;
        RECT 20.445000 75.880000 20.645000 76.080000 ;
        RECT 20.445000 76.285000 20.645000 76.485000 ;
        RECT 20.445000 76.690000 20.645000 76.890000 ;
        RECT 20.445000 77.095000 20.645000 77.295000 ;
        RECT 20.445000 77.500000 20.645000 77.700000 ;
        RECT 20.445000 77.905000 20.645000 78.105000 ;
        RECT 20.445000 78.310000 20.645000 78.510000 ;
        RECT 20.445000 78.715000 20.645000 78.915000 ;
        RECT 20.445000 79.120000 20.645000 79.320000 ;
        RECT 20.445000 79.525000 20.645000 79.725000 ;
        RECT 20.445000 79.930000 20.645000 80.130000 ;
        RECT 20.445000 80.335000 20.645000 80.535000 ;
        RECT 20.445000 80.740000 20.645000 80.940000 ;
        RECT 20.445000 81.145000 20.645000 81.345000 ;
        RECT 20.445000 81.550000 20.645000 81.750000 ;
        RECT 20.445000 81.955000 20.645000 82.155000 ;
        RECT 20.445000 82.360000 20.645000 82.560000 ;
        RECT 20.535000 17.860000 20.735000 18.060000 ;
        RECT 20.535000 18.290000 20.735000 18.490000 ;
        RECT 20.535000 18.720000 20.735000 18.920000 ;
        RECT 20.535000 19.150000 20.735000 19.350000 ;
        RECT 20.535000 19.580000 20.735000 19.780000 ;
        RECT 20.535000 20.010000 20.735000 20.210000 ;
        RECT 20.535000 20.440000 20.735000 20.640000 ;
        RECT 20.535000 20.870000 20.735000 21.070000 ;
        RECT 20.535000 21.300000 20.735000 21.500000 ;
        RECT 20.535000 21.730000 20.735000 21.930000 ;
        RECT 20.535000 22.160000 20.735000 22.360000 ;
        RECT 20.690000 83.010000 20.890000 83.210000 ;
        RECT 20.690000 83.470000 20.890000 83.670000 ;
        RECT 20.690000 83.930000 20.890000 84.130000 ;
        RECT 20.690000 84.395000 20.890000 84.595000 ;
        RECT 20.690000 84.860000 20.890000 85.060000 ;
        RECT 20.690000 85.325000 20.890000 85.525000 ;
        RECT 20.845000 68.125000 21.045000 68.325000 ;
        RECT 20.845000 68.535000 21.045000 68.735000 ;
        RECT 20.845000 68.945000 21.045000 69.145000 ;
        RECT 20.845000 69.355000 21.045000 69.555000 ;
        RECT 20.845000 69.765000 21.045000 69.965000 ;
        RECT 20.845000 70.175000 21.045000 70.375000 ;
        RECT 20.845000 70.585000 21.045000 70.785000 ;
        RECT 20.845000 70.995000 21.045000 71.195000 ;
        RECT 20.845000 71.405000 21.045000 71.605000 ;
        RECT 20.845000 71.815000 21.045000 72.015000 ;
        RECT 20.845000 72.225000 21.045000 72.425000 ;
        RECT 20.845000 72.635000 21.045000 72.835000 ;
        RECT 20.845000 73.045000 21.045000 73.245000 ;
        RECT 20.845000 73.450000 21.045000 73.650000 ;
        RECT 20.845000 73.855000 21.045000 74.055000 ;
        RECT 20.845000 74.260000 21.045000 74.460000 ;
        RECT 20.845000 74.665000 21.045000 74.865000 ;
        RECT 20.845000 75.070000 21.045000 75.270000 ;
        RECT 20.845000 75.475000 21.045000 75.675000 ;
        RECT 20.845000 75.880000 21.045000 76.080000 ;
        RECT 20.845000 76.285000 21.045000 76.485000 ;
        RECT 20.845000 76.690000 21.045000 76.890000 ;
        RECT 20.845000 77.095000 21.045000 77.295000 ;
        RECT 20.845000 77.500000 21.045000 77.700000 ;
        RECT 20.845000 77.905000 21.045000 78.105000 ;
        RECT 20.845000 78.310000 21.045000 78.510000 ;
        RECT 20.845000 78.715000 21.045000 78.915000 ;
        RECT 20.845000 79.120000 21.045000 79.320000 ;
        RECT 20.845000 79.525000 21.045000 79.725000 ;
        RECT 20.845000 79.930000 21.045000 80.130000 ;
        RECT 20.845000 80.335000 21.045000 80.535000 ;
        RECT 20.845000 80.740000 21.045000 80.940000 ;
        RECT 20.845000 81.145000 21.045000 81.345000 ;
        RECT 20.845000 81.550000 21.045000 81.750000 ;
        RECT 20.845000 81.955000 21.045000 82.155000 ;
        RECT 20.845000 82.360000 21.045000 82.560000 ;
        RECT 20.940000 17.860000 21.140000 18.060000 ;
        RECT 20.940000 18.290000 21.140000 18.490000 ;
        RECT 20.940000 18.720000 21.140000 18.920000 ;
        RECT 20.940000 19.150000 21.140000 19.350000 ;
        RECT 20.940000 19.580000 21.140000 19.780000 ;
        RECT 20.940000 20.010000 21.140000 20.210000 ;
        RECT 20.940000 20.440000 21.140000 20.640000 ;
        RECT 20.940000 20.870000 21.140000 21.070000 ;
        RECT 20.940000 21.300000 21.140000 21.500000 ;
        RECT 20.940000 21.730000 21.140000 21.930000 ;
        RECT 20.940000 22.160000 21.140000 22.360000 ;
        RECT 21.170000 83.010000 21.370000 83.210000 ;
        RECT 21.170000 83.470000 21.370000 83.670000 ;
        RECT 21.170000 83.930000 21.370000 84.130000 ;
        RECT 21.170000 84.395000 21.370000 84.595000 ;
        RECT 21.170000 84.860000 21.370000 85.060000 ;
        RECT 21.170000 85.325000 21.370000 85.525000 ;
        RECT 21.245000 68.125000 21.445000 68.325000 ;
        RECT 21.245000 68.535000 21.445000 68.735000 ;
        RECT 21.245000 68.945000 21.445000 69.145000 ;
        RECT 21.245000 69.355000 21.445000 69.555000 ;
        RECT 21.245000 69.765000 21.445000 69.965000 ;
        RECT 21.245000 70.175000 21.445000 70.375000 ;
        RECT 21.245000 70.585000 21.445000 70.785000 ;
        RECT 21.245000 70.995000 21.445000 71.195000 ;
        RECT 21.245000 71.405000 21.445000 71.605000 ;
        RECT 21.245000 71.815000 21.445000 72.015000 ;
        RECT 21.245000 72.225000 21.445000 72.425000 ;
        RECT 21.245000 72.635000 21.445000 72.835000 ;
        RECT 21.245000 73.045000 21.445000 73.245000 ;
        RECT 21.245000 73.450000 21.445000 73.650000 ;
        RECT 21.245000 73.855000 21.445000 74.055000 ;
        RECT 21.245000 74.260000 21.445000 74.460000 ;
        RECT 21.245000 74.665000 21.445000 74.865000 ;
        RECT 21.245000 75.070000 21.445000 75.270000 ;
        RECT 21.245000 75.475000 21.445000 75.675000 ;
        RECT 21.245000 75.880000 21.445000 76.080000 ;
        RECT 21.245000 76.285000 21.445000 76.485000 ;
        RECT 21.245000 76.690000 21.445000 76.890000 ;
        RECT 21.245000 77.095000 21.445000 77.295000 ;
        RECT 21.245000 77.500000 21.445000 77.700000 ;
        RECT 21.245000 77.905000 21.445000 78.105000 ;
        RECT 21.245000 78.310000 21.445000 78.510000 ;
        RECT 21.245000 78.715000 21.445000 78.915000 ;
        RECT 21.245000 79.120000 21.445000 79.320000 ;
        RECT 21.245000 79.525000 21.445000 79.725000 ;
        RECT 21.245000 79.930000 21.445000 80.130000 ;
        RECT 21.245000 80.335000 21.445000 80.535000 ;
        RECT 21.245000 80.740000 21.445000 80.940000 ;
        RECT 21.245000 81.145000 21.445000 81.345000 ;
        RECT 21.245000 81.550000 21.445000 81.750000 ;
        RECT 21.245000 81.955000 21.445000 82.155000 ;
        RECT 21.245000 82.360000 21.445000 82.560000 ;
        RECT 21.345000 17.860000 21.545000 18.060000 ;
        RECT 21.345000 18.290000 21.545000 18.490000 ;
        RECT 21.345000 18.720000 21.545000 18.920000 ;
        RECT 21.345000 19.150000 21.545000 19.350000 ;
        RECT 21.345000 19.580000 21.545000 19.780000 ;
        RECT 21.345000 20.010000 21.545000 20.210000 ;
        RECT 21.345000 20.440000 21.545000 20.640000 ;
        RECT 21.345000 20.870000 21.545000 21.070000 ;
        RECT 21.345000 21.300000 21.545000 21.500000 ;
        RECT 21.345000 21.730000 21.545000 21.930000 ;
        RECT 21.345000 22.160000 21.545000 22.360000 ;
        RECT 21.645000 68.125000 21.845000 68.325000 ;
        RECT 21.645000 68.535000 21.845000 68.735000 ;
        RECT 21.645000 68.945000 21.845000 69.145000 ;
        RECT 21.645000 69.355000 21.845000 69.555000 ;
        RECT 21.645000 69.765000 21.845000 69.965000 ;
        RECT 21.645000 70.175000 21.845000 70.375000 ;
        RECT 21.645000 70.585000 21.845000 70.785000 ;
        RECT 21.645000 70.995000 21.845000 71.195000 ;
        RECT 21.645000 71.405000 21.845000 71.605000 ;
        RECT 21.645000 71.815000 21.845000 72.015000 ;
        RECT 21.645000 72.225000 21.845000 72.425000 ;
        RECT 21.645000 72.635000 21.845000 72.835000 ;
        RECT 21.645000 73.045000 21.845000 73.245000 ;
        RECT 21.645000 73.450000 21.845000 73.650000 ;
        RECT 21.645000 73.855000 21.845000 74.055000 ;
        RECT 21.645000 74.260000 21.845000 74.460000 ;
        RECT 21.645000 74.665000 21.845000 74.865000 ;
        RECT 21.645000 75.070000 21.845000 75.270000 ;
        RECT 21.645000 75.475000 21.845000 75.675000 ;
        RECT 21.645000 75.880000 21.845000 76.080000 ;
        RECT 21.645000 76.285000 21.845000 76.485000 ;
        RECT 21.645000 76.690000 21.845000 76.890000 ;
        RECT 21.645000 77.095000 21.845000 77.295000 ;
        RECT 21.645000 77.500000 21.845000 77.700000 ;
        RECT 21.645000 77.905000 21.845000 78.105000 ;
        RECT 21.645000 78.310000 21.845000 78.510000 ;
        RECT 21.645000 78.715000 21.845000 78.915000 ;
        RECT 21.645000 79.120000 21.845000 79.320000 ;
        RECT 21.645000 79.525000 21.845000 79.725000 ;
        RECT 21.645000 79.930000 21.845000 80.130000 ;
        RECT 21.645000 80.335000 21.845000 80.535000 ;
        RECT 21.645000 80.740000 21.845000 80.940000 ;
        RECT 21.645000 81.145000 21.845000 81.345000 ;
        RECT 21.645000 81.550000 21.845000 81.750000 ;
        RECT 21.645000 81.955000 21.845000 82.155000 ;
        RECT 21.645000 82.360000 21.845000 82.560000 ;
        RECT 21.715000 82.920000 21.915000 83.120000 ;
        RECT 21.715000 83.470000 21.915000 83.670000 ;
        RECT 21.715000 84.020000 21.915000 84.220000 ;
        RECT 21.750000 17.860000 21.950000 18.060000 ;
        RECT 21.750000 18.290000 21.950000 18.490000 ;
        RECT 21.750000 18.720000 21.950000 18.920000 ;
        RECT 21.750000 19.150000 21.950000 19.350000 ;
        RECT 21.750000 19.580000 21.950000 19.780000 ;
        RECT 21.750000 20.010000 21.950000 20.210000 ;
        RECT 21.750000 20.440000 21.950000 20.640000 ;
        RECT 21.750000 20.870000 21.950000 21.070000 ;
        RECT 21.750000 21.300000 21.950000 21.500000 ;
        RECT 21.750000 21.730000 21.950000 21.930000 ;
        RECT 21.750000 22.160000 21.950000 22.360000 ;
        RECT 22.045000 68.125000 22.245000 68.325000 ;
        RECT 22.045000 68.535000 22.245000 68.735000 ;
        RECT 22.045000 68.945000 22.245000 69.145000 ;
        RECT 22.045000 69.355000 22.245000 69.555000 ;
        RECT 22.045000 69.765000 22.245000 69.965000 ;
        RECT 22.045000 70.175000 22.245000 70.375000 ;
        RECT 22.045000 70.585000 22.245000 70.785000 ;
        RECT 22.045000 70.995000 22.245000 71.195000 ;
        RECT 22.045000 71.405000 22.245000 71.605000 ;
        RECT 22.045000 71.815000 22.245000 72.015000 ;
        RECT 22.045000 72.225000 22.245000 72.425000 ;
        RECT 22.045000 72.635000 22.245000 72.835000 ;
        RECT 22.045000 73.045000 22.245000 73.245000 ;
        RECT 22.045000 73.450000 22.245000 73.650000 ;
        RECT 22.045000 73.855000 22.245000 74.055000 ;
        RECT 22.045000 74.260000 22.245000 74.460000 ;
        RECT 22.045000 74.665000 22.245000 74.865000 ;
        RECT 22.045000 75.070000 22.245000 75.270000 ;
        RECT 22.045000 75.475000 22.245000 75.675000 ;
        RECT 22.045000 75.880000 22.245000 76.080000 ;
        RECT 22.045000 76.285000 22.245000 76.485000 ;
        RECT 22.045000 76.690000 22.245000 76.890000 ;
        RECT 22.045000 77.095000 22.245000 77.295000 ;
        RECT 22.045000 77.500000 22.245000 77.700000 ;
        RECT 22.045000 77.905000 22.245000 78.105000 ;
        RECT 22.045000 78.310000 22.245000 78.510000 ;
        RECT 22.045000 78.715000 22.245000 78.915000 ;
        RECT 22.045000 79.120000 22.245000 79.320000 ;
        RECT 22.045000 79.525000 22.245000 79.725000 ;
        RECT 22.045000 79.930000 22.245000 80.130000 ;
        RECT 22.045000 80.335000 22.245000 80.535000 ;
        RECT 22.045000 80.740000 22.245000 80.940000 ;
        RECT 22.045000 81.145000 22.245000 81.345000 ;
        RECT 22.045000 81.550000 22.245000 81.750000 ;
        RECT 22.045000 81.955000 22.245000 82.155000 ;
        RECT 22.045000 82.360000 22.245000 82.560000 ;
        RECT 22.160000 17.860000 22.360000 18.060000 ;
        RECT 22.160000 18.290000 22.360000 18.490000 ;
        RECT 22.160000 18.720000 22.360000 18.920000 ;
        RECT 22.160000 19.150000 22.360000 19.350000 ;
        RECT 22.160000 19.580000 22.360000 19.780000 ;
        RECT 22.160000 20.010000 22.360000 20.210000 ;
        RECT 22.160000 20.440000 22.360000 20.640000 ;
        RECT 22.160000 20.870000 22.360000 21.070000 ;
        RECT 22.160000 21.300000 22.360000 21.500000 ;
        RECT 22.160000 21.730000 22.360000 21.930000 ;
        RECT 22.160000 22.160000 22.360000 22.360000 ;
        RECT 22.445000 68.125000 22.645000 68.325000 ;
        RECT 22.445000 68.535000 22.645000 68.735000 ;
        RECT 22.445000 68.945000 22.645000 69.145000 ;
        RECT 22.445000 69.355000 22.645000 69.555000 ;
        RECT 22.445000 69.765000 22.645000 69.965000 ;
        RECT 22.445000 70.175000 22.645000 70.375000 ;
        RECT 22.445000 70.585000 22.645000 70.785000 ;
        RECT 22.445000 70.995000 22.645000 71.195000 ;
        RECT 22.445000 71.405000 22.645000 71.605000 ;
        RECT 22.445000 71.815000 22.645000 72.015000 ;
        RECT 22.445000 72.225000 22.645000 72.425000 ;
        RECT 22.445000 72.635000 22.645000 72.835000 ;
        RECT 22.445000 73.045000 22.645000 73.245000 ;
        RECT 22.445000 73.450000 22.645000 73.650000 ;
        RECT 22.445000 73.855000 22.645000 74.055000 ;
        RECT 22.445000 74.260000 22.645000 74.460000 ;
        RECT 22.445000 74.665000 22.645000 74.865000 ;
        RECT 22.445000 75.070000 22.645000 75.270000 ;
        RECT 22.445000 75.475000 22.645000 75.675000 ;
        RECT 22.445000 75.880000 22.645000 76.080000 ;
        RECT 22.445000 76.285000 22.645000 76.485000 ;
        RECT 22.445000 76.690000 22.645000 76.890000 ;
        RECT 22.445000 77.095000 22.645000 77.295000 ;
        RECT 22.445000 77.500000 22.645000 77.700000 ;
        RECT 22.445000 77.905000 22.645000 78.105000 ;
        RECT 22.445000 78.310000 22.645000 78.510000 ;
        RECT 22.445000 78.715000 22.645000 78.915000 ;
        RECT 22.445000 79.120000 22.645000 79.320000 ;
        RECT 22.445000 79.525000 22.645000 79.725000 ;
        RECT 22.445000 79.930000 22.645000 80.130000 ;
        RECT 22.445000 80.335000 22.645000 80.535000 ;
        RECT 22.445000 80.740000 22.645000 80.940000 ;
        RECT 22.445000 81.145000 22.645000 81.345000 ;
        RECT 22.445000 81.550000 22.645000 81.750000 ;
        RECT 22.445000 81.955000 22.645000 82.155000 ;
        RECT 22.445000 82.360000 22.645000 82.560000 ;
        RECT 22.505000 82.920000 22.705000 83.120000 ;
        RECT 22.505000 83.470000 22.705000 83.670000 ;
        RECT 22.505000 84.020000 22.705000 84.220000 ;
        RECT 22.570000 17.860000 22.770000 18.060000 ;
        RECT 22.570000 18.290000 22.770000 18.490000 ;
        RECT 22.570000 18.720000 22.770000 18.920000 ;
        RECT 22.570000 19.150000 22.770000 19.350000 ;
        RECT 22.570000 19.580000 22.770000 19.780000 ;
        RECT 22.570000 20.010000 22.770000 20.210000 ;
        RECT 22.570000 20.440000 22.770000 20.640000 ;
        RECT 22.570000 20.870000 22.770000 21.070000 ;
        RECT 22.570000 21.300000 22.770000 21.500000 ;
        RECT 22.570000 21.730000 22.770000 21.930000 ;
        RECT 22.570000 22.160000 22.770000 22.360000 ;
        RECT 22.845000 68.125000 23.045000 68.325000 ;
        RECT 22.845000 68.535000 23.045000 68.735000 ;
        RECT 22.845000 68.945000 23.045000 69.145000 ;
        RECT 22.845000 69.355000 23.045000 69.555000 ;
        RECT 22.845000 69.765000 23.045000 69.965000 ;
        RECT 22.845000 70.175000 23.045000 70.375000 ;
        RECT 22.845000 70.585000 23.045000 70.785000 ;
        RECT 22.845000 70.995000 23.045000 71.195000 ;
        RECT 22.845000 71.405000 23.045000 71.605000 ;
        RECT 22.845000 71.815000 23.045000 72.015000 ;
        RECT 22.845000 72.225000 23.045000 72.425000 ;
        RECT 22.845000 72.635000 23.045000 72.835000 ;
        RECT 22.845000 73.045000 23.045000 73.245000 ;
        RECT 22.845000 73.450000 23.045000 73.650000 ;
        RECT 22.845000 73.855000 23.045000 74.055000 ;
        RECT 22.845000 74.260000 23.045000 74.460000 ;
        RECT 22.845000 74.665000 23.045000 74.865000 ;
        RECT 22.845000 75.070000 23.045000 75.270000 ;
        RECT 22.845000 75.475000 23.045000 75.675000 ;
        RECT 22.845000 75.880000 23.045000 76.080000 ;
        RECT 22.845000 76.285000 23.045000 76.485000 ;
        RECT 22.845000 76.690000 23.045000 76.890000 ;
        RECT 22.845000 77.095000 23.045000 77.295000 ;
        RECT 22.845000 77.500000 23.045000 77.700000 ;
        RECT 22.845000 77.905000 23.045000 78.105000 ;
        RECT 22.845000 78.310000 23.045000 78.510000 ;
        RECT 22.845000 78.715000 23.045000 78.915000 ;
        RECT 22.845000 79.120000 23.045000 79.320000 ;
        RECT 22.845000 79.525000 23.045000 79.725000 ;
        RECT 22.845000 79.930000 23.045000 80.130000 ;
        RECT 22.845000 80.335000 23.045000 80.535000 ;
        RECT 22.845000 80.740000 23.045000 80.940000 ;
        RECT 22.845000 81.145000 23.045000 81.345000 ;
        RECT 22.845000 81.550000 23.045000 81.750000 ;
        RECT 22.845000 81.955000 23.045000 82.155000 ;
        RECT 22.845000 82.360000 23.045000 82.560000 ;
        RECT 22.980000 17.860000 23.180000 18.060000 ;
        RECT 22.980000 18.290000 23.180000 18.490000 ;
        RECT 22.980000 18.720000 23.180000 18.920000 ;
        RECT 22.980000 19.150000 23.180000 19.350000 ;
        RECT 22.980000 19.580000 23.180000 19.780000 ;
        RECT 22.980000 20.010000 23.180000 20.210000 ;
        RECT 22.980000 20.440000 23.180000 20.640000 ;
        RECT 22.980000 20.870000 23.180000 21.070000 ;
        RECT 22.980000 21.300000 23.180000 21.500000 ;
        RECT 22.980000 21.730000 23.180000 21.930000 ;
        RECT 22.980000 22.160000 23.180000 22.360000 ;
        RECT 23.245000 68.125000 23.445000 68.325000 ;
        RECT 23.245000 68.535000 23.445000 68.735000 ;
        RECT 23.245000 68.945000 23.445000 69.145000 ;
        RECT 23.245000 69.355000 23.445000 69.555000 ;
        RECT 23.245000 69.765000 23.445000 69.965000 ;
        RECT 23.245000 70.175000 23.445000 70.375000 ;
        RECT 23.245000 70.585000 23.445000 70.785000 ;
        RECT 23.245000 70.995000 23.445000 71.195000 ;
        RECT 23.245000 71.405000 23.445000 71.605000 ;
        RECT 23.245000 71.815000 23.445000 72.015000 ;
        RECT 23.245000 72.225000 23.445000 72.425000 ;
        RECT 23.245000 72.635000 23.445000 72.835000 ;
        RECT 23.245000 73.045000 23.445000 73.245000 ;
        RECT 23.245000 73.450000 23.445000 73.650000 ;
        RECT 23.245000 73.855000 23.445000 74.055000 ;
        RECT 23.245000 74.260000 23.445000 74.460000 ;
        RECT 23.245000 74.665000 23.445000 74.865000 ;
        RECT 23.245000 75.070000 23.445000 75.270000 ;
        RECT 23.245000 75.475000 23.445000 75.675000 ;
        RECT 23.245000 75.880000 23.445000 76.080000 ;
        RECT 23.245000 76.285000 23.445000 76.485000 ;
        RECT 23.245000 76.690000 23.445000 76.890000 ;
        RECT 23.245000 77.095000 23.445000 77.295000 ;
        RECT 23.245000 77.500000 23.445000 77.700000 ;
        RECT 23.245000 77.905000 23.445000 78.105000 ;
        RECT 23.245000 78.310000 23.445000 78.510000 ;
        RECT 23.245000 78.715000 23.445000 78.915000 ;
        RECT 23.245000 79.120000 23.445000 79.320000 ;
        RECT 23.245000 79.525000 23.445000 79.725000 ;
        RECT 23.245000 79.930000 23.445000 80.130000 ;
        RECT 23.245000 80.335000 23.445000 80.535000 ;
        RECT 23.245000 80.740000 23.445000 80.940000 ;
        RECT 23.245000 81.145000 23.445000 81.345000 ;
        RECT 23.245000 81.550000 23.445000 81.750000 ;
        RECT 23.245000 81.955000 23.445000 82.155000 ;
        RECT 23.245000 82.360000 23.445000 82.560000 ;
        RECT 23.390000 17.860000 23.590000 18.060000 ;
        RECT 23.390000 18.290000 23.590000 18.490000 ;
        RECT 23.390000 18.720000 23.590000 18.920000 ;
        RECT 23.390000 19.150000 23.590000 19.350000 ;
        RECT 23.390000 19.580000 23.590000 19.780000 ;
        RECT 23.390000 20.010000 23.590000 20.210000 ;
        RECT 23.390000 20.440000 23.590000 20.640000 ;
        RECT 23.390000 20.870000 23.590000 21.070000 ;
        RECT 23.390000 21.300000 23.590000 21.500000 ;
        RECT 23.390000 21.730000 23.590000 21.930000 ;
        RECT 23.390000 22.160000 23.590000 22.360000 ;
        RECT 23.645000 68.125000 23.845000 68.325000 ;
        RECT 23.645000 68.535000 23.845000 68.735000 ;
        RECT 23.645000 68.945000 23.845000 69.145000 ;
        RECT 23.645000 69.355000 23.845000 69.555000 ;
        RECT 23.645000 69.765000 23.845000 69.965000 ;
        RECT 23.645000 70.175000 23.845000 70.375000 ;
        RECT 23.645000 70.585000 23.845000 70.785000 ;
        RECT 23.645000 70.995000 23.845000 71.195000 ;
        RECT 23.645000 71.405000 23.845000 71.605000 ;
        RECT 23.645000 71.815000 23.845000 72.015000 ;
        RECT 23.645000 72.225000 23.845000 72.425000 ;
        RECT 23.645000 72.635000 23.845000 72.835000 ;
        RECT 23.645000 73.045000 23.845000 73.245000 ;
        RECT 23.645000 73.450000 23.845000 73.650000 ;
        RECT 23.645000 73.855000 23.845000 74.055000 ;
        RECT 23.645000 74.260000 23.845000 74.460000 ;
        RECT 23.645000 74.665000 23.845000 74.865000 ;
        RECT 23.645000 75.070000 23.845000 75.270000 ;
        RECT 23.645000 75.475000 23.845000 75.675000 ;
        RECT 23.645000 75.880000 23.845000 76.080000 ;
        RECT 23.645000 76.285000 23.845000 76.485000 ;
        RECT 23.645000 76.690000 23.845000 76.890000 ;
        RECT 23.645000 77.095000 23.845000 77.295000 ;
        RECT 23.645000 77.500000 23.845000 77.700000 ;
        RECT 23.645000 77.905000 23.845000 78.105000 ;
        RECT 23.645000 78.310000 23.845000 78.510000 ;
        RECT 23.645000 78.715000 23.845000 78.915000 ;
        RECT 23.645000 79.120000 23.845000 79.320000 ;
        RECT 23.645000 79.525000 23.845000 79.725000 ;
        RECT 23.645000 79.930000 23.845000 80.130000 ;
        RECT 23.645000 80.335000 23.845000 80.535000 ;
        RECT 23.645000 80.740000 23.845000 80.940000 ;
        RECT 23.645000 81.145000 23.845000 81.345000 ;
        RECT 23.645000 81.550000 23.845000 81.750000 ;
        RECT 23.645000 81.955000 23.845000 82.155000 ;
        RECT 23.645000 82.360000 23.845000 82.560000 ;
        RECT 23.800000 17.860000 24.000000 18.060000 ;
        RECT 23.800000 18.290000 24.000000 18.490000 ;
        RECT 23.800000 18.720000 24.000000 18.920000 ;
        RECT 23.800000 19.150000 24.000000 19.350000 ;
        RECT 23.800000 19.580000 24.000000 19.780000 ;
        RECT 23.800000 20.010000 24.000000 20.210000 ;
        RECT 23.800000 20.440000 24.000000 20.640000 ;
        RECT 23.800000 20.870000 24.000000 21.070000 ;
        RECT 23.800000 21.300000 24.000000 21.500000 ;
        RECT 23.800000 21.730000 24.000000 21.930000 ;
        RECT 23.800000 22.160000 24.000000 22.360000 ;
        RECT 24.045000 68.125000 24.245000 68.325000 ;
        RECT 24.045000 68.535000 24.245000 68.735000 ;
        RECT 24.045000 68.945000 24.245000 69.145000 ;
        RECT 24.045000 69.355000 24.245000 69.555000 ;
        RECT 24.045000 69.765000 24.245000 69.965000 ;
        RECT 24.045000 70.175000 24.245000 70.375000 ;
        RECT 24.045000 70.585000 24.245000 70.785000 ;
        RECT 24.045000 70.995000 24.245000 71.195000 ;
        RECT 24.045000 71.405000 24.245000 71.605000 ;
        RECT 24.045000 71.815000 24.245000 72.015000 ;
        RECT 24.045000 72.225000 24.245000 72.425000 ;
        RECT 24.045000 72.635000 24.245000 72.835000 ;
        RECT 24.045000 73.045000 24.245000 73.245000 ;
        RECT 24.045000 73.450000 24.245000 73.650000 ;
        RECT 24.045000 73.855000 24.245000 74.055000 ;
        RECT 24.045000 74.260000 24.245000 74.460000 ;
        RECT 24.045000 74.665000 24.245000 74.865000 ;
        RECT 24.045000 75.070000 24.245000 75.270000 ;
        RECT 24.045000 75.475000 24.245000 75.675000 ;
        RECT 24.045000 75.880000 24.245000 76.080000 ;
        RECT 24.045000 76.285000 24.245000 76.485000 ;
        RECT 24.045000 76.690000 24.245000 76.890000 ;
        RECT 24.045000 77.095000 24.245000 77.295000 ;
        RECT 24.045000 77.500000 24.245000 77.700000 ;
        RECT 24.045000 77.905000 24.245000 78.105000 ;
        RECT 24.045000 78.310000 24.245000 78.510000 ;
        RECT 24.045000 78.715000 24.245000 78.915000 ;
        RECT 24.045000 79.120000 24.245000 79.320000 ;
        RECT 24.045000 79.525000 24.245000 79.725000 ;
        RECT 24.045000 79.930000 24.245000 80.130000 ;
        RECT 24.045000 80.335000 24.245000 80.535000 ;
        RECT 24.045000 80.740000 24.245000 80.940000 ;
        RECT 24.045000 81.145000 24.245000 81.345000 ;
        RECT 24.045000 81.550000 24.245000 81.750000 ;
        RECT 24.045000 81.955000 24.245000 82.155000 ;
        RECT 24.045000 82.360000 24.245000 82.560000 ;
        RECT 24.210000 17.860000 24.410000 18.060000 ;
        RECT 24.210000 18.290000 24.410000 18.490000 ;
        RECT 24.210000 18.720000 24.410000 18.920000 ;
        RECT 24.210000 19.150000 24.410000 19.350000 ;
        RECT 24.210000 19.580000 24.410000 19.780000 ;
        RECT 24.210000 20.010000 24.410000 20.210000 ;
        RECT 24.210000 20.440000 24.410000 20.640000 ;
        RECT 24.210000 20.870000 24.410000 21.070000 ;
        RECT 24.210000 21.300000 24.410000 21.500000 ;
        RECT 24.210000 21.730000 24.410000 21.930000 ;
        RECT 24.210000 22.160000 24.410000 22.360000 ;
        RECT 50.845000 17.860000 51.045000 18.060000 ;
        RECT 50.845000 18.290000 51.045000 18.490000 ;
        RECT 50.845000 18.720000 51.045000 18.920000 ;
        RECT 50.845000 19.150000 51.045000 19.350000 ;
        RECT 50.845000 19.580000 51.045000 19.780000 ;
        RECT 50.845000 20.010000 51.045000 20.210000 ;
        RECT 50.845000 20.440000 51.045000 20.640000 ;
        RECT 50.845000 20.870000 51.045000 21.070000 ;
        RECT 50.845000 21.300000 51.045000 21.500000 ;
        RECT 50.845000 21.730000 51.045000 21.930000 ;
        RECT 50.845000 22.160000 51.045000 22.360000 ;
        RECT 51.010000 68.125000 51.210000 68.325000 ;
        RECT 51.010000 68.535000 51.210000 68.735000 ;
        RECT 51.010000 68.945000 51.210000 69.145000 ;
        RECT 51.010000 69.355000 51.210000 69.555000 ;
        RECT 51.010000 69.765000 51.210000 69.965000 ;
        RECT 51.010000 70.175000 51.210000 70.375000 ;
        RECT 51.010000 70.585000 51.210000 70.785000 ;
        RECT 51.010000 70.995000 51.210000 71.195000 ;
        RECT 51.010000 71.405000 51.210000 71.605000 ;
        RECT 51.010000 71.815000 51.210000 72.015000 ;
        RECT 51.010000 72.225000 51.210000 72.425000 ;
        RECT 51.010000 72.635000 51.210000 72.835000 ;
        RECT 51.010000 73.045000 51.210000 73.245000 ;
        RECT 51.010000 73.450000 51.210000 73.650000 ;
        RECT 51.010000 73.855000 51.210000 74.055000 ;
        RECT 51.010000 74.260000 51.210000 74.460000 ;
        RECT 51.010000 74.665000 51.210000 74.865000 ;
        RECT 51.010000 75.070000 51.210000 75.270000 ;
        RECT 51.010000 75.475000 51.210000 75.675000 ;
        RECT 51.010000 75.880000 51.210000 76.080000 ;
        RECT 51.010000 76.285000 51.210000 76.485000 ;
        RECT 51.010000 76.690000 51.210000 76.890000 ;
        RECT 51.010000 77.095000 51.210000 77.295000 ;
        RECT 51.010000 77.500000 51.210000 77.700000 ;
        RECT 51.010000 77.905000 51.210000 78.105000 ;
        RECT 51.010000 78.310000 51.210000 78.510000 ;
        RECT 51.010000 78.715000 51.210000 78.915000 ;
        RECT 51.010000 79.120000 51.210000 79.320000 ;
        RECT 51.010000 79.525000 51.210000 79.725000 ;
        RECT 51.010000 79.930000 51.210000 80.130000 ;
        RECT 51.010000 80.335000 51.210000 80.535000 ;
        RECT 51.010000 80.740000 51.210000 80.940000 ;
        RECT 51.010000 81.145000 51.210000 81.345000 ;
        RECT 51.010000 81.550000 51.210000 81.750000 ;
        RECT 51.010000 81.955000 51.210000 82.155000 ;
        RECT 51.010000 82.360000 51.210000 82.560000 ;
        RECT 51.250000 17.860000 51.450000 18.060000 ;
        RECT 51.250000 18.290000 51.450000 18.490000 ;
        RECT 51.250000 18.720000 51.450000 18.920000 ;
        RECT 51.250000 19.150000 51.450000 19.350000 ;
        RECT 51.250000 19.580000 51.450000 19.780000 ;
        RECT 51.250000 20.010000 51.450000 20.210000 ;
        RECT 51.250000 20.440000 51.450000 20.640000 ;
        RECT 51.250000 20.870000 51.450000 21.070000 ;
        RECT 51.250000 21.300000 51.450000 21.500000 ;
        RECT 51.250000 21.730000 51.450000 21.930000 ;
        RECT 51.250000 22.160000 51.450000 22.360000 ;
        RECT 51.410000 68.125000 51.610000 68.325000 ;
        RECT 51.410000 68.535000 51.610000 68.735000 ;
        RECT 51.410000 68.945000 51.610000 69.145000 ;
        RECT 51.410000 69.355000 51.610000 69.555000 ;
        RECT 51.410000 69.765000 51.610000 69.965000 ;
        RECT 51.410000 70.175000 51.610000 70.375000 ;
        RECT 51.410000 70.585000 51.610000 70.785000 ;
        RECT 51.410000 70.995000 51.610000 71.195000 ;
        RECT 51.410000 71.405000 51.610000 71.605000 ;
        RECT 51.410000 71.815000 51.610000 72.015000 ;
        RECT 51.410000 72.225000 51.610000 72.425000 ;
        RECT 51.410000 72.635000 51.610000 72.835000 ;
        RECT 51.410000 73.045000 51.610000 73.245000 ;
        RECT 51.410000 73.450000 51.610000 73.650000 ;
        RECT 51.410000 73.855000 51.610000 74.055000 ;
        RECT 51.410000 74.260000 51.610000 74.460000 ;
        RECT 51.410000 74.665000 51.610000 74.865000 ;
        RECT 51.410000 75.070000 51.610000 75.270000 ;
        RECT 51.410000 75.475000 51.610000 75.675000 ;
        RECT 51.410000 75.880000 51.610000 76.080000 ;
        RECT 51.410000 76.285000 51.610000 76.485000 ;
        RECT 51.410000 76.690000 51.610000 76.890000 ;
        RECT 51.410000 77.095000 51.610000 77.295000 ;
        RECT 51.410000 77.500000 51.610000 77.700000 ;
        RECT 51.410000 77.905000 51.610000 78.105000 ;
        RECT 51.410000 78.310000 51.610000 78.510000 ;
        RECT 51.410000 78.715000 51.610000 78.915000 ;
        RECT 51.410000 79.120000 51.610000 79.320000 ;
        RECT 51.410000 79.525000 51.610000 79.725000 ;
        RECT 51.410000 79.930000 51.610000 80.130000 ;
        RECT 51.410000 80.335000 51.610000 80.535000 ;
        RECT 51.410000 80.740000 51.610000 80.940000 ;
        RECT 51.410000 81.145000 51.610000 81.345000 ;
        RECT 51.410000 81.550000 51.610000 81.750000 ;
        RECT 51.410000 81.955000 51.610000 82.155000 ;
        RECT 51.410000 82.360000 51.610000 82.560000 ;
        RECT 51.655000 17.860000 51.855000 18.060000 ;
        RECT 51.655000 18.290000 51.855000 18.490000 ;
        RECT 51.655000 18.720000 51.855000 18.920000 ;
        RECT 51.655000 19.150000 51.855000 19.350000 ;
        RECT 51.655000 19.580000 51.855000 19.780000 ;
        RECT 51.655000 20.010000 51.855000 20.210000 ;
        RECT 51.655000 20.440000 51.855000 20.640000 ;
        RECT 51.655000 20.870000 51.855000 21.070000 ;
        RECT 51.655000 21.300000 51.855000 21.500000 ;
        RECT 51.655000 21.730000 51.855000 21.930000 ;
        RECT 51.655000 22.160000 51.855000 22.360000 ;
        RECT 51.810000 68.125000 52.010000 68.325000 ;
        RECT 51.810000 68.535000 52.010000 68.735000 ;
        RECT 51.810000 68.945000 52.010000 69.145000 ;
        RECT 51.810000 69.355000 52.010000 69.555000 ;
        RECT 51.810000 69.765000 52.010000 69.965000 ;
        RECT 51.810000 70.175000 52.010000 70.375000 ;
        RECT 51.810000 70.585000 52.010000 70.785000 ;
        RECT 51.810000 70.995000 52.010000 71.195000 ;
        RECT 51.810000 71.405000 52.010000 71.605000 ;
        RECT 51.810000 71.815000 52.010000 72.015000 ;
        RECT 51.810000 72.225000 52.010000 72.425000 ;
        RECT 51.810000 72.635000 52.010000 72.835000 ;
        RECT 51.810000 73.045000 52.010000 73.245000 ;
        RECT 51.810000 73.450000 52.010000 73.650000 ;
        RECT 51.810000 73.855000 52.010000 74.055000 ;
        RECT 51.810000 74.260000 52.010000 74.460000 ;
        RECT 51.810000 74.665000 52.010000 74.865000 ;
        RECT 51.810000 75.070000 52.010000 75.270000 ;
        RECT 51.810000 75.475000 52.010000 75.675000 ;
        RECT 51.810000 75.880000 52.010000 76.080000 ;
        RECT 51.810000 76.285000 52.010000 76.485000 ;
        RECT 51.810000 76.690000 52.010000 76.890000 ;
        RECT 51.810000 77.095000 52.010000 77.295000 ;
        RECT 51.810000 77.500000 52.010000 77.700000 ;
        RECT 51.810000 77.905000 52.010000 78.105000 ;
        RECT 51.810000 78.310000 52.010000 78.510000 ;
        RECT 51.810000 78.715000 52.010000 78.915000 ;
        RECT 51.810000 79.120000 52.010000 79.320000 ;
        RECT 51.810000 79.525000 52.010000 79.725000 ;
        RECT 51.810000 79.930000 52.010000 80.130000 ;
        RECT 51.810000 80.335000 52.010000 80.535000 ;
        RECT 51.810000 80.740000 52.010000 80.940000 ;
        RECT 51.810000 81.145000 52.010000 81.345000 ;
        RECT 51.810000 81.550000 52.010000 81.750000 ;
        RECT 51.810000 81.955000 52.010000 82.155000 ;
        RECT 51.810000 82.360000 52.010000 82.560000 ;
        RECT 52.060000 17.860000 52.260000 18.060000 ;
        RECT 52.060000 18.290000 52.260000 18.490000 ;
        RECT 52.060000 18.720000 52.260000 18.920000 ;
        RECT 52.060000 19.150000 52.260000 19.350000 ;
        RECT 52.060000 19.580000 52.260000 19.780000 ;
        RECT 52.060000 20.010000 52.260000 20.210000 ;
        RECT 52.060000 20.440000 52.260000 20.640000 ;
        RECT 52.060000 20.870000 52.260000 21.070000 ;
        RECT 52.060000 21.300000 52.260000 21.500000 ;
        RECT 52.060000 21.730000 52.260000 21.930000 ;
        RECT 52.060000 22.160000 52.260000 22.360000 ;
        RECT 52.210000 68.125000 52.410000 68.325000 ;
        RECT 52.210000 68.535000 52.410000 68.735000 ;
        RECT 52.210000 68.945000 52.410000 69.145000 ;
        RECT 52.210000 69.355000 52.410000 69.555000 ;
        RECT 52.210000 69.765000 52.410000 69.965000 ;
        RECT 52.210000 70.175000 52.410000 70.375000 ;
        RECT 52.210000 70.585000 52.410000 70.785000 ;
        RECT 52.210000 70.995000 52.410000 71.195000 ;
        RECT 52.210000 71.405000 52.410000 71.605000 ;
        RECT 52.210000 71.815000 52.410000 72.015000 ;
        RECT 52.210000 72.225000 52.410000 72.425000 ;
        RECT 52.210000 72.635000 52.410000 72.835000 ;
        RECT 52.210000 73.045000 52.410000 73.245000 ;
        RECT 52.210000 73.450000 52.410000 73.650000 ;
        RECT 52.210000 73.855000 52.410000 74.055000 ;
        RECT 52.210000 74.260000 52.410000 74.460000 ;
        RECT 52.210000 74.665000 52.410000 74.865000 ;
        RECT 52.210000 75.070000 52.410000 75.270000 ;
        RECT 52.210000 75.475000 52.410000 75.675000 ;
        RECT 52.210000 75.880000 52.410000 76.080000 ;
        RECT 52.210000 76.285000 52.410000 76.485000 ;
        RECT 52.210000 76.690000 52.410000 76.890000 ;
        RECT 52.210000 77.095000 52.410000 77.295000 ;
        RECT 52.210000 77.500000 52.410000 77.700000 ;
        RECT 52.210000 77.905000 52.410000 78.105000 ;
        RECT 52.210000 78.310000 52.410000 78.510000 ;
        RECT 52.210000 78.715000 52.410000 78.915000 ;
        RECT 52.210000 79.120000 52.410000 79.320000 ;
        RECT 52.210000 79.525000 52.410000 79.725000 ;
        RECT 52.210000 79.930000 52.410000 80.130000 ;
        RECT 52.210000 80.335000 52.410000 80.535000 ;
        RECT 52.210000 80.740000 52.410000 80.940000 ;
        RECT 52.210000 81.145000 52.410000 81.345000 ;
        RECT 52.210000 81.550000 52.410000 81.750000 ;
        RECT 52.210000 81.955000 52.410000 82.155000 ;
        RECT 52.210000 82.360000 52.410000 82.560000 ;
        RECT 52.465000 17.860000 52.665000 18.060000 ;
        RECT 52.465000 18.290000 52.665000 18.490000 ;
        RECT 52.465000 18.720000 52.665000 18.920000 ;
        RECT 52.465000 19.150000 52.665000 19.350000 ;
        RECT 52.465000 19.580000 52.665000 19.780000 ;
        RECT 52.465000 20.010000 52.665000 20.210000 ;
        RECT 52.465000 20.440000 52.665000 20.640000 ;
        RECT 52.465000 20.870000 52.665000 21.070000 ;
        RECT 52.465000 21.300000 52.665000 21.500000 ;
        RECT 52.465000 21.730000 52.665000 21.930000 ;
        RECT 52.465000 22.160000 52.665000 22.360000 ;
        RECT 52.550000 82.920000 52.750000 83.120000 ;
        RECT 52.550000 83.470000 52.750000 83.670000 ;
        RECT 52.550000 84.020000 52.750000 84.220000 ;
        RECT 52.610000 68.125000 52.810000 68.325000 ;
        RECT 52.610000 68.535000 52.810000 68.735000 ;
        RECT 52.610000 68.945000 52.810000 69.145000 ;
        RECT 52.610000 69.355000 52.810000 69.555000 ;
        RECT 52.610000 69.765000 52.810000 69.965000 ;
        RECT 52.610000 70.175000 52.810000 70.375000 ;
        RECT 52.610000 70.585000 52.810000 70.785000 ;
        RECT 52.610000 70.995000 52.810000 71.195000 ;
        RECT 52.610000 71.405000 52.810000 71.605000 ;
        RECT 52.610000 71.815000 52.810000 72.015000 ;
        RECT 52.610000 72.225000 52.810000 72.425000 ;
        RECT 52.610000 72.635000 52.810000 72.835000 ;
        RECT 52.610000 73.045000 52.810000 73.245000 ;
        RECT 52.610000 73.450000 52.810000 73.650000 ;
        RECT 52.610000 73.855000 52.810000 74.055000 ;
        RECT 52.610000 74.260000 52.810000 74.460000 ;
        RECT 52.610000 74.665000 52.810000 74.865000 ;
        RECT 52.610000 75.070000 52.810000 75.270000 ;
        RECT 52.610000 75.475000 52.810000 75.675000 ;
        RECT 52.610000 75.880000 52.810000 76.080000 ;
        RECT 52.610000 76.285000 52.810000 76.485000 ;
        RECT 52.610000 76.690000 52.810000 76.890000 ;
        RECT 52.610000 77.095000 52.810000 77.295000 ;
        RECT 52.610000 77.500000 52.810000 77.700000 ;
        RECT 52.610000 77.905000 52.810000 78.105000 ;
        RECT 52.610000 78.310000 52.810000 78.510000 ;
        RECT 52.610000 78.715000 52.810000 78.915000 ;
        RECT 52.610000 79.120000 52.810000 79.320000 ;
        RECT 52.610000 79.525000 52.810000 79.725000 ;
        RECT 52.610000 79.930000 52.810000 80.130000 ;
        RECT 52.610000 80.335000 52.810000 80.535000 ;
        RECT 52.610000 80.740000 52.810000 80.940000 ;
        RECT 52.610000 81.145000 52.810000 81.345000 ;
        RECT 52.610000 81.550000 52.810000 81.750000 ;
        RECT 52.610000 81.955000 52.810000 82.155000 ;
        RECT 52.610000 82.360000 52.810000 82.560000 ;
        RECT 52.870000 17.860000 53.070000 18.060000 ;
        RECT 52.870000 18.290000 53.070000 18.490000 ;
        RECT 52.870000 18.720000 53.070000 18.920000 ;
        RECT 52.870000 19.150000 53.070000 19.350000 ;
        RECT 52.870000 19.580000 53.070000 19.780000 ;
        RECT 52.870000 20.010000 53.070000 20.210000 ;
        RECT 52.870000 20.440000 53.070000 20.640000 ;
        RECT 52.870000 20.870000 53.070000 21.070000 ;
        RECT 52.870000 21.300000 53.070000 21.500000 ;
        RECT 52.870000 21.730000 53.070000 21.930000 ;
        RECT 52.870000 22.160000 53.070000 22.360000 ;
        RECT 53.010000 68.125000 53.210000 68.325000 ;
        RECT 53.010000 68.535000 53.210000 68.735000 ;
        RECT 53.010000 68.945000 53.210000 69.145000 ;
        RECT 53.010000 69.355000 53.210000 69.555000 ;
        RECT 53.010000 69.765000 53.210000 69.965000 ;
        RECT 53.010000 70.175000 53.210000 70.375000 ;
        RECT 53.010000 70.585000 53.210000 70.785000 ;
        RECT 53.010000 70.995000 53.210000 71.195000 ;
        RECT 53.010000 71.405000 53.210000 71.605000 ;
        RECT 53.010000 71.815000 53.210000 72.015000 ;
        RECT 53.010000 72.225000 53.210000 72.425000 ;
        RECT 53.010000 72.635000 53.210000 72.835000 ;
        RECT 53.010000 73.045000 53.210000 73.245000 ;
        RECT 53.010000 73.450000 53.210000 73.650000 ;
        RECT 53.010000 73.855000 53.210000 74.055000 ;
        RECT 53.010000 74.260000 53.210000 74.460000 ;
        RECT 53.010000 74.665000 53.210000 74.865000 ;
        RECT 53.010000 75.070000 53.210000 75.270000 ;
        RECT 53.010000 75.475000 53.210000 75.675000 ;
        RECT 53.010000 75.880000 53.210000 76.080000 ;
        RECT 53.010000 76.285000 53.210000 76.485000 ;
        RECT 53.010000 76.690000 53.210000 76.890000 ;
        RECT 53.010000 77.095000 53.210000 77.295000 ;
        RECT 53.010000 77.500000 53.210000 77.700000 ;
        RECT 53.010000 77.905000 53.210000 78.105000 ;
        RECT 53.010000 78.310000 53.210000 78.510000 ;
        RECT 53.010000 78.715000 53.210000 78.915000 ;
        RECT 53.010000 79.120000 53.210000 79.320000 ;
        RECT 53.010000 79.525000 53.210000 79.725000 ;
        RECT 53.010000 79.930000 53.210000 80.130000 ;
        RECT 53.010000 80.335000 53.210000 80.535000 ;
        RECT 53.010000 80.740000 53.210000 80.940000 ;
        RECT 53.010000 81.145000 53.210000 81.345000 ;
        RECT 53.010000 81.550000 53.210000 81.750000 ;
        RECT 53.010000 81.955000 53.210000 82.155000 ;
        RECT 53.010000 82.360000 53.210000 82.560000 ;
        RECT 53.275000 17.860000 53.475000 18.060000 ;
        RECT 53.275000 18.290000 53.475000 18.490000 ;
        RECT 53.275000 18.720000 53.475000 18.920000 ;
        RECT 53.275000 19.150000 53.475000 19.350000 ;
        RECT 53.275000 19.580000 53.475000 19.780000 ;
        RECT 53.275000 20.010000 53.475000 20.210000 ;
        RECT 53.275000 20.440000 53.475000 20.640000 ;
        RECT 53.275000 20.870000 53.475000 21.070000 ;
        RECT 53.275000 21.300000 53.475000 21.500000 ;
        RECT 53.275000 21.730000 53.475000 21.930000 ;
        RECT 53.275000 22.160000 53.475000 22.360000 ;
        RECT 53.340000 82.920000 53.540000 83.120000 ;
        RECT 53.340000 83.470000 53.540000 83.670000 ;
        RECT 53.340000 84.020000 53.540000 84.220000 ;
        RECT 53.410000 68.125000 53.610000 68.325000 ;
        RECT 53.410000 68.535000 53.610000 68.735000 ;
        RECT 53.410000 68.945000 53.610000 69.145000 ;
        RECT 53.410000 69.355000 53.610000 69.555000 ;
        RECT 53.410000 69.765000 53.610000 69.965000 ;
        RECT 53.410000 70.175000 53.610000 70.375000 ;
        RECT 53.410000 70.585000 53.610000 70.785000 ;
        RECT 53.410000 70.995000 53.610000 71.195000 ;
        RECT 53.410000 71.405000 53.610000 71.605000 ;
        RECT 53.410000 71.815000 53.610000 72.015000 ;
        RECT 53.410000 72.225000 53.610000 72.425000 ;
        RECT 53.410000 72.635000 53.610000 72.835000 ;
        RECT 53.410000 73.045000 53.610000 73.245000 ;
        RECT 53.410000 73.450000 53.610000 73.650000 ;
        RECT 53.410000 73.855000 53.610000 74.055000 ;
        RECT 53.410000 74.260000 53.610000 74.460000 ;
        RECT 53.410000 74.665000 53.610000 74.865000 ;
        RECT 53.410000 75.070000 53.610000 75.270000 ;
        RECT 53.410000 75.475000 53.610000 75.675000 ;
        RECT 53.410000 75.880000 53.610000 76.080000 ;
        RECT 53.410000 76.285000 53.610000 76.485000 ;
        RECT 53.410000 76.690000 53.610000 76.890000 ;
        RECT 53.410000 77.095000 53.610000 77.295000 ;
        RECT 53.410000 77.500000 53.610000 77.700000 ;
        RECT 53.410000 77.905000 53.610000 78.105000 ;
        RECT 53.410000 78.310000 53.610000 78.510000 ;
        RECT 53.410000 78.715000 53.610000 78.915000 ;
        RECT 53.410000 79.120000 53.610000 79.320000 ;
        RECT 53.410000 79.525000 53.610000 79.725000 ;
        RECT 53.410000 79.930000 53.610000 80.130000 ;
        RECT 53.410000 80.335000 53.610000 80.535000 ;
        RECT 53.410000 80.740000 53.610000 80.940000 ;
        RECT 53.410000 81.145000 53.610000 81.345000 ;
        RECT 53.410000 81.550000 53.610000 81.750000 ;
        RECT 53.410000 81.955000 53.610000 82.155000 ;
        RECT 53.410000 82.360000 53.610000 82.560000 ;
        RECT 53.680000 17.860000 53.880000 18.060000 ;
        RECT 53.680000 18.290000 53.880000 18.490000 ;
        RECT 53.680000 18.720000 53.880000 18.920000 ;
        RECT 53.680000 19.150000 53.880000 19.350000 ;
        RECT 53.680000 19.580000 53.880000 19.780000 ;
        RECT 53.680000 20.010000 53.880000 20.210000 ;
        RECT 53.680000 20.440000 53.880000 20.640000 ;
        RECT 53.680000 20.870000 53.880000 21.070000 ;
        RECT 53.680000 21.300000 53.880000 21.500000 ;
        RECT 53.680000 21.730000 53.880000 21.930000 ;
        RECT 53.680000 22.160000 53.880000 22.360000 ;
        RECT 53.810000 68.125000 54.010000 68.325000 ;
        RECT 53.810000 68.535000 54.010000 68.735000 ;
        RECT 53.810000 68.945000 54.010000 69.145000 ;
        RECT 53.810000 69.355000 54.010000 69.555000 ;
        RECT 53.810000 69.765000 54.010000 69.965000 ;
        RECT 53.810000 70.175000 54.010000 70.375000 ;
        RECT 53.810000 70.585000 54.010000 70.785000 ;
        RECT 53.810000 70.995000 54.010000 71.195000 ;
        RECT 53.810000 71.405000 54.010000 71.605000 ;
        RECT 53.810000 71.815000 54.010000 72.015000 ;
        RECT 53.810000 72.225000 54.010000 72.425000 ;
        RECT 53.810000 72.635000 54.010000 72.835000 ;
        RECT 53.810000 73.045000 54.010000 73.245000 ;
        RECT 53.810000 73.450000 54.010000 73.650000 ;
        RECT 53.810000 73.855000 54.010000 74.055000 ;
        RECT 53.810000 74.260000 54.010000 74.460000 ;
        RECT 53.810000 74.665000 54.010000 74.865000 ;
        RECT 53.810000 75.070000 54.010000 75.270000 ;
        RECT 53.810000 75.475000 54.010000 75.675000 ;
        RECT 53.810000 75.880000 54.010000 76.080000 ;
        RECT 53.810000 76.285000 54.010000 76.485000 ;
        RECT 53.810000 76.690000 54.010000 76.890000 ;
        RECT 53.810000 77.095000 54.010000 77.295000 ;
        RECT 53.810000 77.500000 54.010000 77.700000 ;
        RECT 53.810000 77.905000 54.010000 78.105000 ;
        RECT 53.810000 78.310000 54.010000 78.510000 ;
        RECT 53.810000 78.715000 54.010000 78.915000 ;
        RECT 53.810000 79.120000 54.010000 79.320000 ;
        RECT 53.810000 79.525000 54.010000 79.725000 ;
        RECT 53.810000 79.930000 54.010000 80.130000 ;
        RECT 53.810000 80.335000 54.010000 80.535000 ;
        RECT 53.810000 80.740000 54.010000 80.940000 ;
        RECT 53.810000 81.145000 54.010000 81.345000 ;
        RECT 53.810000 81.550000 54.010000 81.750000 ;
        RECT 53.810000 81.955000 54.010000 82.155000 ;
        RECT 53.810000 82.360000 54.010000 82.560000 ;
        RECT 53.885000 83.010000 54.085000 83.210000 ;
        RECT 53.885000 83.470000 54.085000 83.670000 ;
        RECT 53.885000 83.930000 54.085000 84.130000 ;
        RECT 53.885000 84.395000 54.085000 84.595000 ;
        RECT 53.885000 84.860000 54.085000 85.060000 ;
        RECT 53.885000 85.325000 54.085000 85.525000 ;
        RECT 54.085000 17.860000 54.285000 18.060000 ;
        RECT 54.085000 18.290000 54.285000 18.490000 ;
        RECT 54.085000 18.720000 54.285000 18.920000 ;
        RECT 54.085000 19.150000 54.285000 19.350000 ;
        RECT 54.085000 19.580000 54.285000 19.780000 ;
        RECT 54.085000 20.010000 54.285000 20.210000 ;
        RECT 54.085000 20.440000 54.285000 20.640000 ;
        RECT 54.085000 20.870000 54.285000 21.070000 ;
        RECT 54.085000 21.300000 54.285000 21.500000 ;
        RECT 54.085000 21.730000 54.285000 21.930000 ;
        RECT 54.085000 22.160000 54.285000 22.360000 ;
        RECT 54.210000 68.125000 54.410000 68.325000 ;
        RECT 54.210000 68.535000 54.410000 68.735000 ;
        RECT 54.210000 68.945000 54.410000 69.145000 ;
        RECT 54.210000 69.355000 54.410000 69.555000 ;
        RECT 54.210000 69.765000 54.410000 69.965000 ;
        RECT 54.210000 70.175000 54.410000 70.375000 ;
        RECT 54.210000 70.585000 54.410000 70.785000 ;
        RECT 54.210000 70.995000 54.410000 71.195000 ;
        RECT 54.210000 71.405000 54.410000 71.605000 ;
        RECT 54.210000 71.815000 54.410000 72.015000 ;
        RECT 54.210000 72.225000 54.410000 72.425000 ;
        RECT 54.210000 72.635000 54.410000 72.835000 ;
        RECT 54.210000 73.045000 54.410000 73.245000 ;
        RECT 54.210000 73.450000 54.410000 73.650000 ;
        RECT 54.210000 73.855000 54.410000 74.055000 ;
        RECT 54.210000 74.260000 54.410000 74.460000 ;
        RECT 54.210000 74.665000 54.410000 74.865000 ;
        RECT 54.210000 75.070000 54.410000 75.270000 ;
        RECT 54.210000 75.475000 54.410000 75.675000 ;
        RECT 54.210000 75.880000 54.410000 76.080000 ;
        RECT 54.210000 76.285000 54.410000 76.485000 ;
        RECT 54.210000 76.690000 54.410000 76.890000 ;
        RECT 54.210000 77.095000 54.410000 77.295000 ;
        RECT 54.210000 77.500000 54.410000 77.700000 ;
        RECT 54.210000 77.905000 54.410000 78.105000 ;
        RECT 54.210000 78.310000 54.410000 78.510000 ;
        RECT 54.210000 78.715000 54.410000 78.915000 ;
        RECT 54.210000 79.120000 54.410000 79.320000 ;
        RECT 54.210000 79.525000 54.410000 79.725000 ;
        RECT 54.210000 79.930000 54.410000 80.130000 ;
        RECT 54.210000 80.335000 54.410000 80.535000 ;
        RECT 54.210000 80.740000 54.410000 80.940000 ;
        RECT 54.210000 81.145000 54.410000 81.345000 ;
        RECT 54.210000 81.550000 54.410000 81.750000 ;
        RECT 54.210000 81.955000 54.410000 82.155000 ;
        RECT 54.210000 82.360000 54.410000 82.560000 ;
        RECT 54.365000 83.010000 54.565000 83.210000 ;
        RECT 54.365000 83.470000 54.565000 83.670000 ;
        RECT 54.365000 83.930000 54.565000 84.130000 ;
        RECT 54.365000 84.395000 54.565000 84.595000 ;
        RECT 54.365000 84.860000 54.565000 85.060000 ;
        RECT 54.365000 85.325000 54.565000 85.525000 ;
        RECT 54.490000 17.860000 54.690000 18.060000 ;
        RECT 54.490000 18.290000 54.690000 18.490000 ;
        RECT 54.490000 18.720000 54.690000 18.920000 ;
        RECT 54.490000 19.150000 54.690000 19.350000 ;
        RECT 54.490000 19.580000 54.690000 19.780000 ;
        RECT 54.490000 20.010000 54.690000 20.210000 ;
        RECT 54.490000 20.440000 54.690000 20.640000 ;
        RECT 54.490000 20.870000 54.690000 21.070000 ;
        RECT 54.490000 21.300000 54.690000 21.500000 ;
        RECT 54.490000 21.730000 54.690000 21.930000 ;
        RECT 54.490000 22.160000 54.690000 22.360000 ;
        RECT 54.610000 68.125000 54.810000 68.325000 ;
        RECT 54.610000 68.535000 54.810000 68.735000 ;
        RECT 54.610000 68.945000 54.810000 69.145000 ;
        RECT 54.610000 69.355000 54.810000 69.555000 ;
        RECT 54.610000 69.765000 54.810000 69.965000 ;
        RECT 54.610000 70.175000 54.810000 70.375000 ;
        RECT 54.610000 70.585000 54.810000 70.785000 ;
        RECT 54.610000 70.995000 54.810000 71.195000 ;
        RECT 54.610000 71.405000 54.810000 71.605000 ;
        RECT 54.610000 71.815000 54.810000 72.015000 ;
        RECT 54.610000 72.225000 54.810000 72.425000 ;
        RECT 54.610000 72.635000 54.810000 72.835000 ;
        RECT 54.610000 73.045000 54.810000 73.245000 ;
        RECT 54.610000 73.450000 54.810000 73.650000 ;
        RECT 54.610000 73.855000 54.810000 74.055000 ;
        RECT 54.610000 74.260000 54.810000 74.460000 ;
        RECT 54.610000 74.665000 54.810000 74.865000 ;
        RECT 54.610000 75.070000 54.810000 75.270000 ;
        RECT 54.610000 75.475000 54.810000 75.675000 ;
        RECT 54.610000 75.880000 54.810000 76.080000 ;
        RECT 54.610000 76.285000 54.810000 76.485000 ;
        RECT 54.610000 76.690000 54.810000 76.890000 ;
        RECT 54.610000 77.095000 54.810000 77.295000 ;
        RECT 54.610000 77.500000 54.810000 77.700000 ;
        RECT 54.610000 77.905000 54.810000 78.105000 ;
        RECT 54.610000 78.310000 54.810000 78.510000 ;
        RECT 54.610000 78.715000 54.810000 78.915000 ;
        RECT 54.610000 79.120000 54.810000 79.320000 ;
        RECT 54.610000 79.525000 54.810000 79.725000 ;
        RECT 54.610000 79.930000 54.810000 80.130000 ;
        RECT 54.610000 80.335000 54.810000 80.535000 ;
        RECT 54.610000 80.740000 54.810000 80.940000 ;
        RECT 54.610000 81.145000 54.810000 81.345000 ;
        RECT 54.610000 81.550000 54.810000 81.750000 ;
        RECT 54.610000 81.955000 54.810000 82.155000 ;
        RECT 54.610000 82.360000 54.810000 82.560000 ;
        RECT 54.845000 83.010000 55.045000 83.210000 ;
        RECT 54.845000 83.470000 55.045000 83.670000 ;
        RECT 54.845000 83.930000 55.045000 84.130000 ;
        RECT 54.845000 84.395000 55.045000 84.595000 ;
        RECT 54.845000 84.860000 55.045000 85.060000 ;
        RECT 54.845000 85.325000 55.045000 85.525000 ;
        RECT 54.895000 17.860000 55.095000 18.060000 ;
        RECT 54.895000 18.290000 55.095000 18.490000 ;
        RECT 54.895000 18.720000 55.095000 18.920000 ;
        RECT 54.895000 19.150000 55.095000 19.350000 ;
        RECT 54.895000 19.580000 55.095000 19.780000 ;
        RECT 54.895000 20.010000 55.095000 20.210000 ;
        RECT 54.895000 20.440000 55.095000 20.640000 ;
        RECT 54.895000 20.870000 55.095000 21.070000 ;
        RECT 54.895000 21.300000 55.095000 21.500000 ;
        RECT 54.895000 21.730000 55.095000 21.930000 ;
        RECT 54.895000 22.160000 55.095000 22.360000 ;
        RECT 55.010000 68.125000 55.210000 68.325000 ;
        RECT 55.010000 68.535000 55.210000 68.735000 ;
        RECT 55.010000 68.945000 55.210000 69.145000 ;
        RECT 55.010000 69.355000 55.210000 69.555000 ;
        RECT 55.010000 69.765000 55.210000 69.965000 ;
        RECT 55.010000 70.175000 55.210000 70.375000 ;
        RECT 55.010000 70.585000 55.210000 70.785000 ;
        RECT 55.010000 70.995000 55.210000 71.195000 ;
        RECT 55.010000 71.405000 55.210000 71.605000 ;
        RECT 55.010000 71.815000 55.210000 72.015000 ;
        RECT 55.010000 72.225000 55.210000 72.425000 ;
        RECT 55.010000 72.635000 55.210000 72.835000 ;
        RECT 55.010000 73.045000 55.210000 73.245000 ;
        RECT 55.010000 73.450000 55.210000 73.650000 ;
        RECT 55.010000 73.855000 55.210000 74.055000 ;
        RECT 55.010000 74.260000 55.210000 74.460000 ;
        RECT 55.010000 74.665000 55.210000 74.865000 ;
        RECT 55.010000 75.070000 55.210000 75.270000 ;
        RECT 55.010000 75.475000 55.210000 75.675000 ;
        RECT 55.010000 75.880000 55.210000 76.080000 ;
        RECT 55.010000 76.285000 55.210000 76.485000 ;
        RECT 55.010000 76.690000 55.210000 76.890000 ;
        RECT 55.010000 77.095000 55.210000 77.295000 ;
        RECT 55.010000 77.500000 55.210000 77.700000 ;
        RECT 55.010000 77.905000 55.210000 78.105000 ;
        RECT 55.010000 78.310000 55.210000 78.510000 ;
        RECT 55.010000 78.715000 55.210000 78.915000 ;
        RECT 55.010000 79.120000 55.210000 79.320000 ;
        RECT 55.010000 79.525000 55.210000 79.725000 ;
        RECT 55.010000 79.930000 55.210000 80.130000 ;
        RECT 55.010000 80.335000 55.210000 80.535000 ;
        RECT 55.010000 80.740000 55.210000 80.940000 ;
        RECT 55.010000 81.145000 55.210000 81.345000 ;
        RECT 55.010000 81.550000 55.210000 81.750000 ;
        RECT 55.010000 81.955000 55.210000 82.155000 ;
        RECT 55.010000 82.360000 55.210000 82.560000 ;
        RECT 55.255000 85.875000 55.455000 86.075000 ;
        RECT 55.255000 86.310000 55.455000 86.510000 ;
        RECT 55.255000 86.750000 55.455000 86.950000 ;
        RECT 55.300000 17.860000 55.500000 18.060000 ;
        RECT 55.300000 18.290000 55.500000 18.490000 ;
        RECT 55.300000 18.720000 55.500000 18.920000 ;
        RECT 55.300000 19.150000 55.500000 19.350000 ;
        RECT 55.300000 19.580000 55.500000 19.780000 ;
        RECT 55.300000 20.010000 55.500000 20.210000 ;
        RECT 55.300000 20.440000 55.500000 20.640000 ;
        RECT 55.300000 20.870000 55.500000 21.070000 ;
        RECT 55.300000 21.300000 55.500000 21.500000 ;
        RECT 55.300000 21.730000 55.500000 21.930000 ;
        RECT 55.300000 22.160000 55.500000 22.360000 ;
        RECT 55.325000 83.010000 55.525000 83.210000 ;
        RECT 55.325000 83.470000 55.525000 83.670000 ;
        RECT 55.325000 83.930000 55.525000 84.130000 ;
        RECT 55.325000 84.395000 55.525000 84.595000 ;
        RECT 55.325000 84.860000 55.525000 85.060000 ;
        RECT 55.325000 85.325000 55.525000 85.525000 ;
        RECT 55.410000 68.125000 55.610000 68.325000 ;
        RECT 55.410000 68.535000 55.610000 68.735000 ;
        RECT 55.410000 68.945000 55.610000 69.145000 ;
        RECT 55.410000 69.355000 55.610000 69.555000 ;
        RECT 55.410000 69.765000 55.610000 69.965000 ;
        RECT 55.410000 70.175000 55.610000 70.375000 ;
        RECT 55.410000 70.585000 55.610000 70.785000 ;
        RECT 55.410000 70.995000 55.610000 71.195000 ;
        RECT 55.410000 71.405000 55.610000 71.605000 ;
        RECT 55.410000 71.815000 55.610000 72.015000 ;
        RECT 55.410000 72.225000 55.610000 72.425000 ;
        RECT 55.410000 72.635000 55.610000 72.835000 ;
        RECT 55.410000 73.045000 55.610000 73.245000 ;
        RECT 55.410000 73.450000 55.610000 73.650000 ;
        RECT 55.410000 73.855000 55.610000 74.055000 ;
        RECT 55.410000 74.260000 55.610000 74.460000 ;
        RECT 55.410000 74.665000 55.610000 74.865000 ;
        RECT 55.410000 75.070000 55.610000 75.270000 ;
        RECT 55.410000 75.475000 55.610000 75.675000 ;
        RECT 55.410000 75.880000 55.610000 76.080000 ;
        RECT 55.410000 76.285000 55.610000 76.485000 ;
        RECT 55.410000 76.690000 55.610000 76.890000 ;
        RECT 55.410000 77.095000 55.610000 77.295000 ;
        RECT 55.410000 77.500000 55.610000 77.700000 ;
        RECT 55.410000 77.905000 55.610000 78.105000 ;
        RECT 55.410000 78.310000 55.610000 78.510000 ;
        RECT 55.410000 78.715000 55.610000 78.915000 ;
        RECT 55.410000 79.120000 55.610000 79.320000 ;
        RECT 55.410000 79.525000 55.610000 79.725000 ;
        RECT 55.410000 79.930000 55.610000 80.130000 ;
        RECT 55.410000 80.335000 55.610000 80.535000 ;
        RECT 55.410000 80.740000 55.610000 80.940000 ;
        RECT 55.410000 81.145000 55.610000 81.345000 ;
        RECT 55.410000 81.550000 55.610000 81.750000 ;
        RECT 55.410000 81.955000 55.610000 82.155000 ;
        RECT 55.410000 82.360000 55.610000 82.560000 ;
        RECT 55.705000 17.860000 55.905000 18.060000 ;
        RECT 55.705000 18.290000 55.905000 18.490000 ;
        RECT 55.705000 18.720000 55.905000 18.920000 ;
        RECT 55.705000 19.150000 55.905000 19.350000 ;
        RECT 55.705000 19.580000 55.905000 19.780000 ;
        RECT 55.705000 20.010000 55.905000 20.210000 ;
        RECT 55.705000 20.440000 55.905000 20.640000 ;
        RECT 55.705000 20.870000 55.905000 21.070000 ;
        RECT 55.705000 21.300000 55.905000 21.500000 ;
        RECT 55.705000 21.730000 55.905000 21.930000 ;
        RECT 55.705000 22.160000 55.905000 22.360000 ;
        RECT 55.805000 83.010000 56.005000 83.210000 ;
        RECT 55.805000 83.470000 56.005000 83.670000 ;
        RECT 55.805000 83.930000 56.005000 84.130000 ;
        RECT 55.805000 84.395000 56.005000 84.595000 ;
        RECT 55.805000 84.860000 56.005000 85.060000 ;
        RECT 55.805000 85.325000 56.005000 85.525000 ;
        RECT 55.810000 68.125000 56.010000 68.325000 ;
        RECT 55.810000 68.535000 56.010000 68.735000 ;
        RECT 55.810000 68.945000 56.010000 69.145000 ;
        RECT 55.810000 69.355000 56.010000 69.555000 ;
        RECT 55.810000 69.765000 56.010000 69.965000 ;
        RECT 55.810000 70.175000 56.010000 70.375000 ;
        RECT 55.810000 70.585000 56.010000 70.785000 ;
        RECT 55.810000 70.995000 56.010000 71.195000 ;
        RECT 55.810000 71.405000 56.010000 71.605000 ;
        RECT 55.810000 71.815000 56.010000 72.015000 ;
        RECT 55.810000 72.225000 56.010000 72.425000 ;
        RECT 55.810000 72.635000 56.010000 72.835000 ;
        RECT 55.810000 73.045000 56.010000 73.245000 ;
        RECT 55.810000 73.450000 56.010000 73.650000 ;
        RECT 55.810000 73.855000 56.010000 74.055000 ;
        RECT 55.810000 74.260000 56.010000 74.460000 ;
        RECT 55.810000 74.665000 56.010000 74.865000 ;
        RECT 55.810000 75.070000 56.010000 75.270000 ;
        RECT 55.810000 75.475000 56.010000 75.675000 ;
        RECT 55.810000 75.880000 56.010000 76.080000 ;
        RECT 55.810000 76.285000 56.010000 76.485000 ;
        RECT 55.810000 76.690000 56.010000 76.890000 ;
        RECT 55.810000 77.095000 56.010000 77.295000 ;
        RECT 55.810000 77.500000 56.010000 77.700000 ;
        RECT 55.810000 77.905000 56.010000 78.105000 ;
        RECT 55.810000 78.310000 56.010000 78.510000 ;
        RECT 55.810000 78.715000 56.010000 78.915000 ;
        RECT 55.810000 79.120000 56.010000 79.320000 ;
        RECT 55.810000 79.525000 56.010000 79.725000 ;
        RECT 55.810000 79.930000 56.010000 80.130000 ;
        RECT 55.810000 80.335000 56.010000 80.535000 ;
        RECT 55.810000 80.740000 56.010000 80.940000 ;
        RECT 55.810000 81.145000 56.010000 81.345000 ;
        RECT 55.810000 81.550000 56.010000 81.750000 ;
        RECT 55.810000 81.955000 56.010000 82.155000 ;
        RECT 55.810000 82.360000 56.010000 82.560000 ;
        RECT 55.995000 85.875000 56.195000 86.075000 ;
        RECT 55.995000 86.310000 56.195000 86.510000 ;
        RECT 55.995000 86.750000 56.195000 86.950000 ;
        RECT 56.110000 17.860000 56.310000 18.060000 ;
        RECT 56.110000 18.290000 56.310000 18.490000 ;
        RECT 56.110000 18.720000 56.310000 18.920000 ;
        RECT 56.110000 19.150000 56.310000 19.350000 ;
        RECT 56.110000 19.580000 56.310000 19.780000 ;
        RECT 56.110000 20.010000 56.310000 20.210000 ;
        RECT 56.110000 20.440000 56.310000 20.640000 ;
        RECT 56.110000 20.870000 56.310000 21.070000 ;
        RECT 56.110000 21.300000 56.310000 21.500000 ;
        RECT 56.110000 21.730000 56.310000 21.930000 ;
        RECT 56.110000 22.160000 56.310000 22.360000 ;
        RECT 56.210000 68.125000 56.410000 68.325000 ;
        RECT 56.210000 68.535000 56.410000 68.735000 ;
        RECT 56.210000 68.945000 56.410000 69.145000 ;
        RECT 56.210000 69.355000 56.410000 69.555000 ;
        RECT 56.210000 69.765000 56.410000 69.965000 ;
        RECT 56.210000 70.175000 56.410000 70.375000 ;
        RECT 56.210000 70.585000 56.410000 70.785000 ;
        RECT 56.210000 70.995000 56.410000 71.195000 ;
        RECT 56.210000 71.405000 56.410000 71.605000 ;
        RECT 56.210000 71.815000 56.410000 72.015000 ;
        RECT 56.210000 72.225000 56.410000 72.425000 ;
        RECT 56.210000 72.635000 56.410000 72.835000 ;
        RECT 56.210000 73.045000 56.410000 73.245000 ;
        RECT 56.210000 73.450000 56.410000 73.650000 ;
        RECT 56.210000 73.855000 56.410000 74.055000 ;
        RECT 56.210000 74.260000 56.410000 74.460000 ;
        RECT 56.210000 74.665000 56.410000 74.865000 ;
        RECT 56.210000 75.070000 56.410000 75.270000 ;
        RECT 56.210000 75.475000 56.410000 75.675000 ;
        RECT 56.210000 75.880000 56.410000 76.080000 ;
        RECT 56.210000 76.285000 56.410000 76.485000 ;
        RECT 56.210000 76.690000 56.410000 76.890000 ;
        RECT 56.210000 77.095000 56.410000 77.295000 ;
        RECT 56.210000 77.500000 56.410000 77.700000 ;
        RECT 56.210000 77.905000 56.410000 78.105000 ;
        RECT 56.210000 78.310000 56.410000 78.510000 ;
        RECT 56.210000 78.715000 56.410000 78.915000 ;
        RECT 56.210000 79.120000 56.410000 79.320000 ;
        RECT 56.210000 79.525000 56.410000 79.725000 ;
        RECT 56.210000 79.930000 56.410000 80.130000 ;
        RECT 56.210000 80.335000 56.410000 80.535000 ;
        RECT 56.210000 80.740000 56.410000 80.940000 ;
        RECT 56.210000 81.145000 56.410000 81.345000 ;
        RECT 56.210000 81.550000 56.410000 81.750000 ;
        RECT 56.210000 81.955000 56.410000 82.155000 ;
        RECT 56.210000 82.360000 56.410000 82.560000 ;
        RECT 56.490000 83.055000 56.690000 83.255000 ;
        RECT 56.490000 83.455000 56.690000 83.655000 ;
        RECT 56.490000 83.855000 56.690000 84.055000 ;
        RECT 56.490000 84.255000 56.690000 84.455000 ;
        RECT 56.490000 84.655000 56.690000 84.855000 ;
        RECT 56.490000 85.055000 56.690000 85.255000 ;
        RECT 56.490000 85.455000 56.690000 85.655000 ;
        RECT 56.490000 85.855000 56.690000 86.055000 ;
        RECT 56.490000 86.255000 56.690000 86.455000 ;
        RECT 56.490000 86.660000 56.690000 86.860000 ;
        RECT 56.490000 87.065000 56.690000 87.265000 ;
        RECT 56.490000 87.470000 56.690000 87.670000 ;
        RECT 56.490000 87.875000 56.690000 88.075000 ;
        RECT 56.515000 17.860000 56.715000 18.060000 ;
        RECT 56.515000 18.290000 56.715000 18.490000 ;
        RECT 56.515000 18.720000 56.715000 18.920000 ;
        RECT 56.515000 19.150000 56.715000 19.350000 ;
        RECT 56.515000 19.580000 56.715000 19.780000 ;
        RECT 56.515000 20.010000 56.715000 20.210000 ;
        RECT 56.515000 20.440000 56.715000 20.640000 ;
        RECT 56.515000 20.870000 56.715000 21.070000 ;
        RECT 56.515000 21.300000 56.715000 21.500000 ;
        RECT 56.515000 21.730000 56.715000 21.930000 ;
        RECT 56.515000 22.160000 56.715000 22.360000 ;
        RECT 56.610000 68.125000 56.810000 68.325000 ;
        RECT 56.610000 68.535000 56.810000 68.735000 ;
        RECT 56.610000 68.945000 56.810000 69.145000 ;
        RECT 56.610000 69.355000 56.810000 69.555000 ;
        RECT 56.610000 69.765000 56.810000 69.965000 ;
        RECT 56.610000 70.175000 56.810000 70.375000 ;
        RECT 56.610000 70.585000 56.810000 70.785000 ;
        RECT 56.610000 70.995000 56.810000 71.195000 ;
        RECT 56.610000 71.405000 56.810000 71.605000 ;
        RECT 56.610000 71.815000 56.810000 72.015000 ;
        RECT 56.610000 72.225000 56.810000 72.425000 ;
        RECT 56.610000 72.635000 56.810000 72.835000 ;
        RECT 56.610000 73.045000 56.810000 73.245000 ;
        RECT 56.610000 73.450000 56.810000 73.650000 ;
        RECT 56.610000 73.855000 56.810000 74.055000 ;
        RECT 56.610000 74.260000 56.810000 74.460000 ;
        RECT 56.610000 74.665000 56.810000 74.865000 ;
        RECT 56.610000 75.070000 56.810000 75.270000 ;
        RECT 56.610000 75.475000 56.810000 75.675000 ;
        RECT 56.610000 75.880000 56.810000 76.080000 ;
        RECT 56.610000 76.285000 56.810000 76.485000 ;
        RECT 56.610000 76.690000 56.810000 76.890000 ;
        RECT 56.610000 77.095000 56.810000 77.295000 ;
        RECT 56.610000 77.500000 56.810000 77.700000 ;
        RECT 56.610000 77.905000 56.810000 78.105000 ;
        RECT 56.610000 78.310000 56.810000 78.510000 ;
        RECT 56.610000 78.715000 56.810000 78.915000 ;
        RECT 56.610000 79.120000 56.810000 79.320000 ;
        RECT 56.610000 79.525000 56.810000 79.725000 ;
        RECT 56.610000 79.930000 56.810000 80.130000 ;
        RECT 56.610000 80.335000 56.810000 80.535000 ;
        RECT 56.610000 80.740000 56.810000 80.940000 ;
        RECT 56.610000 81.145000 56.810000 81.345000 ;
        RECT 56.610000 81.550000 56.810000 81.750000 ;
        RECT 56.610000 81.955000 56.810000 82.155000 ;
        RECT 56.610000 82.360000 56.810000 82.560000 ;
        RECT 56.900000 83.055000 57.100000 83.255000 ;
        RECT 56.900000 83.455000 57.100000 83.655000 ;
        RECT 56.900000 83.855000 57.100000 84.055000 ;
        RECT 56.900000 84.255000 57.100000 84.455000 ;
        RECT 56.900000 84.655000 57.100000 84.855000 ;
        RECT 56.900000 85.055000 57.100000 85.255000 ;
        RECT 56.900000 85.455000 57.100000 85.655000 ;
        RECT 56.900000 85.855000 57.100000 86.055000 ;
        RECT 56.900000 86.255000 57.100000 86.455000 ;
        RECT 56.900000 86.660000 57.100000 86.860000 ;
        RECT 56.900000 87.065000 57.100000 87.265000 ;
        RECT 56.900000 87.470000 57.100000 87.670000 ;
        RECT 56.900000 87.875000 57.100000 88.075000 ;
        RECT 56.920000 17.860000 57.120000 18.060000 ;
        RECT 56.920000 18.290000 57.120000 18.490000 ;
        RECT 56.920000 18.720000 57.120000 18.920000 ;
        RECT 56.920000 19.150000 57.120000 19.350000 ;
        RECT 56.920000 19.580000 57.120000 19.780000 ;
        RECT 56.920000 20.010000 57.120000 20.210000 ;
        RECT 56.920000 20.440000 57.120000 20.640000 ;
        RECT 56.920000 20.870000 57.120000 21.070000 ;
        RECT 56.920000 21.300000 57.120000 21.500000 ;
        RECT 56.920000 21.730000 57.120000 21.930000 ;
        RECT 56.920000 22.160000 57.120000 22.360000 ;
        RECT 57.010000 68.125000 57.210000 68.325000 ;
        RECT 57.010000 68.535000 57.210000 68.735000 ;
        RECT 57.010000 68.945000 57.210000 69.145000 ;
        RECT 57.010000 69.355000 57.210000 69.555000 ;
        RECT 57.010000 69.765000 57.210000 69.965000 ;
        RECT 57.010000 70.175000 57.210000 70.375000 ;
        RECT 57.010000 70.585000 57.210000 70.785000 ;
        RECT 57.010000 70.995000 57.210000 71.195000 ;
        RECT 57.010000 71.405000 57.210000 71.605000 ;
        RECT 57.010000 71.815000 57.210000 72.015000 ;
        RECT 57.010000 72.225000 57.210000 72.425000 ;
        RECT 57.010000 72.635000 57.210000 72.835000 ;
        RECT 57.010000 73.045000 57.210000 73.245000 ;
        RECT 57.010000 73.450000 57.210000 73.650000 ;
        RECT 57.010000 73.855000 57.210000 74.055000 ;
        RECT 57.010000 74.260000 57.210000 74.460000 ;
        RECT 57.010000 74.665000 57.210000 74.865000 ;
        RECT 57.010000 75.070000 57.210000 75.270000 ;
        RECT 57.010000 75.475000 57.210000 75.675000 ;
        RECT 57.010000 75.880000 57.210000 76.080000 ;
        RECT 57.010000 76.285000 57.210000 76.485000 ;
        RECT 57.010000 76.690000 57.210000 76.890000 ;
        RECT 57.010000 77.095000 57.210000 77.295000 ;
        RECT 57.010000 77.500000 57.210000 77.700000 ;
        RECT 57.010000 77.905000 57.210000 78.105000 ;
        RECT 57.010000 78.310000 57.210000 78.510000 ;
        RECT 57.010000 78.715000 57.210000 78.915000 ;
        RECT 57.010000 79.120000 57.210000 79.320000 ;
        RECT 57.010000 79.525000 57.210000 79.725000 ;
        RECT 57.010000 79.930000 57.210000 80.130000 ;
        RECT 57.010000 80.335000 57.210000 80.535000 ;
        RECT 57.010000 80.740000 57.210000 80.940000 ;
        RECT 57.010000 81.145000 57.210000 81.345000 ;
        RECT 57.010000 81.550000 57.210000 81.750000 ;
        RECT 57.010000 81.955000 57.210000 82.155000 ;
        RECT 57.010000 82.360000 57.210000 82.560000 ;
        RECT 57.310000 83.055000 57.510000 83.255000 ;
        RECT 57.310000 83.455000 57.510000 83.655000 ;
        RECT 57.310000 83.855000 57.510000 84.055000 ;
        RECT 57.310000 84.255000 57.510000 84.455000 ;
        RECT 57.310000 84.655000 57.510000 84.855000 ;
        RECT 57.310000 85.055000 57.510000 85.255000 ;
        RECT 57.310000 85.455000 57.510000 85.655000 ;
        RECT 57.310000 85.855000 57.510000 86.055000 ;
        RECT 57.310000 86.255000 57.510000 86.455000 ;
        RECT 57.310000 86.660000 57.510000 86.860000 ;
        RECT 57.310000 87.065000 57.510000 87.265000 ;
        RECT 57.310000 87.470000 57.510000 87.670000 ;
        RECT 57.310000 87.875000 57.510000 88.075000 ;
        RECT 57.325000 17.860000 57.525000 18.060000 ;
        RECT 57.325000 18.290000 57.525000 18.490000 ;
        RECT 57.325000 18.720000 57.525000 18.920000 ;
        RECT 57.325000 19.150000 57.525000 19.350000 ;
        RECT 57.325000 19.580000 57.525000 19.780000 ;
        RECT 57.325000 20.010000 57.525000 20.210000 ;
        RECT 57.325000 20.440000 57.525000 20.640000 ;
        RECT 57.325000 20.870000 57.525000 21.070000 ;
        RECT 57.325000 21.300000 57.525000 21.500000 ;
        RECT 57.325000 21.730000 57.525000 21.930000 ;
        RECT 57.325000 22.160000 57.525000 22.360000 ;
        RECT 57.410000 68.125000 57.610000 68.325000 ;
        RECT 57.410000 68.535000 57.610000 68.735000 ;
        RECT 57.410000 68.945000 57.610000 69.145000 ;
        RECT 57.410000 69.355000 57.610000 69.555000 ;
        RECT 57.410000 69.765000 57.610000 69.965000 ;
        RECT 57.410000 70.175000 57.610000 70.375000 ;
        RECT 57.410000 70.585000 57.610000 70.785000 ;
        RECT 57.410000 70.995000 57.610000 71.195000 ;
        RECT 57.410000 71.405000 57.610000 71.605000 ;
        RECT 57.410000 71.815000 57.610000 72.015000 ;
        RECT 57.410000 72.225000 57.610000 72.425000 ;
        RECT 57.410000 72.635000 57.610000 72.835000 ;
        RECT 57.410000 73.045000 57.610000 73.245000 ;
        RECT 57.410000 73.450000 57.610000 73.650000 ;
        RECT 57.410000 73.855000 57.610000 74.055000 ;
        RECT 57.410000 74.260000 57.610000 74.460000 ;
        RECT 57.410000 74.665000 57.610000 74.865000 ;
        RECT 57.410000 75.070000 57.610000 75.270000 ;
        RECT 57.410000 75.475000 57.610000 75.675000 ;
        RECT 57.410000 75.880000 57.610000 76.080000 ;
        RECT 57.410000 76.285000 57.610000 76.485000 ;
        RECT 57.410000 76.690000 57.610000 76.890000 ;
        RECT 57.410000 77.095000 57.610000 77.295000 ;
        RECT 57.410000 77.500000 57.610000 77.700000 ;
        RECT 57.410000 77.905000 57.610000 78.105000 ;
        RECT 57.410000 78.310000 57.610000 78.510000 ;
        RECT 57.410000 78.715000 57.610000 78.915000 ;
        RECT 57.410000 79.120000 57.610000 79.320000 ;
        RECT 57.410000 79.525000 57.610000 79.725000 ;
        RECT 57.410000 79.930000 57.610000 80.130000 ;
        RECT 57.410000 80.335000 57.610000 80.535000 ;
        RECT 57.410000 80.740000 57.610000 80.940000 ;
        RECT 57.410000 81.145000 57.610000 81.345000 ;
        RECT 57.410000 81.550000 57.610000 81.750000 ;
        RECT 57.410000 81.955000 57.610000 82.155000 ;
        RECT 57.410000 82.360000 57.610000 82.560000 ;
        RECT 57.720000 83.055000 57.920000 83.255000 ;
        RECT 57.720000 83.455000 57.920000 83.655000 ;
        RECT 57.720000 83.855000 57.920000 84.055000 ;
        RECT 57.720000 84.255000 57.920000 84.455000 ;
        RECT 57.720000 84.655000 57.920000 84.855000 ;
        RECT 57.720000 85.055000 57.920000 85.255000 ;
        RECT 57.720000 85.455000 57.920000 85.655000 ;
        RECT 57.720000 85.855000 57.920000 86.055000 ;
        RECT 57.720000 86.255000 57.920000 86.455000 ;
        RECT 57.720000 86.660000 57.920000 86.860000 ;
        RECT 57.720000 87.065000 57.920000 87.265000 ;
        RECT 57.720000 87.470000 57.920000 87.670000 ;
        RECT 57.720000 87.875000 57.920000 88.075000 ;
        RECT 57.730000 17.860000 57.930000 18.060000 ;
        RECT 57.730000 18.290000 57.930000 18.490000 ;
        RECT 57.730000 18.720000 57.930000 18.920000 ;
        RECT 57.730000 19.150000 57.930000 19.350000 ;
        RECT 57.730000 19.580000 57.930000 19.780000 ;
        RECT 57.730000 20.010000 57.930000 20.210000 ;
        RECT 57.730000 20.440000 57.930000 20.640000 ;
        RECT 57.730000 20.870000 57.930000 21.070000 ;
        RECT 57.730000 21.300000 57.930000 21.500000 ;
        RECT 57.730000 21.730000 57.930000 21.930000 ;
        RECT 57.730000 22.160000 57.930000 22.360000 ;
        RECT 57.795000 88.430000 57.995000 88.630000 ;
        RECT 57.795000 88.845000 57.995000 89.045000 ;
        RECT 57.795000 89.265000 57.995000 89.465000 ;
        RECT 57.810000 68.125000 58.010000 68.325000 ;
        RECT 57.810000 68.535000 58.010000 68.735000 ;
        RECT 57.810000 68.945000 58.010000 69.145000 ;
        RECT 57.810000 69.355000 58.010000 69.555000 ;
        RECT 57.810000 69.765000 58.010000 69.965000 ;
        RECT 57.810000 70.175000 58.010000 70.375000 ;
        RECT 57.810000 70.585000 58.010000 70.785000 ;
        RECT 57.810000 70.995000 58.010000 71.195000 ;
        RECT 57.810000 71.405000 58.010000 71.605000 ;
        RECT 57.810000 71.815000 58.010000 72.015000 ;
        RECT 57.810000 72.225000 58.010000 72.425000 ;
        RECT 57.810000 72.635000 58.010000 72.835000 ;
        RECT 57.810000 73.045000 58.010000 73.245000 ;
        RECT 57.810000 73.450000 58.010000 73.650000 ;
        RECT 57.810000 73.855000 58.010000 74.055000 ;
        RECT 57.810000 74.260000 58.010000 74.460000 ;
        RECT 57.810000 74.665000 58.010000 74.865000 ;
        RECT 57.810000 75.070000 58.010000 75.270000 ;
        RECT 57.810000 75.475000 58.010000 75.675000 ;
        RECT 57.810000 75.880000 58.010000 76.080000 ;
        RECT 57.810000 76.285000 58.010000 76.485000 ;
        RECT 57.810000 76.690000 58.010000 76.890000 ;
        RECT 57.810000 77.095000 58.010000 77.295000 ;
        RECT 57.810000 77.500000 58.010000 77.700000 ;
        RECT 57.810000 77.905000 58.010000 78.105000 ;
        RECT 57.810000 78.310000 58.010000 78.510000 ;
        RECT 57.810000 78.715000 58.010000 78.915000 ;
        RECT 57.810000 79.120000 58.010000 79.320000 ;
        RECT 57.810000 79.525000 58.010000 79.725000 ;
        RECT 57.810000 79.930000 58.010000 80.130000 ;
        RECT 57.810000 80.335000 58.010000 80.535000 ;
        RECT 57.810000 80.740000 58.010000 80.940000 ;
        RECT 57.810000 81.145000 58.010000 81.345000 ;
        RECT 57.810000 81.550000 58.010000 81.750000 ;
        RECT 57.810000 81.955000 58.010000 82.155000 ;
        RECT 57.810000 82.360000 58.010000 82.560000 ;
        RECT 58.130000 83.055000 58.330000 83.255000 ;
        RECT 58.130000 83.455000 58.330000 83.655000 ;
        RECT 58.130000 83.855000 58.330000 84.055000 ;
        RECT 58.130000 84.255000 58.330000 84.455000 ;
        RECT 58.130000 84.655000 58.330000 84.855000 ;
        RECT 58.130000 85.055000 58.330000 85.255000 ;
        RECT 58.130000 85.455000 58.330000 85.655000 ;
        RECT 58.130000 85.855000 58.330000 86.055000 ;
        RECT 58.130000 86.255000 58.330000 86.455000 ;
        RECT 58.130000 86.660000 58.330000 86.860000 ;
        RECT 58.130000 87.065000 58.330000 87.265000 ;
        RECT 58.130000 87.470000 58.330000 87.670000 ;
        RECT 58.130000 87.875000 58.330000 88.075000 ;
        RECT 58.135000 17.860000 58.335000 18.060000 ;
        RECT 58.135000 18.290000 58.335000 18.490000 ;
        RECT 58.135000 18.720000 58.335000 18.920000 ;
        RECT 58.135000 19.150000 58.335000 19.350000 ;
        RECT 58.135000 19.580000 58.335000 19.780000 ;
        RECT 58.135000 20.010000 58.335000 20.210000 ;
        RECT 58.135000 20.440000 58.335000 20.640000 ;
        RECT 58.135000 20.870000 58.335000 21.070000 ;
        RECT 58.135000 21.300000 58.335000 21.500000 ;
        RECT 58.135000 21.730000 58.335000 21.930000 ;
        RECT 58.135000 22.160000 58.335000 22.360000 ;
        RECT 58.210000 68.125000 58.410000 68.325000 ;
        RECT 58.210000 68.535000 58.410000 68.735000 ;
        RECT 58.210000 68.945000 58.410000 69.145000 ;
        RECT 58.210000 69.355000 58.410000 69.555000 ;
        RECT 58.210000 69.765000 58.410000 69.965000 ;
        RECT 58.210000 70.175000 58.410000 70.375000 ;
        RECT 58.210000 70.585000 58.410000 70.785000 ;
        RECT 58.210000 70.995000 58.410000 71.195000 ;
        RECT 58.210000 71.405000 58.410000 71.605000 ;
        RECT 58.210000 71.815000 58.410000 72.015000 ;
        RECT 58.210000 72.225000 58.410000 72.425000 ;
        RECT 58.210000 72.635000 58.410000 72.835000 ;
        RECT 58.210000 73.045000 58.410000 73.245000 ;
        RECT 58.210000 73.450000 58.410000 73.650000 ;
        RECT 58.210000 73.855000 58.410000 74.055000 ;
        RECT 58.210000 74.260000 58.410000 74.460000 ;
        RECT 58.210000 74.665000 58.410000 74.865000 ;
        RECT 58.210000 75.070000 58.410000 75.270000 ;
        RECT 58.210000 75.475000 58.410000 75.675000 ;
        RECT 58.210000 75.880000 58.410000 76.080000 ;
        RECT 58.210000 76.285000 58.410000 76.485000 ;
        RECT 58.210000 76.690000 58.410000 76.890000 ;
        RECT 58.210000 77.095000 58.410000 77.295000 ;
        RECT 58.210000 77.500000 58.410000 77.700000 ;
        RECT 58.210000 77.905000 58.410000 78.105000 ;
        RECT 58.210000 78.310000 58.410000 78.510000 ;
        RECT 58.210000 78.715000 58.410000 78.915000 ;
        RECT 58.210000 79.120000 58.410000 79.320000 ;
        RECT 58.210000 79.525000 58.410000 79.725000 ;
        RECT 58.210000 79.930000 58.410000 80.130000 ;
        RECT 58.210000 80.335000 58.410000 80.535000 ;
        RECT 58.210000 80.740000 58.410000 80.940000 ;
        RECT 58.210000 81.145000 58.410000 81.345000 ;
        RECT 58.210000 81.550000 58.410000 81.750000 ;
        RECT 58.210000 81.955000 58.410000 82.155000 ;
        RECT 58.210000 82.360000 58.410000 82.560000 ;
        RECT 58.540000 17.860000 58.740000 18.060000 ;
        RECT 58.540000 18.290000 58.740000 18.490000 ;
        RECT 58.540000 18.720000 58.740000 18.920000 ;
        RECT 58.540000 19.150000 58.740000 19.350000 ;
        RECT 58.540000 19.580000 58.740000 19.780000 ;
        RECT 58.540000 20.010000 58.740000 20.210000 ;
        RECT 58.540000 20.440000 58.740000 20.640000 ;
        RECT 58.540000 20.870000 58.740000 21.070000 ;
        RECT 58.540000 21.300000 58.740000 21.500000 ;
        RECT 58.540000 21.730000 58.740000 21.930000 ;
        RECT 58.540000 22.160000 58.740000 22.360000 ;
        RECT 58.540000 83.055000 58.740000 83.255000 ;
        RECT 58.540000 83.455000 58.740000 83.655000 ;
        RECT 58.540000 83.855000 58.740000 84.055000 ;
        RECT 58.540000 84.255000 58.740000 84.455000 ;
        RECT 58.540000 84.655000 58.740000 84.855000 ;
        RECT 58.540000 85.055000 58.740000 85.255000 ;
        RECT 58.540000 85.455000 58.740000 85.655000 ;
        RECT 58.540000 85.855000 58.740000 86.055000 ;
        RECT 58.540000 86.255000 58.740000 86.455000 ;
        RECT 58.540000 86.660000 58.740000 86.860000 ;
        RECT 58.540000 87.065000 58.740000 87.265000 ;
        RECT 58.540000 87.470000 58.740000 87.670000 ;
        RECT 58.540000 87.875000 58.740000 88.075000 ;
        RECT 58.575000 88.430000 58.775000 88.630000 ;
        RECT 58.575000 88.845000 58.775000 89.045000 ;
        RECT 58.575000 89.265000 58.775000 89.465000 ;
        RECT 58.610000 68.125000 58.810000 68.325000 ;
        RECT 58.610000 68.535000 58.810000 68.735000 ;
        RECT 58.610000 68.945000 58.810000 69.145000 ;
        RECT 58.610000 69.355000 58.810000 69.555000 ;
        RECT 58.610000 69.765000 58.810000 69.965000 ;
        RECT 58.610000 70.175000 58.810000 70.375000 ;
        RECT 58.610000 70.585000 58.810000 70.785000 ;
        RECT 58.610000 70.995000 58.810000 71.195000 ;
        RECT 58.610000 71.405000 58.810000 71.605000 ;
        RECT 58.610000 71.815000 58.810000 72.015000 ;
        RECT 58.610000 72.225000 58.810000 72.425000 ;
        RECT 58.610000 72.635000 58.810000 72.835000 ;
        RECT 58.610000 73.045000 58.810000 73.245000 ;
        RECT 58.610000 73.450000 58.810000 73.650000 ;
        RECT 58.610000 73.855000 58.810000 74.055000 ;
        RECT 58.610000 74.260000 58.810000 74.460000 ;
        RECT 58.610000 74.665000 58.810000 74.865000 ;
        RECT 58.610000 75.070000 58.810000 75.270000 ;
        RECT 58.610000 75.475000 58.810000 75.675000 ;
        RECT 58.610000 75.880000 58.810000 76.080000 ;
        RECT 58.610000 76.285000 58.810000 76.485000 ;
        RECT 58.610000 76.690000 58.810000 76.890000 ;
        RECT 58.610000 77.095000 58.810000 77.295000 ;
        RECT 58.610000 77.500000 58.810000 77.700000 ;
        RECT 58.610000 77.905000 58.810000 78.105000 ;
        RECT 58.610000 78.310000 58.810000 78.510000 ;
        RECT 58.610000 78.715000 58.810000 78.915000 ;
        RECT 58.610000 79.120000 58.810000 79.320000 ;
        RECT 58.610000 79.525000 58.810000 79.725000 ;
        RECT 58.610000 79.930000 58.810000 80.130000 ;
        RECT 58.610000 80.335000 58.810000 80.535000 ;
        RECT 58.610000 80.740000 58.810000 80.940000 ;
        RECT 58.610000 81.145000 58.810000 81.345000 ;
        RECT 58.610000 81.550000 58.810000 81.750000 ;
        RECT 58.610000 81.955000 58.810000 82.155000 ;
        RECT 58.610000 82.360000 58.810000 82.560000 ;
        RECT 58.945000 17.860000 59.145000 18.060000 ;
        RECT 58.945000 18.290000 59.145000 18.490000 ;
        RECT 58.945000 18.720000 59.145000 18.920000 ;
        RECT 58.945000 19.150000 59.145000 19.350000 ;
        RECT 58.945000 19.580000 59.145000 19.780000 ;
        RECT 58.945000 20.010000 59.145000 20.210000 ;
        RECT 58.945000 20.440000 59.145000 20.640000 ;
        RECT 58.945000 20.870000 59.145000 21.070000 ;
        RECT 58.945000 21.300000 59.145000 21.500000 ;
        RECT 58.945000 21.730000 59.145000 21.930000 ;
        RECT 58.945000 22.160000 59.145000 22.360000 ;
        RECT 58.950000 83.055000 59.150000 83.255000 ;
        RECT 58.950000 83.455000 59.150000 83.655000 ;
        RECT 58.950000 83.855000 59.150000 84.055000 ;
        RECT 58.950000 84.255000 59.150000 84.455000 ;
        RECT 58.950000 84.655000 59.150000 84.855000 ;
        RECT 58.950000 85.055000 59.150000 85.255000 ;
        RECT 58.950000 85.455000 59.150000 85.655000 ;
        RECT 58.950000 85.855000 59.150000 86.055000 ;
        RECT 58.950000 86.255000 59.150000 86.455000 ;
        RECT 58.950000 86.660000 59.150000 86.860000 ;
        RECT 58.950000 87.065000 59.150000 87.265000 ;
        RECT 58.950000 87.470000 59.150000 87.670000 ;
        RECT 58.950000 87.875000 59.150000 88.075000 ;
        RECT 59.010000 68.125000 59.210000 68.325000 ;
        RECT 59.010000 68.535000 59.210000 68.735000 ;
        RECT 59.010000 68.945000 59.210000 69.145000 ;
        RECT 59.010000 69.355000 59.210000 69.555000 ;
        RECT 59.010000 69.765000 59.210000 69.965000 ;
        RECT 59.010000 70.175000 59.210000 70.375000 ;
        RECT 59.010000 70.585000 59.210000 70.785000 ;
        RECT 59.010000 70.995000 59.210000 71.195000 ;
        RECT 59.010000 71.405000 59.210000 71.605000 ;
        RECT 59.010000 71.815000 59.210000 72.015000 ;
        RECT 59.010000 72.225000 59.210000 72.425000 ;
        RECT 59.010000 72.635000 59.210000 72.835000 ;
        RECT 59.010000 73.045000 59.210000 73.245000 ;
        RECT 59.010000 73.450000 59.210000 73.650000 ;
        RECT 59.010000 73.855000 59.210000 74.055000 ;
        RECT 59.010000 74.260000 59.210000 74.460000 ;
        RECT 59.010000 74.665000 59.210000 74.865000 ;
        RECT 59.010000 75.070000 59.210000 75.270000 ;
        RECT 59.010000 75.475000 59.210000 75.675000 ;
        RECT 59.010000 75.880000 59.210000 76.080000 ;
        RECT 59.010000 76.285000 59.210000 76.485000 ;
        RECT 59.010000 76.690000 59.210000 76.890000 ;
        RECT 59.010000 77.095000 59.210000 77.295000 ;
        RECT 59.010000 77.500000 59.210000 77.700000 ;
        RECT 59.010000 77.905000 59.210000 78.105000 ;
        RECT 59.010000 78.310000 59.210000 78.510000 ;
        RECT 59.010000 78.715000 59.210000 78.915000 ;
        RECT 59.010000 79.120000 59.210000 79.320000 ;
        RECT 59.010000 79.525000 59.210000 79.725000 ;
        RECT 59.010000 79.930000 59.210000 80.130000 ;
        RECT 59.010000 80.335000 59.210000 80.535000 ;
        RECT 59.010000 80.740000 59.210000 80.940000 ;
        RECT 59.010000 81.145000 59.210000 81.345000 ;
        RECT 59.010000 81.550000 59.210000 81.750000 ;
        RECT 59.010000 81.955000 59.210000 82.155000 ;
        RECT 59.010000 82.360000 59.210000 82.560000 ;
        RECT 59.075000 88.410000 59.275000 88.610000 ;
        RECT 59.075000 88.835000 59.275000 89.035000 ;
        RECT 59.075000 89.265000 59.275000 89.465000 ;
        RECT 59.075000 89.695000 59.275000 89.895000 ;
        RECT 59.075000 90.125000 59.275000 90.325000 ;
        RECT 59.075000 90.555000 59.275000 90.755000 ;
        RECT 59.350000 17.860000 59.550000 18.060000 ;
        RECT 59.350000 18.290000 59.550000 18.490000 ;
        RECT 59.350000 18.720000 59.550000 18.920000 ;
        RECT 59.350000 19.150000 59.550000 19.350000 ;
        RECT 59.350000 19.580000 59.550000 19.780000 ;
        RECT 59.350000 20.010000 59.550000 20.210000 ;
        RECT 59.350000 20.440000 59.550000 20.640000 ;
        RECT 59.350000 20.870000 59.550000 21.070000 ;
        RECT 59.350000 21.300000 59.550000 21.500000 ;
        RECT 59.350000 21.730000 59.550000 21.930000 ;
        RECT 59.350000 22.160000 59.550000 22.360000 ;
        RECT 59.360000 83.055000 59.560000 83.255000 ;
        RECT 59.360000 83.455000 59.560000 83.655000 ;
        RECT 59.360000 83.855000 59.560000 84.055000 ;
        RECT 59.360000 84.255000 59.560000 84.455000 ;
        RECT 59.360000 84.655000 59.560000 84.855000 ;
        RECT 59.360000 85.055000 59.560000 85.255000 ;
        RECT 59.360000 85.455000 59.560000 85.655000 ;
        RECT 59.360000 85.855000 59.560000 86.055000 ;
        RECT 59.360000 86.255000 59.560000 86.455000 ;
        RECT 59.360000 86.660000 59.560000 86.860000 ;
        RECT 59.360000 87.065000 59.560000 87.265000 ;
        RECT 59.360000 87.470000 59.560000 87.670000 ;
        RECT 59.360000 87.875000 59.560000 88.075000 ;
        RECT 59.410000 68.125000 59.610000 68.325000 ;
        RECT 59.410000 68.535000 59.610000 68.735000 ;
        RECT 59.410000 68.945000 59.610000 69.145000 ;
        RECT 59.410000 69.355000 59.610000 69.555000 ;
        RECT 59.410000 69.765000 59.610000 69.965000 ;
        RECT 59.410000 70.175000 59.610000 70.375000 ;
        RECT 59.410000 70.585000 59.610000 70.785000 ;
        RECT 59.410000 70.995000 59.610000 71.195000 ;
        RECT 59.410000 71.405000 59.610000 71.605000 ;
        RECT 59.410000 71.815000 59.610000 72.015000 ;
        RECT 59.410000 72.225000 59.610000 72.425000 ;
        RECT 59.410000 72.635000 59.610000 72.835000 ;
        RECT 59.410000 73.045000 59.610000 73.245000 ;
        RECT 59.410000 73.450000 59.610000 73.650000 ;
        RECT 59.410000 73.855000 59.610000 74.055000 ;
        RECT 59.410000 74.260000 59.610000 74.460000 ;
        RECT 59.410000 74.665000 59.610000 74.865000 ;
        RECT 59.410000 75.070000 59.610000 75.270000 ;
        RECT 59.410000 75.475000 59.610000 75.675000 ;
        RECT 59.410000 75.880000 59.610000 76.080000 ;
        RECT 59.410000 76.285000 59.610000 76.485000 ;
        RECT 59.410000 76.690000 59.610000 76.890000 ;
        RECT 59.410000 77.095000 59.610000 77.295000 ;
        RECT 59.410000 77.500000 59.610000 77.700000 ;
        RECT 59.410000 77.905000 59.610000 78.105000 ;
        RECT 59.410000 78.310000 59.610000 78.510000 ;
        RECT 59.410000 78.715000 59.610000 78.915000 ;
        RECT 59.410000 79.120000 59.610000 79.320000 ;
        RECT 59.410000 79.525000 59.610000 79.725000 ;
        RECT 59.410000 79.930000 59.610000 80.130000 ;
        RECT 59.410000 80.335000 59.610000 80.535000 ;
        RECT 59.410000 80.740000 59.610000 80.940000 ;
        RECT 59.410000 81.145000 59.610000 81.345000 ;
        RECT 59.410000 81.550000 59.610000 81.750000 ;
        RECT 59.410000 81.955000 59.610000 82.155000 ;
        RECT 59.410000 82.360000 59.610000 82.560000 ;
        RECT 59.485000 88.410000 59.685000 88.610000 ;
        RECT 59.485000 88.835000 59.685000 89.035000 ;
        RECT 59.485000 89.265000 59.685000 89.465000 ;
        RECT 59.485000 89.695000 59.685000 89.895000 ;
        RECT 59.485000 90.125000 59.685000 90.325000 ;
        RECT 59.485000 90.555000 59.685000 90.755000 ;
        RECT 59.755000 17.860000 59.955000 18.060000 ;
        RECT 59.755000 18.290000 59.955000 18.490000 ;
        RECT 59.755000 18.720000 59.955000 18.920000 ;
        RECT 59.755000 19.150000 59.955000 19.350000 ;
        RECT 59.755000 19.580000 59.955000 19.780000 ;
        RECT 59.755000 20.010000 59.955000 20.210000 ;
        RECT 59.755000 20.440000 59.955000 20.640000 ;
        RECT 59.755000 20.870000 59.955000 21.070000 ;
        RECT 59.755000 21.300000 59.955000 21.500000 ;
        RECT 59.755000 21.730000 59.955000 21.930000 ;
        RECT 59.755000 22.160000 59.955000 22.360000 ;
        RECT 59.770000 83.055000 59.970000 83.255000 ;
        RECT 59.770000 83.455000 59.970000 83.655000 ;
        RECT 59.770000 83.855000 59.970000 84.055000 ;
        RECT 59.770000 84.255000 59.970000 84.455000 ;
        RECT 59.770000 84.655000 59.970000 84.855000 ;
        RECT 59.770000 85.055000 59.970000 85.255000 ;
        RECT 59.770000 85.455000 59.970000 85.655000 ;
        RECT 59.770000 85.855000 59.970000 86.055000 ;
        RECT 59.770000 86.255000 59.970000 86.455000 ;
        RECT 59.770000 86.660000 59.970000 86.860000 ;
        RECT 59.770000 87.065000 59.970000 87.265000 ;
        RECT 59.770000 87.470000 59.970000 87.670000 ;
        RECT 59.770000 87.875000 59.970000 88.075000 ;
        RECT 59.810000 68.125000 60.010000 68.325000 ;
        RECT 59.810000 68.535000 60.010000 68.735000 ;
        RECT 59.810000 68.945000 60.010000 69.145000 ;
        RECT 59.810000 69.355000 60.010000 69.555000 ;
        RECT 59.810000 69.765000 60.010000 69.965000 ;
        RECT 59.810000 70.175000 60.010000 70.375000 ;
        RECT 59.810000 70.585000 60.010000 70.785000 ;
        RECT 59.810000 70.995000 60.010000 71.195000 ;
        RECT 59.810000 71.405000 60.010000 71.605000 ;
        RECT 59.810000 71.815000 60.010000 72.015000 ;
        RECT 59.810000 72.225000 60.010000 72.425000 ;
        RECT 59.810000 72.635000 60.010000 72.835000 ;
        RECT 59.810000 73.045000 60.010000 73.245000 ;
        RECT 59.810000 73.450000 60.010000 73.650000 ;
        RECT 59.810000 73.855000 60.010000 74.055000 ;
        RECT 59.810000 74.260000 60.010000 74.460000 ;
        RECT 59.810000 74.665000 60.010000 74.865000 ;
        RECT 59.810000 75.070000 60.010000 75.270000 ;
        RECT 59.810000 75.475000 60.010000 75.675000 ;
        RECT 59.810000 75.880000 60.010000 76.080000 ;
        RECT 59.810000 76.285000 60.010000 76.485000 ;
        RECT 59.810000 76.690000 60.010000 76.890000 ;
        RECT 59.810000 77.095000 60.010000 77.295000 ;
        RECT 59.810000 77.500000 60.010000 77.700000 ;
        RECT 59.810000 77.905000 60.010000 78.105000 ;
        RECT 59.810000 78.310000 60.010000 78.510000 ;
        RECT 59.810000 78.715000 60.010000 78.915000 ;
        RECT 59.810000 79.120000 60.010000 79.320000 ;
        RECT 59.810000 79.525000 60.010000 79.725000 ;
        RECT 59.810000 79.930000 60.010000 80.130000 ;
        RECT 59.810000 80.335000 60.010000 80.535000 ;
        RECT 59.810000 80.740000 60.010000 80.940000 ;
        RECT 59.810000 81.145000 60.010000 81.345000 ;
        RECT 59.810000 81.550000 60.010000 81.750000 ;
        RECT 59.810000 81.955000 60.010000 82.155000 ;
        RECT 59.810000 82.360000 60.010000 82.560000 ;
        RECT 59.895000 88.410000 60.095000 88.610000 ;
        RECT 59.895000 88.835000 60.095000 89.035000 ;
        RECT 59.895000 89.265000 60.095000 89.465000 ;
        RECT 59.895000 89.695000 60.095000 89.895000 ;
        RECT 59.895000 90.125000 60.095000 90.325000 ;
        RECT 59.895000 90.555000 60.095000 90.755000 ;
        RECT 59.955000 91.015000 60.155000 91.215000 ;
        RECT 59.955000 91.445000 60.155000 91.645000 ;
        RECT 60.160000 17.860000 60.360000 18.060000 ;
        RECT 60.160000 18.290000 60.360000 18.490000 ;
        RECT 60.160000 18.720000 60.360000 18.920000 ;
        RECT 60.160000 19.150000 60.360000 19.350000 ;
        RECT 60.160000 19.580000 60.360000 19.780000 ;
        RECT 60.160000 20.010000 60.360000 20.210000 ;
        RECT 60.160000 20.440000 60.360000 20.640000 ;
        RECT 60.160000 20.870000 60.360000 21.070000 ;
        RECT 60.160000 21.300000 60.360000 21.500000 ;
        RECT 60.160000 21.730000 60.360000 21.930000 ;
        RECT 60.160000 22.160000 60.360000 22.360000 ;
        RECT 60.180000 83.055000 60.380000 83.255000 ;
        RECT 60.180000 83.455000 60.380000 83.655000 ;
        RECT 60.180000 83.855000 60.380000 84.055000 ;
        RECT 60.180000 84.255000 60.380000 84.455000 ;
        RECT 60.180000 84.655000 60.380000 84.855000 ;
        RECT 60.180000 85.055000 60.380000 85.255000 ;
        RECT 60.180000 85.455000 60.380000 85.655000 ;
        RECT 60.180000 85.855000 60.380000 86.055000 ;
        RECT 60.180000 86.255000 60.380000 86.455000 ;
        RECT 60.180000 86.660000 60.380000 86.860000 ;
        RECT 60.180000 87.065000 60.380000 87.265000 ;
        RECT 60.180000 87.470000 60.380000 87.670000 ;
        RECT 60.180000 87.875000 60.380000 88.075000 ;
        RECT 60.210000 68.125000 60.410000 68.325000 ;
        RECT 60.210000 68.535000 60.410000 68.735000 ;
        RECT 60.210000 68.945000 60.410000 69.145000 ;
        RECT 60.210000 69.355000 60.410000 69.555000 ;
        RECT 60.210000 69.765000 60.410000 69.965000 ;
        RECT 60.210000 70.175000 60.410000 70.375000 ;
        RECT 60.210000 70.585000 60.410000 70.785000 ;
        RECT 60.210000 70.995000 60.410000 71.195000 ;
        RECT 60.210000 71.405000 60.410000 71.605000 ;
        RECT 60.210000 71.815000 60.410000 72.015000 ;
        RECT 60.210000 72.225000 60.410000 72.425000 ;
        RECT 60.210000 72.635000 60.410000 72.835000 ;
        RECT 60.210000 73.045000 60.410000 73.245000 ;
        RECT 60.210000 73.450000 60.410000 73.650000 ;
        RECT 60.210000 73.855000 60.410000 74.055000 ;
        RECT 60.210000 74.260000 60.410000 74.460000 ;
        RECT 60.210000 74.665000 60.410000 74.865000 ;
        RECT 60.210000 75.070000 60.410000 75.270000 ;
        RECT 60.210000 75.475000 60.410000 75.675000 ;
        RECT 60.210000 75.880000 60.410000 76.080000 ;
        RECT 60.210000 76.285000 60.410000 76.485000 ;
        RECT 60.210000 76.690000 60.410000 76.890000 ;
        RECT 60.210000 77.095000 60.410000 77.295000 ;
        RECT 60.210000 77.500000 60.410000 77.700000 ;
        RECT 60.210000 77.905000 60.410000 78.105000 ;
        RECT 60.210000 78.310000 60.410000 78.510000 ;
        RECT 60.210000 78.715000 60.410000 78.915000 ;
        RECT 60.210000 79.120000 60.410000 79.320000 ;
        RECT 60.210000 79.525000 60.410000 79.725000 ;
        RECT 60.210000 79.930000 60.410000 80.130000 ;
        RECT 60.210000 80.335000 60.410000 80.535000 ;
        RECT 60.210000 80.740000 60.410000 80.940000 ;
        RECT 60.210000 81.145000 60.410000 81.345000 ;
        RECT 60.210000 81.550000 60.410000 81.750000 ;
        RECT 60.210000 81.955000 60.410000 82.155000 ;
        RECT 60.210000 82.360000 60.410000 82.560000 ;
        RECT 60.305000 88.410000 60.505000 88.610000 ;
        RECT 60.305000 88.835000 60.505000 89.035000 ;
        RECT 60.305000 89.265000 60.505000 89.465000 ;
        RECT 60.305000 89.695000 60.505000 89.895000 ;
        RECT 60.305000 90.125000 60.505000 90.325000 ;
        RECT 60.305000 90.555000 60.505000 90.755000 ;
        RECT 60.565000 17.860000 60.765000 18.060000 ;
        RECT 60.565000 18.290000 60.765000 18.490000 ;
        RECT 60.565000 18.720000 60.765000 18.920000 ;
        RECT 60.565000 19.150000 60.765000 19.350000 ;
        RECT 60.565000 19.580000 60.765000 19.780000 ;
        RECT 60.565000 20.010000 60.765000 20.210000 ;
        RECT 60.565000 20.440000 60.765000 20.640000 ;
        RECT 60.565000 20.870000 60.765000 21.070000 ;
        RECT 60.565000 21.300000 60.765000 21.500000 ;
        RECT 60.565000 21.730000 60.765000 21.930000 ;
        RECT 60.565000 22.160000 60.765000 22.360000 ;
        RECT 60.590000 83.055000 60.790000 83.255000 ;
        RECT 60.590000 83.455000 60.790000 83.655000 ;
        RECT 60.590000 83.855000 60.790000 84.055000 ;
        RECT 60.590000 84.255000 60.790000 84.455000 ;
        RECT 60.590000 84.655000 60.790000 84.855000 ;
        RECT 60.590000 85.055000 60.790000 85.255000 ;
        RECT 60.590000 85.455000 60.790000 85.655000 ;
        RECT 60.590000 85.855000 60.790000 86.055000 ;
        RECT 60.590000 86.255000 60.790000 86.455000 ;
        RECT 60.590000 86.660000 60.790000 86.860000 ;
        RECT 60.590000 87.065000 60.790000 87.265000 ;
        RECT 60.590000 87.470000 60.790000 87.670000 ;
        RECT 60.590000 87.875000 60.790000 88.075000 ;
        RECT 60.610000 68.125000 60.810000 68.325000 ;
        RECT 60.610000 68.535000 60.810000 68.735000 ;
        RECT 60.610000 68.945000 60.810000 69.145000 ;
        RECT 60.610000 69.355000 60.810000 69.555000 ;
        RECT 60.610000 69.765000 60.810000 69.965000 ;
        RECT 60.610000 70.175000 60.810000 70.375000 ;
        RECT 60.610000 70.585000 60.810000 70.785000 ;
        RECT 60.610000 70.995000 60.810000 71.195000 ;
        RECT 60.610000 71.405000 60.810000 71.605000 ;
        RECT 60.610000 71.815000 60.810000 72.015000 ;
        RECT 60.610000 72.225000 60.810000 72.425000 ;
        RECT 60.610000 72.635000 60.810000 72.835000 ;
        RECT 60.610000 73.045000 60.810000 73.245000 ;
        RECT 60.610000 73.450000 60.810000 73.650000 ;
        RECT 60.610000 73.855000 60.810000 74.055000 ;
        RECT 60.610000 74.260000 60.810000 74.460000 ;
        RECT 60.610000 74.665000 60.810000 74.865000 ;
        RECT 60.610000 75.070000 60.810000 75.270000 ;
        RECT 60.610000 75.475000 60.810000 75.675000 ;
        RECT 60.610000 75.880000 60.810000 76.080000 ;
        RECT 60.610000 76.285000 60.810000 76.485000 ;
        RECT 60.610000 76.690000 60.810000 76.890000 ;
        RECT 60.610000 77.095000 60.810000 77.295000 ;
        RECT 60.610000 77.500000 60.810000 77.700000 ;
        RECT 60.610000 77.905000 60.810000 78.105000 ;
        RECT 60.610000 78.310000 60.810000 78.510000 ;
        RECT 60.610000 78.715000 60.810000 78.915000 ;
        RECT 60.610000 79.120000 60.810000 79.320000 ;
        RECT 60.610000 79.525000 60.810000 79.725000 ;
        RECT 60.610000 79.930000 60.810000 80.130000 ;
        RECT 60.610000 80.335000 60.810000 80.535000 ;
        RECT 60.610000 80.740000 60.810000 80.940000 ;
        RECT 60.610000 81.145000 60.810000 81.345000 ;
        RECT 60.610000 81.550000 60.810000 81.750000 ;
        RECT 60.610000 81.955000 60.810000 82.155000 ;
        RECT 60.610000 82.360000 60.810000 82.560000 ;
        RECT 60.715000 88.410000 60.915000 88.610000 ;
        RECT 60.715000 88.835000 60.915000 89.035000 ;
        RECT 60.715000 89.265000 60.915000 89.465000 ;
        RECT 60.715000 89.695000 60.915000 89.895000 ;
        RECT 60.715000 90.125000 60.915000 90.325000 ;
        RECT 60.715000 90.555000 60.915000 90.755000 ;
        RECT 60.735000 91.015000 60.935000 91.215000 ;
        RECT 60.735000 91.445000 60.935000 91.645000 ;
        RECT 60.970000 17.860000 61.170000 18.060000 ;
        RECT 60.970000 18.290000 61.170000 18.490000 ;
        RECT 60.970000 18.720000 61.170000 18.920000 ;
        RECT 60.970000 19.150000 61.170000 19.350000 ;
        RECT 60.970000 19.580000 61.170000 19.780000 ;
        RECT 60.970000 20.010000 61.170000 20.210000 ;
        RECT 60.970000 20.440000 61.170000 20.640000 ;
        RECT 60.970000 20.870000 61.170000 21.070000 ;
        RECT 60.970000 21.300000 61.170000 21.500000 ;
        RECT 60.970000 21.730000 61.170000 21.930000 ;
        RECT 60.970000 22.160000 61.170000 22.360000 ;
        RECT 61.010000 68.125000 61.210000 68.325000 ;
        RECT 61.010000 68.535000 61.210000 68.735000 ;
        RECT 61.010000 68.945000 61.210000 69.145000 ;
        RECT 61.010000 69.355000 61.210000 69.555000 ;
        RECT 61.010000 69.765000 61.210000 69.965000 ;
        RECT 61.010000 70.175000 61.210000 70.375000 ;
        RECT 61.010000 70.585000 61.210000 70.785000 ;
        RECT 61.010000 70.995000 61.210000 71.195000 ;
        RECT 61.010000 71.405000 61.210000 71.605000 ;
        RECT 61.010000 71.815000 61.210000 72.015000 ;
        RECT 61.010000 72.225000 61.210000 72.425000 ;
        RECT 61.010000 72.635000 61.210000 72.835000 ;
        RECT 61.010000 73.045000 61.210000 73.245000 ;
        RECT 61.010000 73.450000 61.210000 73.650000 ;
        RECT 61.010000 73.855000 61.210000 74.055000 ;
        RECT 61.010000 74.260000 61.210000 74.460000 ;
        RECT 61.010000 74.665000 61.210000 74.865000 ;
        RECT 61.010000 75.070000 61.210000 75.270000 ;
        RECT 61.010000 75.475000 61.210000 75.675000 ;
        RECT 61.010000 75.880000 61.210000 76.080000 ;
        RECT 61.010000 76.285000 61.210000 76.485000 ;
        RECT 61.010000 76.690000 61.210000 76.890000 ;
        RECT 61.010000 77.095000 61.210000 77.295000 ;
        RECT 61.010000 77.500000 61.210000 77.700000 ;
        RECT 61.010000 77.905000 61.210000 78.105000 ;
        RECT 61.010000 78.310000 61.210000 78.510000 ;
        RECT 61.010000 78.715000 61.210000 78.915000 ;
        RECT 61.010000 79.120000 61.210000 79.320000 ;
        RECT 61.010000 79.525000 61.210000 79.725000 ;
        RECT 61.010000 79.930000 61.210000 80.130000 ;
        RECT 61.010000 80.335000 61.210000 80.535000 ;
        RECT 61.010000 80.740000 61.210000 80.940000 ;
        RECT 61.010000 81.145000 61.210000 81.345000 ;
        RECT 61.010000 81.550000 61.210000 81.750000 ;
        RECT 61.010000 81.955000 61.210000 82.155000 ;
        RECT 61.010000 82.360000 61.210000 82.560000 ;
        RECT 61.215000 82.855000 61.415000 83.055000 ;
        RECT 61.215000 83.265000 61.415000 83.465000 ;
        RECT 61.215000 83.675000 61.415000 83.875000 ;
        RECT 61.215000 84.085000 61.415000 84.285000 ;
        RECT 61.215000 84.495000 61.415000 84.695000 ;
        RECT 61.215000 84.905000 61.415000 85.105000 ;
        RECT 61.215000 85.315000 61.415000 85.515000 ;
        RECT 61.215000 85.725000 61.415000 85.925000 ;
        RECT 61.215000 86.135000 61.415000 86.335000 ;
        RECT 61.215000 86.545000 61.415000 86.745000 ;
        RECT 61.215000 86.955000 61.415000 87.155000 ;
        RECT 61.215000 87.365000 61.415000 87.565000 ;
        RECT 61.215000 87.775000 61.415000 87.975000 ;
        RECT 61.215000 88.185000 61.415000 88.385000 ;
        RECT 61.215000 88.595000 61.415000 88.795000 ;
        RECT 61.215000 89.005000 61.415000 89.205000 ;
        RECT 61.215000 89.415000 61.415000 89.615000 ;
        RECT 61.215000 89.825000 61.415000 90.025000 ;
        RECT 61.215000 90.235000 61.415000 90.435000 ;
        RECT 61.215000 90.645000 61.415000 90.845000 ;
        RECT 61.215000 91.055000 61.415000 91.255000 ;
        RECT 61.215000 91.465000 61.415000 91.665000 ;
        RECT 61.215000 91.875000 61.415000 92.075000 ;
        RECT 61.215000 92.285000 61.415000 92.485000 ;
        RECT 61.215000 92.695000 61.415000 92.895000 ;
        RECT 61.375000 17.860000 61.575000 18.060000 ;
        RECT 61.375000 18.290000 61.575000 18.490000 ;
        RECT 61.375000 18.720000 61.575000 18.920000 ;
        RECT 61.375000 19.150000 61.575000 19.350000 ;
        RECT 61.375000 19.580000 61.575000 19.780000 ;
        RECT 61.375000 20.010000 61.575000 20.210000 ;
        RECT 61.375000 20.440000 61.575000 20.640000 ;
        RECT 61.375000 20.870000 61.575000 21.070000 ;
        RECT 61.375000 21.300000 61.575000 21.500000 ;
        RECT 61.375000 21.730000 61.575000 21.930000 ;
        RECT 61.375000 22.160000 61.575000 22.360000 ;
        RECT 61.410000 68.125000 61.610000 68.325000 ;
        RECT 61.410000 68.535000 61.610000 68.735000 ;
        RECT 61.410000 68.945000 61.610000 69.145000 ;
        RECT 61.410000 69.355000 61.610000 69.555000 ;
        RECT 61.410000 69.765000 61.610000 69.965000 ;
        RECT 61.410000 70.175000 61.610000 70.375000 ;
        RECT 61.410000 70.585000 61.610000 70.785000 ;
        RECT 61.410000 70.995000 61.610000 71.195000 ;
        RECT 61.410000 71.405000 61.610000 71.605000 ;
        RECT 61.410000 71.815000 61.610000 72.015000 ;
        RECT 61.410000 72.225000 61.610000 72.425000 ;
        RECT 61.410000 72.635000 61.610000 72.835000 ;
        RECT 61.410000 73.045000 61.610000 73.245000 ;
        RECT 61.410000 73.450000 61.610000 73.650000 ;
        RECT 61.410000 73.855000 61.610000 74.055000 ;
        RECT 61.410000 74.260000 61.610000 74.460000 ;
        RECT 61.410000 74.665000 61.610000 74.865000 ;
        RECT 61.410000 75.070000 61.610000 75.270000 ;
        RECT 61.410000 75.475000 61.610000 75.675000 ;
        RECT 61.410000 75.880000 61.610000 76.080000 ;
        RECT 61.410000 76.285000 61.610000 76.485000 ;
        RECT 61.410000 76.690000 61.610000 76.890000 ;
        RECT 61.410000 77.095000 61.610000 77.295000 ;
        RECT 61.410000 77.500000 61.610000 77.700000 ;
        RECT 61.410000 77.905000 61.610000 78.105000 ;
        RECT 61.410000 78.310000 61.610000 78.510000 ;
        RECT 61.410000 78.715000 61.610000 78.915000 ;
        RECT 61.410000 79.120000 61.610000 79.320000 ;
        RECT 61.410000 79.525000 61.610000 79.725000 ;
        RECT 61.410000 79.930000 61.610000 80.130000 ;
        RECT 61.410000 80.335000 61.610000 80.535000 ;
        RECT 61.410000 80.740000 61.610000 80.940000 ;
        RECT 61.410000 81.145000 61.610000 81.345000 ;
        RECT 61.410000 81.550000 61.610000 81.750000 ;
        RECT 61.410000 81.955000 61.610000 82.155000 ;
        RECT 61.410000 82.360000 61.610000 82.560000 ;
        RECT 61.620000 82.855000 61.820000 83.055000 ;
        RECT 61.620000 83.265000 61.820000 83.465000 ;
        RECT 61.620000 83.675000 61.820000 83.875000 ;
        RECT 61.620000 84.085000 61.820000 84.285000 ;
        RECT 61.620000 84.495000 61.820000 84.695000 ;
        RECT 61.620000 84.905000 61.820000 85.105000 ;
        RECT 61.620000 85.315000 61.820000 85.515000 ;
        RECT 61.620000 85.725000 61.820000 85.925000 ;
        RECT 61.620000 86.135000 61.820000 86.335000 ;
        RECT 61.620000 86.545000 61.820000 86.745000 ;
        RECT 61.620000 86.955000 61.820000 87.155000 ;
        RECT 61.620000 87.365000 61.820000 87.565000 ;
        RECT 61.620000 87.775000 61.820000 87.975000 ;
        RECT 61.620000 88.185000 61.820000 88.385000 ;
        RECT 61.620000 88.595000 61.820000 88.795000 ;
        RECT 61.620000 89.005000 61.820000 89.205000 ;
        RECT 61.620000 89.415000 61.820000 89.615000 ;
        RECT 61.620000 89.825000 61.820000 90.025000 ;
        RECT 61.620000 90.235000 61.820000 90.435000 ;
        RECT 61.620000 90.645000 61.820000 90.845000 ;
        RECT 61.620000 91.055000 61.820000 91.255000 ;
        RECT 61.620000 91.465000 61.820000 91.665000 ;
        RECT 61.620000 91.875000 61.820000 92.075000 ;
        RECT 61.620000 92.285000 61.820000 92.485000 ;
        RECT 61.620000 92.695000 61.820000 92.895000 ;
        RECT 61.780000 17.860000 61.980000 18.060000 ;
        RECT 61.780000 18.290000 61.980000 18.490000 ;
        RECT 61.780000 18.720000 61.980000 18.920000 ;
        RECT 61.780000 19.150000 61.980000 19.350000 ;
        RECT 61.780000 19.580000 61.980000 19.780000 ;
        RECT 61.780000 20.010000 61.980000 20.210000 ;
        RECT 61.780000 20.440000 61.980000 20.640000 ;
        RECT 61.780000 20.870000 61.980000 21.070000 ;
        RECT 61.780000 21.300000 61.980000 21.500000 ;
        RECT 61.780000 21.730000 61.980000 21.930000 ;
        RECT 61.780000 22.160000 61.980000 22.360000 ;
        RECT 61.810000 68.125000 62.010000 68.325000 ;
        RECT 61.810000 68.535000 62.010000 68.735000 ;
        RECT 61.810000 68.945000 62.010000 69.145000 ;
        RECT 61.810000 69.355000 62.010000 69.555000 ;
        RECT 61.810000 69.765000 62.010000 69.965000 ;
        RECT 61.810000 70.175000 62.010000 70.375000 ;
        RECT 61.810000 70.585000 62.010000 70.785000 ;
        RECT 61.810000 70.995000 62.010000 71.195000 ;
        RECT 61.810000 71.405000 62.010000 71.605000 ;
        RECT 61.810000 71.815000 62.010000 72.015000 ;
        RECT 61.810000 72.225000 62.010000 72.425000 ;
        RECT 61.810000 72.635000 62.010000 72.835000 ;
        RECT 61.810000 73.045000 62.010000 73.245000 ;
        RECT 61.810000 73.450000 62.010000 73.650000 ;
        RECT 61.810000 73.855000 62.010000 74.055000 ;
        RECT 61.810000 74.260000 62.010000 74.460000 ;
        RECT 61.810000 74.665000 62.010000 74.865000 ;
        RECT 61.810000 75.070000 62.010000 75.270000 ;
        RECT 61.810000 75.475000 62.010000 75.675000 ;
        RECT 61.810000 75.880000 62.010000 76.080000 ;
        RECT 61.810000 76.285000 62.010000 76.485000 ;
        RECT 61.810000 76.690000 62.010000 76.890000 ;
        RECT 61.810000 77.095000 62.010000 77.295000 ;
        RECT 61.810000 77.500000 62.010000 77.700000 ;
        RECT 61.810000 77.905000 62.010000 78.105000 ;
        RECT 61.810000 78.310000 62.010000 78.510000 ;
        RECT 61.810000 78.715000 62.010000 78.915000 ;
        RECT 61.810000 79.120000 62.010000 79.320000 ;
        RECT 61.810000 79.525000 62.010000 79.725000 ;
        RECT 61.810000 79.930000 62.010000 80.130000 ;
        RECT 61.810000 80.335000 62.010000 80.535000 ;
        RECT 61.810000 80.740000 62.010000 80.940000 ;
        RECT 61.810000 81.145000 62.010000 81.345000 ;
        RECT 61.810000 81.550000 62.010000 81.750000 ;
        RECT 61.810000 81.955000 62.010000 82.155000 ;
        RECT 61.810000 82.360000 62.010000 82.560000 ;
        RECT 62.025000 82.855000 62.225000 83.055000 ;
        RECT 62.025000 83.265000 62.225000 83.465000 ;
        RECT 62.025000 83.675000 62.225000 83.875000 ;
        RECT 62.025000 84.085000 62.225000 84.285000 ;
        RECT 62.025000 84.495000 62.225000 84.695000 ;
        RECT 62.025000 84.905000 62.225000 85.105000 ;
        RECT 62.025000 85.315000 62.225000 85.515000 ;
        RECT 62.025000 85.725000 62.225000 85.925000 ;
        RECT 62.025000 86.135000 62.225000 86.335000 ;
        RECT 62.025000 86.545000 62.225000 86.745000 ;
        RECT 62.025000 86.955000 62.225000 87.155000 ;
        RECT 62.025000 87.365000 62.225000 87.565000 ;
        RECT 62.025000 87.775000 62.225000 87.975000 ;
        RECT 62.025000 88.185000 62.225000 88.385000 ;
        RECT 62.025000 88.595000 62.225000 88.795000 ;
        RECT 62.025000 89.005000 62.225000 89.205000 ;
        RECT 62.025000 89.415000 62.225000 89.615000 ;
        RECT 62.025000 89.825000 62.225000 90.025000 ;
        RECT 62.025000 90.235000 62.225000 90.435000 ;
        RECT 62.025000 90.645000 62.225000 90.845000 ;
        RECT 62.025000 91.055000 62.225000 91.255000 ;
        RECT 62.025000 91.465000 62.225000 91.665000 ;
        RECT 62.025000 91.875000 62.225000 92.075000 ;
        RECT 62.025000 92.285000 62.225000 92.485000 ;
        RECT 62.025000 92.695000 62.225000 92.895000 ;
        RECT 62.185000 17.860000 62.385000 18.060000 ;
        RECT 62.185000 18.290000 62.385000 18.490000 ;
        RECT 62.185000 18.720000 62.385000 18.920000 ;
        RECT 62.185000 19.150000 62.385000 19.350000 ;
        RECT 62.185000 19.580000 62.385000 19.780000 ;
        RECT 62.185000 20.010000 62.385000 20.210000 ;
        RECT 62.185000 20.440000 62.385000 20.640000 ;
        RECT 62.185000 20.870000 62.385000 21.070000 ;
        RECT 62.185000 21.300000 62.385000 21.500000 ;
        RECT 62.185000 21.730000 62.385000 21.930000 ;
        RECT 62.185000 22.160000 62.385000 22.360000 ;
        RECT 62.210000 68.125000 62.410000 68.325000 ;
        RECT 62.210000 68.535000 62.410000 68.735000 ;
        RECT 62.210000 68.945000 62.410000 69.145000 ;
        RECT 62.210000 69.355000 62.410000 69.555000 ;
        RECT 62.210000 69.765000 62.410000 69.965000 ;
        RECT 62.210000 70.175000 62.410000 70.375000 ;
        RECT 62.210000 70.585000 62.410000 70.785000 ;
        RECT 62.210000 70.995000 62.410000 71.195000 ;
        RECT 62.210000 71.405000 62.410000 71.605000 ;
        RECT 62.210000 71.815000 62.410000 72.015000 ;
        RECT 62.210000 72.225000 62.410000 72.425000 ;
        RECT 62.210000 72.635000 62.410000 72.835000 ;
        RECT 62.210000 73.045000 62.410000 73.245000 ;
        RECT 62.210000 73.450000 62.410000 73.650000 ;
        RECT 62.210000 73.855000 62.410000 74.055000 ;
        RECT 62.210000 74.260000 62.410000 74.460000 ;
        RECT 62.210000 74.665000 62.410000 74.865000 ;
        RECT 62.210000 75.070000 62.410000 75.270000 ;
        RECT 62.210000 75.475000 62.410000 75.675000 ;
        RECT 62.210000 75.880000 62.410000 76.080000 ;
        RECT 62.210000 76.285000 62.410000 76.485000 ;
        RECT 62.210000 76.690000 62.410000 76.890000 ;
        RECT 62.210000 77.095000 62.410000 77.295000 ;
        RECT 62.210000 77.500000 62.410000 77.700000 ;
        RECT 62.210000 77.905000 62.410000 78.105000 ;
        RECT 62.210000 78.310000 62.410000 78.510000 ;
        RECT 62.210000 78.715000 62.410000 78.915000 ;
        RECT 62.210000 79.120000 62.410000 79.320000 ;
        RECT 62.210000 79.525000 62.410000 79.725000 ;
        RECT 62.210000 79.930000 62.410000 80.130000 ;
        RECT 62.210000 80.335000 62.410000 80.535000 ;
        RECT 62.210000 80.740000 62.410000 80.940000 ;
        RECT 62.210000 81.145000 62.410000 81.345000 ;
        RECT 62.210000 81.550000 62.410000 81.750000 ;
        RECT 62.210000 81.955000 62.410000 82.155000 ;
        RECT 62.210000 82.360000 62.410000 82.560000 ;
        RECT 62.430000 82.855000 62.630000 83.055000 ;
        RECT 62.430000 83.265000 62.630000 83.465000 ;
        RECT 62.430000 83.675000 62.630000 83.875000 ;
        RECT 62.430000 84.085000 62.630000 84.285000 ;
        RECT 62.430000 84.495000 62.630000 84.695000 ;
        RECT 62.430000 84.905000 62.630000 85.105000 ;
        RECT 62.430000 85.315000 62.630000 85.515000 ;
        RECT 62.430000 85.725000 62.630000 85.925000 ;
        RECT 62.430000 86.135000 62.630000 86.335000 ;
        RECT 62.430000 86.545000 62.630000 86.745000 ;
        RECT 62.430000 86.955000 62.630000 87.155000 ;
        RECT 62.430000 87.365000 62.630000 87.565000 ;
        RECT 62.430000 87.775000 62.630000 87.975000 ;
        RECT 62.430000 88.185000 62.630000 88.385000 ;
        RECT 62.430000 88.595000 62.630000 88.795000 ;
        RECT 62.430000 89.005000 62.630000 89.205000 ;
        RECT 62.430000 89.415000 62.630000 89.615000 ;
        RECT 62.430000 89.825000 62.630000 90.025000 ;
        RECT 62.430000 90.235000 62.630000 90.435000 ;
        RECT 62.430000 90.645000 62.630000 90.845000 ;
        RECT 62.430000 91.055000 62.630000 91.255000 ;
        RECT 62.430000 91.465000 62.630000 91.665000 ;
        RECT 62.430000 91.875000 62.630000 92.075000 ;
        RECT 62.430000 92.285000 62.630000 92.485000 ;
        RECT 62.430000 92.695000 62.630000 92.895000 ;
        RECT 62.590000 17.860000 62.790000 18.060000 ;
        RECT 62.590000 18.290000 62.790000 18.490000 ;
        RECT 62.590000 18.720000 62.790000 18.920000 ;
        RECT 62.590000 19.150000 62.790000 19.350000 ;
        RECT 62.590000 19.580000 62.790000 19.780000 ;
        RECT 62.590000 20.010000 62.790000 20.210000 ;
        RECT 62.590000 20.440000 62.790000 20.640000 ;
        RECT 62.590000 20.870000 62.790000 21.070000 ;
        RECT 62.590000 21.300000 62.790000 21.500000 ;
        RECT 62.590000 21.730000 62.790000 21.930000 ;
        RECT 62.590000 22.160000 62.790000 22.360000 ;
        RECT 62.610000 68.125000 62.810000 68.325000 ;
        RECT 62.610000 68.535000 62.810000 68.735000 ;
        RECT 62.610000 68.945000 62.810000 69.145000 ;
        RECT 62.610000 69.355000 62.810000 69.555000 ;
        RECT 62.610000 69.765000 62.810000 69.965000 ;
        RECT 62.610000 70.175000 62.810000 70.375000 ;
        RECT 62.610000 70.585000 62.810000 70.785000 ;
        RECT 62.610000 70.995000 62.810000 71.195000 ;
        RECT 62.610000 71.405000 62.810000 71.605000 ;
        RECT 62.610000 71.815000 62.810000 72.015000 ;
        RECT 62.610000 72.225000 62.810000 72.425000 ;
        RECT 62.610000 72.635000 62.810000 72.835000 ;
        RECT 62.610000 73.045000 62.810000 73.245000 ;
        RECT 62.610000 73.450000 62.810000 73.650000 ;
        RECT 62.610000 73.855000 62.810000 74.055000 ;
        RECT 62.610000 74.260000 62.810000 74.460000 ;
        RECT 62.610000 74.665000 62.810000 74.865000 ;
        RECT 62.610000 75.070000 62.810000 75.270000 ;
        RECT 62.610000 75.475000 62.810000 75.675000 ;
        RECT 62.610000 75.880000 62.810000 76.080000 ;
        RECT 62.610000 76.285000 62.810000 76.485000 ;
        RECT 62.610000 76.690000 62.810000 76.890000 ;
        RECT 62.610000 77.095000 62.810000 77.295000 ;
        RECT 62.610000 77.500000 62.810000 77.700000 ;
        RECT 62.610000 77.905000 62.810000 78.105000 ;
        RECT 62.610000 78.310000 62.810000 78.510000 ;
        RECT 62.610000 78.715000 62.810000 78.915000 ;
        RECT 62.610000 79.120000 62.810000 79.320000 ;
        RECT 62.610000 79.525000 62.810000 79.725000 ;
        RECT 62.610000 79.930000 62.810000 80.130000 ;
        RECT 62.610000 80.335000 62.810000 80.535000 ;
        RECT 62.610000 80.740000 62.810000 80.940000 ;
        RECT 62.610000 81.145000 62.810000 81.345000 ;
        RECT 62.610000 81.550000 62.810000 81.750000 ;
        RECT 62.610000 81.955000 62.810000 82.155000 ;
        RECT 62.610000 82.360000 62.810000 82.560000 ;
        RECT 62.840000 82.855000 63.040000 83.055000 ;
        RECT 62.840000 83.265000 63.040000 83.465000 ;
        RECT 62.840000 83.675000 63.040000 83.875000 ;
        RECT 62.840000 84.085000 63.040000 84.285000 ;
        RECT 62.840000 84.495000 63.040000 84.695000 ;
        RECT 62.840000 84.905000 63.040000 85.105000 ;
        RECT 62.840000 85.315000 63.040000 85.515000 ;
        RECT 62.840000 85.725000 63.040000 85.925000 ;
        RECT 62.840000 86.135000 63.040000 86.335000 ;
        RECT 62.840000 86.545000 63.040000 86.745000 ;
        RECT 62.840000 86.955000 63.040000 87.155000 ;
        RECT 62.840000 87.365000 63.040000 87.565000 ;
        RECT 62.840000 87.775000 63.040000 87.975000 ;
        RECT 62.840000 88.185000 63.040000 88.385000 ;
        RECT 62.840000 88.595000 63.040000 88.795000 ;
        RECT 62.840000 89.005000 63.040000 89.205000 ;
        RECT 62.840000 89.415000 63.040000 89.615000 ;
        RECT 62.840000 89.825000 63.040000 90.025000 ;
        RECT 62.840000 90.235000 63.040000 90.435000 ;
        RECT 62.840000 90.645000 63.040000 90.845000 ;
        RECT 62.840000 91.055000 63.040000 91.255000 ;
        RECT 62.840000 91.465000 63.040000 91.665000 ;
        RECT 62.840000 91.875000 63.040000 92.075000 ;
        RECT 62.840000 92.285000 63.040000 92.485000 ;
        RECT 62.840000 92.695000 63.040000 92.895000 ;
        RECT 62.995000 17.860000 63.195000 18.060000 ;
        RECT 62.995000 18.290000 63.195000 18.490000 ;
        RECT 62.995000 18.720000 63.195000 18.920000 ;
        RECT 62.995000 19.150000 63.195000 19.350000 ;
        RECT 62.995000 19.580000 63.195000 19.780000 ;
        RECT 62.995000 20.010000 63.195000 20.210000 ;
        RECT 62.995000 20.440000 63.195000 20.640000 ;
        RECT 62.995000 20.870000 63.195000 21.070000 ;
        RECT 62.995000 21.300000 63.195000 21.500000 ;
        RECT 62.995000 21.730000 63.195000 21.930000 ;
        RECT 62.995000 22.160000 63.195000 22.360000 ;
        RECT 63.010000 68.125000 63.210000 68.325000 ;
        RECT 63.010000 68.535000 63.210000 68.735000 ;
        RECT 63.010000 68.945000 63.210000 69.145000 ;
        RECT 63.010000 69.355000 63.210000 69.555000 ;
        RECT 63.010000 69.765000 63.210000 69.965000 ;
        RECT 63.010000 70.175000 63.210000 70.375000 ;
        RECT 63.010000 70.585000 63.210000 70.785000 ;
        RECT 63.010000 70.995000 63.210000 71.195000 ;
        RECT 63.010000 71.405000 63.210000 71.605000 ;
        RECT 63.010000 71.815000 63.210000 72.015000 ;
        RECT 63.010000 72.225000 63.210000 72.425000 ;
        RECT 63.010000 72.635000 63.210000 72.835000 ;
        RECT 63.010000 73.045000 63.210000 73.245000 ;
        RECT 63.010000 73.450000 63.210000 73.650000 ;
        RECT 63.010000 73.855000 63.210000 74.055000 ;
        RECT 63.010000 74.260000 63.210000 74.460000 ;
        RECT 63.010000 74.665000 63.210000 74.865000 ;
        RECT 63.010000 75.070000 63.210000 75.270000 ;
        RECT 63.010000 75.475000 63.210000 75.675000 ;
        RECT 63.010000 75.880000 63.210000 76.080000 ;
        RECT 63.010000 76.285000 63.210000 76.485000 ;
        RECT 63.010000 76.690000 63.210000 76.890000 ;
        RECT 63.010000 77.095000 63.210000 77.295000 ;
        RECT 63.010000 77.500000 63.210000 77.700000 ;
        RECT 63.010000 77.905000 63.210000 78.105000 ;
        RECT 63.010000 78.310000 63.210000 78.510000 ;
        RECT 63.010000 78.715000 63.210000 78.915000 ;
        RECT 63.010000 79.120000 63.210000 79.320000 ;
        RECT 63.010000 79.525000 63.210000 79.725000 ;
        RECT 63.010000 79.930000 63.210000 80.130000 ;
        RECT 63.010000 80.335000 63.210000 80.535000 ;
        RECT 63.010000 80.740000 63.210000 80.940000 ;
        RECT 63.010000 81.145000 63.210000 81.345000 ;
        RECT 63.010000 81.550000 63.210000 81.750000 ;
        RECT 63.010000 81.955000 63.210000 82.155000 ;
        RECT 63.010000 82.360000 63.210000 82.560000 ;
        RECT 63.250000 82.855000 63.450000 83.055000 ;
        RECT 63.250000 83.265000 63.450000 83.465000 ;
        RECT 63.250000 83.675000 63.450000 83.875000 ;
        RECT 63.250000 84.085000 63.450000 84.285000 ;
        RECT 63.250000 84.495000 63.450000 84.695000 ;
        RECT 63.250000 84.905000 63.450000 85.105000 ;
        RECT 63.250000 85.315000 63.450000 85.515000 ;
        RECT 63.250000 85.725000 63.450000 85.925000 ;
        RECT 63.250000 86.135000 63.450000 86.335000 ;
        RECT 63.250000 86.545000 63.450000 86.745000 ;
        RECT 63.250000 86.955000 63.450000 87.155000 ;
        RECT 63.250000 87.365000 63.450000 87.565000 ;
        RECT 63.250000 87.775000 63.450000 87.975000 ;
        RECT 63.250000 88.185000 63.450000 88.385000 ;
        RECT 63.250000 88.595000 63.450000 88.795000 ;
        RECT 63.250000 89.005000 63.450000 89.205000 ;
        RECT 63.250000 89.415000 63.450000 89.615000 ;
        RECT 63.250000 89.825000 63.450000 90.025000 ;
        RECT 63.250000 90.235000 63.450000 90.435000 ;
        RECT 63.250000 90.645000 63.450000 90.845000 ;
        RECT 63.250000 91.055000 63.450000 91.255000 ;
        RECT 63.250000 91.465000 63.450000 91.665000 ;
        RECT 63.250000 91.875000 63.450000 92.075000 ;
        RECT 63.250000 92.285000 63.450000 92.485000 ;
        RECT 63.250000 92.695000 63.450000 92.895000 ;
        RECT 63.400000 17.860000 63.600000 18.060000 ;
        RECT 63.400000 18.290000 63.600000 18.490000 ;
        RECT 63.400000 18.720000 63.600000 18.920000 ;
        RECT 63.400000 19.150000 63.600000 19.350000 ;
        RECT 63.400000 19.580000 63.600000 19.780000 ;
        RECT 63.400000 20.010000 63.600000 20.210000 ;
        RECT 63.400000 20.440000 63.600000 20.640000 ;
        RECT 63.400000 20.870000 63.600000 21.070000 ;
        RECT 63.400000 21.300000 63.600000 21.500000 ;
        RECT 63.400000 21.730000 63.600000 21.930000 ;
        RECT 63.400000 22.160000 63.600000 22.360000 ;
        RECT 63.410000 68.125000 63.610000 68.325000 ;
        RECT 63.410000 68.535000 63.610000 68.735000 ;
        RECT 63.410000 68.945000 63.610000 69.145000 ;
        RECT 63.410000 69.355000 63.610000 69.555000 ;
        RECT 63.410000 69.765000 63.610000 69.965000 ;
        RECT 63.410000 70.175000 63.610000 70.375000 ;
        RECT 63.410000 70.585000 63.610000 70.785000 ;
        RECT 63.410000 70.995000 63.610000 71.195000 ;
        RECT 63.410000 71.405000 63.610000 71.605000 ;
        RECT 63.410000 71.815000 63.610000 72.015000 ;
        RECT 63.410000 72.225000 63.610000 72.425000 ;
        RECT 63.410000 72.635000 63.610000 72.835000 ;
        RECT 63.410000 73.045000 63.610000 73.245000 ;
        RECT 63.410000 73.450000 63.610000 73.650000 ;
        RECT 63.410000 73.855000 63.610000 74.055000 ;
        RECT 63.410000 74.260000 63.610000 74.460000 ;
        RECT 63.410000 74.665000 63.610000 74.865000 ;
        RECT 63.410000 75.070000 63.610000 75.270000 ;
        RECT 63.410000 75.475000 63.610000 75.675000 ;
        RECT 63.410000 75.880000 63.610000 76.080000 ;
        RECT 63.410000 76.285000 63.610000 76.485000 ;
        RECT 63.410000 76.690000 63.610000 76.890000 ;
        RECT 63.410000 77.095000 63.610000 77.295000 ;
        RECT 63.410000 77.500000 63.610000 77.700000 ;
        RECT 63.410000 77.905000 63.610000 78.105000 ;
        RECT 63.410000 78.310000 63.610000 78.510000 ;
        RECT 63.410000 78.715000 63.610000 78.915000 ;
        RECT 63.410000 79.120000 63.610000 79.320000 ;
        RECT 63.410000 79.525000 63.610000 79.725000 ;
        RECT 63.410000 79.930000 63.610000 80.130000 ;
        RECT 63.410000 80.335000 63.610000 80.535000 ;
        RECT 63.410000 80.740000 63.610000 80.940000 ;
        RECT 63.410000 81.145000 63.610000 81.345000 ;
        RECT 63.410000 81.550000 63.610000 81.750000 ;
        RECT 63.410000 81.955000 63.610000 82.155000 ;
        RECT 63.410000 82.360000 63.610000 82.560000 ;
        RECT 63.660000 82.855000 63.860000 83.055000 ;
        RECT 63.660000 83.265000 63.860000 83.465000 ;
        RECT 63.660000 83.675000 63.860000 83.875000 ;
        RECT 63.660000 84.085000 63.860000 84.285000 ;
        RECT 63.660000 84.495000 63.860000 84.695000 ;
        RECT 63.660000 84.905000 63.860000 85.105000 ;
        RECT 63.660000 85.315000 63.860000 85.515000 ;
        RECT 63.660000 85.725000 63.860000 85.925000 ;
        RECT 63.660000 86.135000 63.860000 86.335000 ;
        RECT 63.660000 86.545000 63.860000 86.745000 ;
        RECT 63.660000 86.955000 63.860000 87.155000 ;
        RECT 63.660000 87.365000 63.860000 87.565000 ;
        RECT 63.660000 87.775000 63.860000 87.975000 ;
        RECT 63.660000 88.185000 63.860000 88.385000 ;
        RECT 63.660000 88.595000 63.860000 88.795000 ;
        RECT 63.660000 89.005000 63.860000 89.205000 ;
        RECT 63.660000 89.415000 63.860000 89.615000 ;
        RECT 63.660000 89.825000 63.860000 90.025000 ;
        RECT 63.660000 90.235000 63.860000 90.435000 ;
        RECT 63.660000 90.645000 63.860000 90.845000 ;
        RECT 63.660000 91.055000 63.860000 91.255000 ;
        RECT 63.660000 91.465000 63.860000 91.665000 ;
        RECT 63.660000 91.875000 63.860000 92.075000 ;
        RECT 63.660000 92.285000 63.860000 92.485000 ;
        RECT 63.660000 92.695000 63.860000 92.895000 ;
        RECT 63.805000 17.860000 64.005000 18.060000 ;
        RECT 63.805000 18.290000 64.005000 18.490000 ;
        RECT 63.805000 18.720000 64.005000 18.920000 ;
        RECT 63.805000 19.150000 64.005000 19.350000 ;
        RECT 63.805000 19.580000 64.005000 19.780000 ;
        RECT 63.805000 20.010000 64.005000 20.210000 ;
        RECT 63.805000 20.440000 64.005000 20.640000 ;
        RECT 63.805000 20.870000 64.005000 21.070000 ;
        RECT 63.805000 21.300000 64.005000 21.500000 ;
        RECT 63.805000 21.730000 64.005000 21.930000 ;
        RECT 63.805000 22.160000 64.005000 22.360000 ;
        RECT 63.810000 68.125000 64.010000 68.325000 ;
        RECT 63.810000 68.535000 64.010000 68.735000 ;
        RECT 63.810000 68.945000 64.010000 69.145000 ;
        RECT 63.810000 69.355000 64.010000 69.555000 ;
        RECT 63.810000 69.765000 64.010000 69.965000 ;
        RECT 63.810000 70.175000 64.010000 70.375000 ;
        RECT 63.810000 70.585000 64.010000 70.785000 ;
        RECT 63.810000 70.995000 64.010000 71.195000 ;
        RECT 63.810000 71.405000 64.010000 71.605000 ;
        RECT 63.810000 71.815000 64.010000 72.015000 ;
        RECT 63.810000 72.225000 64.010000 72.425000 ;
        RECT 63.810000 72.635000 64.010000 72.835000 ;
        RECT 63.810000 73.045000 64.010000 73.245000 ;
        RECT 63.810000 73.450000 64.010000 73.650000 ;
        RECT 63.810000 73.855000 64.010000 74.055000 ;
        RECT 63.810000 74.260000 64.010000 74.460000 ;
        RECT 63.810000 74.665000 64.010000 74.865000 ;
        RECT 63.810000 75.070000 64.010000 75.270000 ;
        RECT 63.810000 75.475000 64.010000 75.675000 ;
        RECT 63.810000 75.880000 64.010000 76.080000 ;
        RECT 63.810000 76.285000 64.010000 76.485000 ;
        RECT 63.810000 76.690000 64.010000 76.890000 ;
        RECT 63.810000 77.095000 64.010000 77.295000 ;
        RECT 63.810000 77.500000 64.010000 77.700000 ;
        RECT 63.810000 77.905000 64.010000 78.105000 ;
        RECT 63.810000 78.310000 64.010000 78.510000 ;
        RECT 63.810000 78.715000 64.010000 78.915000 ;
        RECT 63.810000 79.120000 64.010000 79.320000 ;
        RECT 63.810000 79.525000 64.010000 79.725000 ;
        RECT 63.810000 79.930000 64.010000 80.130000 ;
        RECT 63.810000 80.335000 64.010000 80.535000 ;
        RECT 63.810000 80.740000 64.010000 80.940000 ;
        RECT 63.810000 81.145000 64.010000 81.345000 ;
        RECT 63.810000 81.550000 64.010000 81.750000 ;
        RECT 63.810000 81.955000 64.010000 82.155000 ;
        RECT 63.810000 82.360000 64.010000 82.560000 ;
        RECT 64.070000 82.855000 64.270000 83.055000 ;
        RECT 64.070000 83.265000 64.270000 83.465000 ;
        RECT 64.070000 83.675000 64.270000 83.875000 ;
        RECT 64.070000 84.085000 64.270000 84.285000 ;
        RECT 64.070000 84.495000 64.270000 84.695000 ;
        RECT 64.070000 84.905000 64.270000 85.105000 ;
        RECT 64.070000 85.315000 64.270000 85.515000 ;
        RECT 64.070000 85.725000 64.270000 85.925000 ;
        RECT 64.070000 86.135000 64.270000 86.335000 ;
        RECT 64.070000 86.545000 64.270000 86.745000 ;
        RECT 64.070000 86.955000 64.270000 87.155000 ;
        RECT 64.070000 87.365000 64.270000 87.565000 ;
        RECT 64.070000 87.775000 64.270000 87.975000 ;
        RECT 64.070000 88.185000 64.270000 88.385000 ;
        RECT 64.070000 88.595000 64.270000 88.795000 ;
        RECT 64.070000 89.005000 64.270000 89.205000 ;
        RECT 64.070000 89.415000 64.270000 89.615000 ;
        RECT 64.070000 89.825000 64.270000 90.025000 ;
        RECT 64.070000 90.235000 64.270000 90.435000 ;
        RECT 64.070000 90.645000 64.270000 90.845000 ;
        RECT 64.070000 91.055000 64.270000 91.255000 ;
        RECT 64.070000 91.465000 64.270000 91.665000 ;
        RECT 64.070000 91.875000 64.270000 92.075000 ;
        RECT 64.070000 92.285000 64.270000 92.485000 ;
        RECT 64.070000 92.695000 64.270000 92.895000 ;
        RECT 64.210000 17.860000 64.410000 18.060000 ;
        RECT 64.210000 18.290000 64.410000 18.490000 ;
        RECT 64.210000 18.720000 64.410000 18.920000 ;
        RECT 64.210000 19.150000 64.410000 19.350000 ;
        RECT 64.210000 19.580000 64.410000 19.780000 ;
        RECT 64.210000 20.010000 64.410000 20.210000 ;
        RECT 64.210000 20.440000 64.410000 20.640000 ;
        RECT 64.210000 20.870000 64.410000 21.070000 ;
        RECT 64.210000 21.300000 64.410000 21.500000 ;
        RECT 64.210000 21.730000 64.410000 21.930000 ;
        RECT 64.210000 22.160000 64.410000 22.360000 ;
        RECT 64.210000 68.125000 64.410000 68.325000 ;
        RECT 64.210000 68.535000 64.410000 68.735000 ;
        RECT 64.210000 68.945000 64.410000 69.145000 ;
        RECT 64.210000 69.355000 64.410000 69.555000 ;
        RECT 64.210000 69.765000 64.410000 69.965000 ;
        RECT 64.210000 70.175000 64.410000 70.375000 ;
        RECT 64.210000 70.585000 64.410000 70.785000 ;
        RECT 64.210000 70.995000 64.410000 71.195000 ;
        RECT 64.210000 71.405000 64.410000 71.605000 ;
        RECT 64.210000 71.815000 64.410000 72.015000 ;
        RECT 64.210000 72.225000 64.410000 72.425000 ;
        RECT 64.210000 72.635000 64.410000 72.835000 ;
        RECT 64.210000 73.045000 64.410000 73.245000 ;
        RECT 64.210000 73.450000 64.410000 73.650000 ;
        RECT 64.210000 73.855000 64.410000 74.055000 ;
        RECT 64.210000 74.260000 64.410000 74.460000 ;
        RECT 64.210000 74.665000 64.410000 74.865000 ;
        RECT 64.210000 75.070000 64.410000 75.270000 ;
        RECT 64.210000 75.475000 64.410000 75.675000 ;
        RECT 64.210000 75.880000 64.410000 76.080000 ;
        RECT 64.210000 76.285000 64.410000 76.485000 ;
        RECT 64.210000 76.690000 64.410000 76.890000 ;
        RECT 64.210000 77.095000 64.410000 77.295000 ;
        RECT 64.210000 77.500000 64.410000 77.700000 ;
        RECT 64.210000 77.905000 64.410000 78.105000 ;
        RECT 64.210000 78.310000 64.410000 78.510000 ;
        RECT 64.210000 78.715000 64.410000 78.915000 ;
        RECT 64.210000 79.120000 64.410000 79.320000 ;
        RECT 64.210000 79.525000 64.410000 79.725000 ;
        RECT 64.210000 79.930000 64.410000 80.130000 ;
        RECT 64.210000 80.335000 64.410000 80.535000 ;
        RECT 64.210000 80.740000 64.410000 80.940000 ;
        RECT 64.210000 81.145000 64.410000 81.345000 ;
        RECT 64.210000 81.550000 64.410000 81.750000 ;
        RECT 64.210000 81.955000 64.410000 82.155000 ;
        RECT 64.210000 82.360000 64.410000 82.560000 ;
        RECT 64.480000 82.855000 64.680000 83.055000 ;
        RECT 64.480000 83.265000 64.680000 83.465000 ;
        RECT 64.480000 83.675000 64.680000 83.875000 ;
        RECT 64.480000 84.085000 64.680000 84.285000 ;
        RECT 64.480000 84.495000 64.680000 84.695000 ;
        RECT 64.480000 84.905000 64.680000 85.105000 ;
        RECT 64.480000 85.315000 64.680000 85.515000 ;
        RECT 64.480000 85.725000 64.680000 85.925000 ;
        RECT 64.480000 86.135000 64.680000 86.335000 ;
        RECT 64.480000 86.545000 64.680000 86.745000 ;
        RECT 64.480000 86.955000 64.680000 87.155000 ;
        RECT 64.480000 87.365000 64.680000 87.565000 ;
        RECT 64.480000 87.775000 64.680000 87.975000 ;
        RECT 64.480000 88.185000 64.680000 88.385000 ;
        RECT 64.480000 88.595000 64.680000 88.795000 ;
        RECT 64.480000 89.005000 64.680000 89.205000 ;
        RECT 64.480000 89.415000 64.680000 89.615000 ;
        RECT 64.480000 89.825000 64.680000 90.025000 ;
        RECT 64.480000 90.235000 64.680000 90.435000 ;
        RECT 64.480000 90.645000 64.680000 90.845000 ;
        RECT 64.480000 91.055000 64.680000 91.255000 ;
        RECT 64.480000 91.465000 64.680000 91.665000 ;
        RECT 64.480000 91.875000 64.680000 92.075000 ;
        RECT 64.480000 92.285000 64.680000 92.485000 ;
        RECT 64.480000 92.695000 64.680000 92.895000 ;
        RECT 64.610000 68.125000 64.810000 68.325000 ;
        RECT 64.610000 68.535000 64.810000 68.735000 ;
        RECT 64.610000 68.945000 64.810000 69.145000 ;
        RECT 64.610000 69.355000 64.810000 69.555000 ;
        RECT 64.610000 69.765000 64.810000 69.965000 ;
        RECT 64.610000 70.175000 64.810000 70.375000 ;
        RECT 64.610000 70.585000 64.810000 70.785000 ;
        RECT 64.610000 70.995000 64.810000 71.195000 ;
        RECT 64.610000 71.405000 64.810000 71.605000 ;
        RECT 64.610000 71.815000 64.810000 72.015000 ;
        RECT 64.610000 72.225000 64.810000 72.425000 ;
        RECT 64.610000 72.635000 64.810000 72.835000 ;
        RECT 64.610000 73.045000 64.810000 73.245000 ;
        RECT 64.610000 73.450000 64.810000 73.650000 ;
        RECT 64.610000 73.855000 64.810000 74.055000 ;
        RECT 64.610000 74.260000 64.810000 74.460000 ;
        RECT 64.610000 74.665000 64.810000 74.865000 ;
        RECT 64.610000 75.070000 64.810000 75.270000 ;
        RECT 64.610000 75.475000 64.810000 75.675000 ;
        RECT 64.610000 75.880000 64.810000 76.080000 ;
        RECT 64.610000 76.285000 64.810000 76.485000 ;
        RECT 64.610000 76.690000 64.810000 76.890000 ;
        RECT 64.610000 77.095000 64.810000 77.295000 ;
        RECT 64.610000 77.500000 64.810000 77.700000 ;
        RECT 64.610000 77.905000 64.810000 78.105000 ;
        RECT 64.610000 78.310000 64.810000 78.510000 ;
        RECT 64.610000 78.715000 64.810000 78.915000 ;
        RECT 64.610000 79.120000 64.810000 79.320000 ;
        RECT 64.610000 79.525000 64.810000 79.725000 ;
        RECT 64.610000 79.930000 64.810000 80.130000 ;
        RECT 64.610000 80.335000 64.810000 80.535000 ;
        RECT 64.610000 80.740000 64.810000 80.940000 ;
        RECT 64.610000 81.145000 64.810000 81.345000 ;
        RECT 64.610000 81.550000 64.810000 81.750000 ;
        RECT 64.610000 81.955000 64.810000 82.155000 ;
        RECT 64.610000 82.360000 64.810000 82.560000 ;
        RECT 64.615000 17.860000 64.815000 18.060000 ;
        RECT 64.615000 18.290000 64.815000 18.490000 ;
        RECT 64.615000 18.720000 64.815000 18.920000 ;
        RECT 64.615000 19.150000 64.815000 19.350000 ;
        RECT 64.615000 19.580000 64.815000 19.780000 ;
        RECT 64.615000 20.010000 64.815000 20.210000 ;
        RECT 64.615000 20.440000 64.815000 20.640000 ;
        RECT 64.615000 20.870000 64.815000 21.070000 ;
        RECT 64.615000 21.300000 64.815000 21.500000 ;
        RECT 64.615000 21.730000 64.815000 21.930000 ;
        RECT 64.615000 22.160000 64.815000 22.360000 ;
        RECT 64.890000 82.855000 65.090000 83.055000 ;
        RECT 64.890000 83.265000 65.090000 83.465000 ;
        RECT 64.890000 83.675000 65.090000 83.875000 ;
        RECT 64.890000 84.085000 65.090000 84.285000 ;
        RECT 64.890000 84.495000 65.090000 84.695000 ;
        RECT 64.890000 84.905000 65.090000 85.105000 ;
        RECT 64.890000 85.315000 65.090000 85.515000 ;
        RECT 64.890000 85.725000 65.090000 85.925000 ;
        RECT 64.890000 86.135000 65.090000 86.335000 ;
        RECT 64.890000 86.545000 65.090000 86.745000 ;
        RECT 64.890000 86.955000 65.090000 87.155000 ;
        RECT 64.890000 87.365000 65.090000 87.565000 ;
        RECT 64.890000 87.775000 65.090000 87.975000 ;
        RECT 64.890000 88.185000 65.090000 88.385000 ;
        RECT 64.890000 88.595000 65.090000 88.795000 ;
        RECT 64.890000 89.005000 65.090000 89.205000 ;
        RECT 64.890000 89.415000 65.090000 89.615000 ;
        RECT 64.890000 89.825000 65.090000 90.025000 ;
        RECT 64.890000 90.235000 65.090000 90.435000 ;
        RECT 64.890000 90.645000 65.090000 90.845000 ;
        RECT 64.890000 91.055000 65.090000 91.255000 ;
        RECT 64.890000 91.465000 65.090000 91.665000 ;
        RECT 64.890000 91.875000 65.090000 92.075000 ;
        RECT 64.890000 92.285000 65.090000 92.485000 ;
        RECT 64.890000 92.695000 65.090000 92.895000 ;
        RECT 65.010000 68.125000 65.210000 68.325000 ;
        RECT 65.010000 68.535000 65.210000 68.735000 ;
        RECT 65.010000 68.945000 65.210000 69.145000 ;
        RECT 65.010000 69.355000 65.210000 69.555000 ;
        RECT 65.010000 69.765000 65.210000 69.965000 ;
        RECT 65.010000 70.175000 65.210000 70.375000 ;
        RECT 65.010000 70.585000 65.210000 70.785000 ;
        RECT 65.010000 70.995000 65.210000 71.195000 ;
        RECT 65.010000 71.405000 65.210000 71.605000 ;
        RECT 65.010000 71.815000 65.210000 72.015000 ;
        RECT 65.010000 72.225000 65.210000 72.425000 ;
        RECT 65.010000 72.635000 65.210000 72.835000 ;
        RECT 65.010000 73.045000 65.210000 73.245000 ;
        RECT 65.010000 73.450000 65.210000 73.650000 ;
        RECT 65.010000 73.855000 65.210000 74.055000 ;
        RECT 65.010000 74.260000 65.210000 74.460000 ;
        RECT 65.010000 74.665000 65.210000 74.865000 ;
        RECT 65.010000 75.070000 65.210000 75.270000 ;
        RECT 65.010000 75.475000 65.210000 75.675000 ;
        RECT 65.010000 75.880000 65.210000 76.080000 ;
        RECT 65.010000 76.285000 65.210000 76.485000 ;
        RECT 65.010000 76.690000 65.210000 76.890000 ;
        RECT 65.010000 77.095000 65.210000 77.295000 ;
        RECT 65.010000 77.500000 65.210000 77.700000 ;
        RECT 65.010000 77.905000 65.210000 78.105000 ;
        RECT 65.010000 78.310000 65.210000 78.510000 ;
        RECT 65.010000 78.715000 65.210000 78.915000 ;
        RECT 65.010000 79.120000 65.210000 79.320000 ;
        RECT 65.010000 79.525000 65.210000 79.725000 ;
        RECT 65.010000 79.930000 65.210000 80.130000 ;
        RECT 65.010000 80.335000 65.210000 80.535000 ;
        RECT 65.010000 80.740000 65.210000 80.940000 ;
        RECT 65.010000 81.145000 65.210000 81.345000 ;
        RECT 65.010000 81.550000 65.210000 81.750000 ;
        RECT 65.010000 81.955000 65.210000 82.155000 ;
        RECT 65.010000 82.360000 65.210000 82.560000 ;
        RECT 65.020000 17.860000 65.220000 18.060000 ;
        RECT 65.020000 18.290000 65.220000 18.490000 ;
        RECT 65.020000 18.720000 65.220000 18.920000 ;
        RECT 65.020000 19.150000 65.220000 19.350000 ;
        RECT 65.020000 19.580000 65.220000 19.780000 ;
        RECT 65.020000 20.010000 65.220000 20.210000 ;
        RECT 65.020000 20.440000 65.220000 20.640000 ;
        RECT 65.020000 20.870000 65.220000 21.070000 ;
        RECT 65.020000 21.300000 65.220000 21.500000 ;
        RECT 65.020000 21.730000 65.220000 21.930000 ;
        RECT 65.020000 22.160000 65.220000 22.360000 ;
        RECT 65.300000 82.855000 65.500000 83.055000 ;
        RECT 65.300000 83.265000 65.500000 83.465000 ;
        RECT 65.300000 83.675000 65.500000 83.875000 ;
        RECT 65.300000 84.085000 65.500000 84.285000 ;
        RECT 65.300000 84.495000 65.500000 84.695000 ;
        RECT 65.300000 84.905000 65.500000 85.105000 ;
        RECT 65.300000 85.315000 65.500000 85.515000 ;
        RECT 65.300000 85.725000 65.500000 85.925000 ;
        RECT 65.300000 86.135000 65.500000 86.335000 ;
        RECT 65.300000 86.545000 65.500000 86.745000 ;
        RECT 65.300000 86.955000 65.500000 87.155000 ;
        RECT 65.300000 87.365000 65.500000 87.565000 ;
        RECT 65.300000 87.775000 65.500000 87.975000 ;
        RECT 65.300000 88.185000 65.500000 88.385000 ;
        RECT 65.300000 88.595000 65.500000 88.795000 ;
        RECT 65.300000 89.005000 65.500000 89.205000 ;
        RECT 65.300000 89.415000 65.500000 89.615000 ;
        RECT 65.300000 89.825000 65.500000 90.025000 ;
        RECT 65.300000 90.235000 65.500000 90.435000 ;
        RECT 65.300000 90.645000 65.500000 90.845000 ;
        RECT 65.300000 91.055000 65.500000 91.255000 ;
        RECT 65.300000 91.465000 65.500000 91.665000 ;
        RECT 65.300000 91.875000 65.500000 92.075000 ;
        RECT 65.300000 92.285000 65.500000 92.485000 ;
        RECT 65.300000 92.695000 65.500000 92.895000 ;
        RECT 65.410000 68.125000 65.610000 68.325000 ;
        RECT 65.410000 68.535000 65.610000 68.735000 ;
        RECT 65.410000 68.945000 65.610000 69.145000 ;
        RECT 65.410000 69.355000 65.610000 69.555000 ;
        RECT 65.410000 69.765000 65.610000 69.965000 ;
        RECT 65.410000 70.175000 65.610000 70.375000 ;
        RECT 65.410000 70.585000 65.610000 70.785000 ;
        RECT 65.410000 70.995000 65.610000 71.195000 ;
        RECT 65.410000 71.405000 65.610000 71.605000 ;
        RECT 65.410000 71.815000 65.610000 72.015000 ;
        RECT 65.410000 72.225000 65.610000 72.425000 ;
        RECT 65.410000 72.635000 65.610000 72.835000 ;
        RECT 65.410000 73.045000 65.610000 73.245000 ;
        RECT 65.410000 73.450000 65.610000 73.650000 ;
        RECT 65.410000 73.855000 65.610000 74.055000 ;
        RECT 65.410000 74.260000 65.610000 74.460000 ;
        RECT 65.410000 74.665000 65.610000 74.865000 ;
        RECT 65.410000 75.070000 65.610000 75.270000 ;
        RECT 65.410000 75.475000 65.610000 75.675000 ;
        RECT 65.410000 75.880000 65.610000 76.080000 ;
        RECT 65.410000 76.285000 65.610000 76.485000 ;
        RECT 65.410000 76.690000 65.610000 76.890000 ;
        RECT 65.410000 77.095000 65.610000 77.295000 ;
        RECT 65.410000 77.500000 65.610000 77.700000 ;
        RECT 65.410000 77.905000 65.610000 78.105000 ;
        RECT 65.410000 78.310000 65.610000 78.510000 ;
        RECT 65.410000 78.715000 65.610000 78.915000 ;
        RECT 65.410000 79.120000 65.610000 79.320000 ;
        RECT 65.410000 79.525000 65.610000 79.725000 ;
        RECT 65.410000 79.930000 65.610000 80.130000 ;
        RECT 65.410000 80.335000 65.610000 80.535000 ;
        RECT 65.410000 80.740000 65.610000 80.940000 ;
        RECT 65.410000 81.145000 65.610000 81.345000 ;
        RECT 65.410000 81.550000 65.610000 81.750000 ;
        RECT 65.410000 81.955000 65.610000 82.155000 ;
        RECT 65.410000 82.360000 65.610000 82.560000 ;
        RECT 65.425000 17.860000 65.625000 18.060000 ;
        RECT 65.425000 18.290000 65.625000 18.490000 ;
        RECT 65.425000 18.720000 65.625000 18.920000 ;
        RECT 65.425000 19.150000 65.625000 19.350000 ;
        RECT 65.425000 19.580000 65.625000 19.780000 ;
        RECT 65.425000 20.010000 65.625000 20.210000 ;
        RECT 65.425000 20.440000 65.625000 20.640000 ;
        RECT 65.425000 20.870000 65.625000 21.070000 ;
        RECT 65.425000 21.300000 65.625000 21.500000 ;
        RECT 65.425000 21.730000 65.625000 21.930000 ;
        RECT 65.425000 22.160000 65.625000 22.360000 ;
        RECT 65.710000 82.855000 65.910000 83.055000 ;
        RECT 65.710000 83.265000 65.910000 83.465000 ;
        RECT 65.710000 83.675000 65.910000 83.875000 ;
        RECT 65.710000 84.085000 65.910000 84.285000 ;
        RECT 65.710000 84.495000 65.910000 84.695000 ;
        RECT 65.710000 84.905000 65.910000 85.105000 ;
        RECT 65.710000 85.315000 65.910000 85.515000 ;
        RECT 65.710000 85.725000 65.910000 85.925000 ;
        RECT 65.710000 86.135000 65.910000 86.335000 ;
        RECT 65.710000 86.545000 65.910000 86.745000 ;
        RECT 65.710000 86.955000 65.910000 87.155000 ;
        RECT 65.710000 87.365000 65.910000 87.565000 ;
        RECT 65.710000 87.775000 65.910000 87.975000 ;
        RECT 65.710000 88.185000 65.910000 88.385000 ;
        RECT 65.710000 88.595000 65.910000 88.795000 ;
        RECT 65.710000 89.005000 65.910000 89.205000 ;
        RECT 65.710000 89.415000 65.910000 89.615000 ;
        RECT 65.710000 89.825000 65.910000 90.025000 ;
        RECT 65.710000 90.235000 65.910000 90.435000 ;
        RECT 65.710000 90.645000 65.910000 90.845000 ;
        RECT 65.710000 91.055000 65.910000 91.255000 ;
        RECT 65.710000 91.465000 65.910000 91.665000 ;
        RECT 65.710000 91.875000 65.910000 92.075000 ;
        RECT 65.710000 92.285000 65.910000 92.485000 ;
        RECT 65.710000 92.695000 65.910000 92.895000 ;
        RECT 65.810000 68.125000 66.010000 68.325000 ;
        RECT 65.810000 68.535000 66.010000 68.735000 ;
        RECT 65.810000 68.945000 66.010000 69.145000 ;
        RECT 65.810000 69.355000 66.010000 69.555000 ;
        RECT 65.810000 69.765000 66.010000 69.965000 ;
        RECT 65.810000 70.175000 66.010000 70.375000 ;
        RECT 65.810000 70.585000 66.010000 70.785000 ;
        RECT 65.810000 70.995000 66.010000 71.195000 ;
        RECT 65.810000 71.405000 66.010000 71.605000 ;
        RECT 65.810000 71.815000 66.010000 72.015000 ;
        RECT 65.810000 72.225000 66.010000 72.425000 ;
        RECT 65.810000 72.635000 66.010000 72.835000 ;
        RECT 65.810000 73.045000 66.010000 73.245000 ;
        RECT 65.810000 73.450000 66.010000 73.650000 ;
        RECT 65.810000 73.855000 66.010000 74.055000 ;
        RECT 65.810000 74.260000 66.010000 74.460000 ;
        RECT 65.810000 74.665000 66.010000 74.865000 ;
        RECT 65.810000 75.070000 66.010000 75.270000 ;
        RECT 65.810000 75.475000 66.010000 75.675000 ;
        RECT 65.810000 75.880000 66.010000 76.080000 ;
        RECT 65.810000 76.285000 66.010000 76.485000 ;
        RECT 65.810000 76.690000 66.010000 76.890000 ;
        RECT 65.810000 77.095000 66.010000 77.295000 ;
        RECT 65.810000 77.500000 66.010000 77.700000 ;
        RECT 65.810000 77.905000 66.010000 78.105000 ;
        RECT 65.810000 78.310000 66.010000 78.510000 ;
        RECT 65.810000 78.715000 66.010000 78.915000 ;
        RECT 65.810000 79.120000 66.010000 79.320000 ;
        RECT 65.810000 79.525000 66.010000 79.725000 ;
        RECT 65.810000 79.930000 66.010000 80.130000 ;
        RECT 65.810000 80.335000 66.010000 80.535000 ;
        RECT 65.810000 80.740000 66.010000 80.940000 ;
        RECT 65.810000 81.145000 66.010000 81.345000 ;
        RECT 65.810000 81.550000 66.010000 81.750000 ;
        RECT 65.810000 81.955000 66.010000 82.155000 ;
        RECT 65.810000 82.360000 66.010000 82.560000 ;
        RECT 65.830000 17.860000 66.030000 18.060000 ;
        RECT 65.830000 18.290000 66.030000 18.490000 ;
        RECT 65.830000 18.720000 66.030000 18.920000 ;
        RECT 65.830000 19.150000 66.030000 19.350000 ;
        RECT 65.830000 19.580000 66.030000 19.780000 ;
        RECT 65.830000 20.010000 66.030000 20.210000 ;
        RECT 65.830000 20.440000 66.030000 20.640000 ;
        RECT 65.830000 20.870000 66.030000 21.070000 ;
        RECT 65.830000 21.300000 66.030000 21.500000 ;
        RECT 65.830000 21.730000 66.030000 21.930000 ;
        RECT 65.830000 22.160000 66.030000 22.360000 ;
        RECT 66.120000 82.855000 66.320000 83.055000 ;
        RECT 66.120000 83.265000 66.320000 83.465000 ;
        RECT 66.120000 83.675000 66.320000 83.875000 ;
        RECT 66.120000 84.085000 66.320000 84.285000 ;
        RECT 66.120000 84.495000 66.320000 84.695000 ;
        RECT 66.120000 84.905000 66.320000 85.105000 ;
        RECT 66.120000 85.315000 66.320000 85.515000 ;
        RECT 66.120000 85.725000 66.320000 85.925000 ;
        RECT 66.120000 86.135000 66.320000 86.335000 ;
        RECT 66.120000 86.545000 66.320000 86.745000 ;
        RECT 66.120000 86.955000 66.320000 87.155000 ;
        RECT 66.120000 87.365000 66.320000 87.565000 ;
        RECT 66.120000 87.775000 66.320000 87.975000 ;
        RECT 66.120000 88.185000 66.320000 88.385000 ;
        RECT 66.120000 88.595000 66.320000 88.795000 ;
        RECT 66.120000 89.005000 66.320000 89.205000 ;
        RECT 66.120000 89.415000 66.320000 89.615000 ;
        RECT 66.120000 89.825000 66.320000 90.025000 ;
        RECT 66.120000 90.235000 66.320000 90.435000 ;
        RECT 66.120000 90.645000 66.320000 90.845000 ;
        RECT 66.120000 91.055000 66.320000 91.255000 ;
        RECT 66.120000 91.465000 66.320000 91.665000 ;
        RECT 66.120000 91.875000 66.320000 92.075000 ;
        RECT 66.120000 92.285000 66.320000 92.485000 ;
        RECT 66.120000 92.695000 66.320000 92.895000 ;
        RECT 66.210000 68.125000 66.410000 68.325000 ;
        RECT 66.210000 68.535000 66.410000 68.735000 ;
        RECT 66.210000 68.945000 66.410000 69.145000 ;
        RECT 66.210000 69.355000 66.410000 69.555000 ;
        RECT 66.210000 69.765000 66.410000 69.965000 ;
        RECT 66.210000 70.175000 66.410000 70.375000 ;
        RECT 66.210000 70.585000 66.410000 70.785000 ;
        RECT 66.210000 70.995000 66.410000 71.195000 ;
        RECT 66.210000 71.405000 66.410000 71.605000 ;
        RECT 66.210000 71.815000 66.410000 72.015000 ;
        RECT 66.210000 72.225000 66.410000 72.425000 ;
        RECT 66.210000 72.635000 66.410000 72.835000 ;
        RECT 66.210000 73.045000 66.410000 73.245000 ;
        RECT 66.210000 73.450000 66.410000 73.650000 ;
        RECT 66.210000 73.855000 66.410000 74.055000 ;
        RECT 66.210000 74.260000 66.410000 74.460000 ;
        RECT 66.210000 74.665000 66.410000 74.865000 ;
        RECT 66.210000 75.070000 66.410000 75.270000 ;
        RECT 66.210000 75.475000 66.410000 75.675000 ;
        RECT 66.210000 75.880000 66.410000 76.080000 ;
        RECT 66.210000 76.285000 66.410000 76.485000 ;
        RECT 66.210000 76.690000 66.410000 76.890000 ;
        RECT 66.210000 77.095000 66.410000 77.295000 ;
        RECT 66.210000 77.500000 66.410000 77.700000 ;
        RECT 66.210000 77.905000 66.410000 78.105000 ;
        RECT 66.210000 78.310000 66.410000 78.510000 ;
        RECT 66.210000 78.715000 66.410000 78.915000 ;
        RECT 66.210000 79.120000 66.410000 79.320000 ;
        RECT 66.210000 79.525000 66.410000 79.725000 ;
        RECT 66.210000 79.930000 66.410000 80.130000 ;
        RECT 66.210000 80.335000 66.410000 80.535000 ;
        RECT 66.210000 80.740000 66.410000 80.940000 ;
        RECT 66.210000 81.145000 66.410000 81.345000 ;
        RECT 66.210000 81.550000 66.410000 81.750000 ;
        RECT 66.210000 81.955000 66.410000 82.155000 ;
        RECT 66.210000 82.360000 66.410000 82.560000 ;
        RECT 66.235000 17.860000 66.435000 18.060000 ;
        RECT 66.235000 18.290000 66.435000 18.490000 ;
        RECT 66.235000 18.720000 66.435000 18.920000 ;
        RECT 66.235000 19.150000 66.435000 19.350000 ;
        RECT 66.235000 19.580000 66.435000 19.780000 ;
        RECT 66.235000 20.010000 66.435000 20.210000 ;
        RECT 66.235000 20.440000 66.435000 20.640000 ;
        RECT 66.235000 20.870000 66.435000 21.070000 ;
        RECT 66.235000 21.300000 66.435000 21.500000 ;
        RECT 66.235000 21.730000 66.435000 21.930000 ;
        RECT 66.235000 22.160000 66.435000 22.360000 ;
        RECT 66.530000 82.855000 66.730000 83.055000 ;
        RECT 66.530000 83.265000 66.730000 83.465000 ;
        RECT 66.530000 83.675000 66.730000 83.875000 ;
        RECT 66.530000 84.085000 66.730000 84.285000 ;
        RECT 66.530000 84.495000 66.730000 84.695000 ;
        RECT 66.530000 84.905000 66.730000 85.105000 ;
        RECT 66.530000 85.315000 66.730000 85.515000 ;
        RECT 66.530000 85.725000 66.730000 85.925000 ;
        RECT 66.530000 86.135000 66.730000 86.335000 ;
        RECT 66.530000 86.545000 66.730000 86.745000 ;
        RECT 66.530000 86.955000 66.730000 87.155000 ;
        RECT 66.530000 87.365000 66.730000 87.565000 ;
        RECT 66.530000 87.775000 66.730000 87.975000 ;
        RECT 66.530000 88.185000 66.730000 88.385000 ;
        RECT 66.530000 88.595000 66.730000 88.795000 ;
        RECT 66.530000 89.005000 66.730000 89.205000 ;
        RECT 66.530000 89.415000 66.730000 89.615000 ;
        RECT 66.530000 89.825000 66.730000 90.025000 ;
        RECT 66.530000 90.235000 66.730000 90.435000 ;
        RECT 66.530000 90.645000 66.730000 90.845000 ;
        RECT 66.530000 91.055000 66.730000 91.255000 ;
        RECT 66.530000 91.465000 66.730000 91.665000 ;
        RECT 66.530000 91.875000 66.730000 92.075000 ;
        RECT 66.530000 92.285000 66.730000 92.485000 ;
        RECT 66.530000 92.695000 66.730000 92.895000 ;
        RECT 66.610000 68.125000 66.810000 68.325000 ;
        RECT 66.610000 68.535000 66.810000 68.735000 ;
        RECT 66.610000 68.945000 66.810000 69.145000 ;
        RECT 66.610000 69.355000 66.810000 69.555000 ;
        RECT 66.610000 69.765000 66.810000 69.965000 ;
        RECT 66.610000 70.175000 66.810000 70.375000 ;
        RECT 66.610000 70.585000 66.810000 70.785000 ;
        RECT 66.610000 70.995000 66.810000 71.195000 ;
        RECT 66.610000 71.405000 66.810000 71.605000 ;
        RECT 66.610000 71.815000 66.810000 72.015000 ;
        RECT 66.610000 72.225000 66.810000 72.425000 ;
        RECT 66.610000 72.635000 66.810000 72.835000 ;
        RECT 66.610000 73.045000 66.810000 73.245000 ;
        RECT 66.610000 73.450000 66.810000 73.650000 ;
        RECT 66.610000 73.855000 66.810000 74.055000 ;
        RECT 66.610000 74.260000 66.810000 74.460000 ;
        RECT 66.610000 74.665000 66.810000 74.865000 ;
        RECT 66.610000 75.070000 66.810000 75.270000 ;
        RECT 66.610000 75.475000 66.810000 75.675000 ;
        RECT 66.610000 75.880000 66.810000 76.080000 ;
        RECT 66.610000 76.285000 66.810000 76.485000 ;
        RECT 66.610000 76.690000 66.810000 76.890000 ;
        RECT 66.610000 77.095000 66.810000 77.295000 ;
        RECT 66.610000 77.500000 66.810000 77.700000 ;
        RECT 66.610000 77.905000 66.810000 78.105000 ;
        RECT 66.610000 78.310000 66.810000 78.510000 ;
        RECT 66.610000 78.715000 66.810000 78.915000 ;
        RECT 66.610000 79.120000 66.810000 79.320000 ;
        RECT 66.610000 79.525000 66.810000 79.725000 ;
        RECT 66.610000 79.930000 66.810000 80.130000 ;
        RECT 66.610000 80.335000 66.810000 80.535000 ;
        RECT 66.610000 80.740000 66.810000 80.940000 ;
        RECT 66.610000 81.145000 66.810000 81.345000 ;
        RECT 66.610000 81.550000 66.810000 81.750000 ;
        RECT 66.610000 81.955000 66.810000 82.155000 ;
        RECT 66.610000 82.360000 66.810000 82.560000 ;
        RECT 66.640000 17.860000 66.840000 18.060000 ;
        RECT 66.640000 18.290000 66.840000 18.490000 ;
        RECT 66.640000 18.720000 66.840000 18.920000 ;
        RECT 66.640000 19.150000 66.840000 19.350000 ;
        RECT 66.640000 19.580000 66.840000 19.780000 ;
        RECT 66.640000 20.010000 66.840000 20.210000 ;
        RECT 66.640000 20.440000 66.840000 20.640000 ;
        RECT 66.640000 20.870000 66.840000 21.070000 ;
        RECT 66.640000 21.300000 66.840000 21.500000 ;
        RECT 66.640000 21.730000 66.840000 21.930000 ;
        RECT 66.640000 22.160000 66.840000 22.360000 ;
        RECT 66.940000 82.855000 67.140000 83.055000 ;
        RECT 66.940000 83.265000 67.140000 83.465000 ;
        RECT 66.940000 83.675000 67.140000 83.875000 ;
        RECT 66.940000 84.085000 67.140000 84.285000 ;
        RECT 66.940000 84.495000 67.140000 84.695000 ;
        RECT 66.940000 84.905000 67.140000 85.105000 ;
        RECT 66.940000 85.315000 67.140000 85.515000 ;
        RECT 66.940000 85.725000 67.140000 85.925000 ;
        RECT 66.940000 86.135000 67.140000 86.335000 ;
        RECT 66.940000 86.545000 67.140000 86.745000 ;
        RECT 66.940000 86.955000 67.140000 87.155000 ;
        RECT 66.940000 87.365000 67.140000 87.565000 ;
        RECT 66.940000 87.775000 67.140000 87.975000 ;
        RECT 66.940000 88.185000 67.140000 88.385000 ;
        RECT 66.940000 88.595000 67.140000 88.795000 ;
        RECT 66.940000 89.005000 67.140000 89.205000 ;
        RECT 66.940000 89.415000 67.140000 89.615000 ;
        RECT 66.940000 89.825000 67.140000 90.025000 ;
        RECT 66.940000 90.235000 67.140000 90.435000 ;
        RECT 66.940000 90.645000 67.140000 90.845000 ;
        RECT 66.940000 91.055000 67.140000 91.255000 ;
        RECT 66.940000 91.465000 67.140000 91.665000 ;
        RECT 66.940000 91.875000 67.140000 92.075000 ;
        RECT 66.940000 92.285000 67.140000 92.485000 ;
        RECT 66.940000 92.695000 67.140000 92.895000 ;
        RECT 67.010000 68.125000 67.210000 68.325000 ;
        RECT 67.010000 68.535000 67.210000 68.735000 ;
        RECT 67.010000 68.945000 67.210000 69.145000 ;
        RECT 67.010000 69.355000 67.210000 69.555000 ;
        RECT 67.010000 69.765000 67.210000 69.965000 ;
        RECT 67.010000 70.175000 67.210000 70.375000 ;
        RECT 67.010000 70.585000 67.210000 70.785000 ;
        RECT 67.010000 70.995000 67.210000 71.195000 ;
        RECT 67.010000 71.405000 67.210000 71.605000 ;
        RECT 67.010000 71.815000 67.210000 72.015000 ;
        RECT 67.010000 72.225000 67.210000 72.425000 ;
        RECT 67.010000 72.635000 67.210000 72.835000 ;
        RECT 67.010000 73.045000 67.210000 73.245000 ;
        RECT 67.010000 73.450000 67.210000 73.650000 ;
        RECT 67.010000 73.855000 67.210000 74.055000 ;
        RECT 67.010000 74.260000 67.210000 74.460000 ;
        RECT 67.010000 74.665000 67.210000 74.865000 ;
        RECT 67.010000 75.070000 67.210000 75.270000 ;
        RECT 67.010000 75.475000 67.210000 75.675000 ;
        RECT 67.010000 75.880000 67.210000 76.080000 ;
        RECT 67.010000 76.285000 67.210000 76.485000 ;
        RECT 67.010000 76.690000 67.210000 76.890000 ;
        RECT 67.010000 77.095000 67.210000 77.295000 ;
        RECT 67.010000 77.500000 67.210000 77.700000 ;
        RECT 67.010000 77.905000 67.210000 78.105000 ;
        RECT 67.010000 78.310000 67.210000 78.510000 ;
        RECT 67.010000 78.715000 67.210000 78.915000 ;
        RECT 67.010000 79.120000 67.210000 79.320000 ;
        RECT 67.010000 79.525000 67.210000 79.725000 ;
        RECT 67.010000 79.930000 67.210000 80.130000 ;
        RECT 67.010000 80.335000 67.210000 80.535000 ;
        RECT 67.010000 80.740000 67.210000 80.940000 ;
        RECT 67.010000 81.145000 67.210000 81.345000 ;
        RECT 67.010000 81.550000 67.210000 81.750000 ;
        RECT 67.010000 81.955000 67.210000 82.155000 ;
        RECT 67.010000 82.360000 67.210000 82.560000 ;
        RECT 67.045000 17.860000 67.245000 18.060000 ;
        RECT 67.045000 18.290000 67.245000 18.490000 ;
        RECT 67.045000 18.720000 67.245000 18.920000 ;
        RECT 67.045000 19.150000 67.245000 19.350000 ;
        RECT 67.045000 19.580000 67.245000 19.780000 ;
        RECT 67.045000 20.010000 67.245000 20.210000 ;
        RECT 67.045000 20.440000 67.245000 20.640000 ;
        RECT 67.045000 20.870000 67.245000 21.070000 ;
        RECT 67.045000 21.300000 67.245000 21.500000 ;
        RECT 67.045000 21.730000 67.245000 21.930000 ;
        RECT 67.045000 22.160000 67.245000 22.360000 ;
        RECT 67.350000 82.855000 67.550000 83.055000 ;
        RECT 67.350000 83.265000 67.550000 83.465000 ;
        RECT 67.350000 83.675000 67.550000 83.875000 ;
        RECT 67.350000 84.085000 67.550000 84.285000 ;
        RECT 67.350000 84.495000 67.550000 84.695000 ;
        RECT 67.350000 84.905000 67.550000 85.105000 ;
        RECT 67.350000 85.315000 67.550000 85.515000 ;
        RECT 67.350000 85.725000 67.550000 85.925000 ;
        RECT 67.350000 86.135000 67.550000 86.335000 ;
        RECT 67.350000 86.545000 67.550000 86.745000 ;
        RECT 67.350000 86.955000 67.550000 87.155000 ;
        RECT 67.350000 87.365000 67.550000 87.565000 ;
        RECT 67.350000 87.775000 67.550000 87.975000 ;
        RECT 67.350000 88.185000 67.550000 88.385000 ;
        RECT 67.350000 88.595000 67.550000 88.795000 ;
        RECT 67.350000 89.005000 67.550000 89.205000 ;
        RECT 67.350000 89.415000 67.550000 89.615000 ;
        RECT 67.350000 89.825000 67.550000 90.025000 ;
        RECT 67.350000 90.235000 67.550000 90.435000 ;
        RECT 67.350000 90.645000 67.550000 90.845000 ;
        RECT 67.350000 91.055000 67.550000 91.255000 ;
        RECT 67.350000 91.465000 67.550000 91.665000 ;
        RECT 67.350000 91.875000 67.550000 92.075000 ;
        RECT 67.350000 92.285000 67.550000 92.485000 ;
        RECT 67.350000 92.695000 67.550000 92.895000 ;
        RECT 67.410000 68.125000 67.610000 68.325000 ;
        RECT 67.410000 68.535000 67.610000 68.735000 ;
        RECT 67.410000 68.945000 67.610000 69.145000 ;
        RECT 67.410000 69.355000 67.610000 69.555000 ;
        RECT 67.410000 69.765000 67.610000 69.965000 ;
        RECT 67.410000 70.175000 67.610000 70.375000 ;
        RECT 67.410000 70.585000 67.610000 70.785000 ;
        RECT 67.410000 70.995000 67.610000 71.195000 ;
        RECT 67.410000 71.405000 67.610000 71.605000 ;
        RECT 67.410000 71.815000 67.610000 72.015000 ;
        RECT 67.410000 72.225000 67.610000 72.425000 ;
        RECT 67.410000 72.635000 67.610000 72.835000 ;
        RECT 67.410000 73.045000 67.610000 73.245000 ;
        RECT 67.410000 73.450000 67.610000 73.650000 ;
        RECT 67.410000 73.855000 67.610000 74.055000 ;
        RECT 67.410000 74.260000 67.610000 74.460000 ;
        RECT 67.410000 74.665000 67.610000 74.865000 ;
        RECT 67.410000 75.070000 67.610000 75.270000 ;
        RECT 67.410000 75.475000 67.610000 75.675000 ;
        RECT 67.410000 75.880000 67.610000 76.080000 ;
        RECT 67.410000 76.285000 67.610000 76.485000 ;
        RECT 67.410000 76.690000 67.610000 76.890000 ;
        RECT 67.410000 77.095000 67.610000 77.295000 ;
        RECT 67.410000 77.500000 67.610000 77.700000 ;
        RECT 67.410000 77.905000 67.610000 78.105000 ;
        RECT 67.410000 78.310000 67.610000 78.510000 ;
        RECT 67.410000 78.715000 67.610000 78.915000 ;
        RECT 67.410000 79.120000 67.610000 79.320000 ;
        RECT 67.410000 79.525000 67.610000 79.725000 ;
        RECT 67.410000 79.930000 67.610000 80.130000 ;
        RECT 67.410000 80.335000 67.610000 80.535000 ;
        RECT 67.410000 80.740000 67.610000 80.940000 ;
        RECT 67.410000 81.145000 67.610000 81.345000 ;
        RECT 67.410000 81.550000 67.610000 81.750000 ;
        RECT 67.410000 81.955000 67.610000 82.155000 ;
        RECT 67.410000 82.360000 67.610000 82.560000 ;
        RECT 67.450000 17.860000 67.650000 18.060000 ;
        RECT 67.450000 18.290000 67.650000 18.490000 ;
        RECT 67.450000 18.720000 67.650000 18.920000 ;
        RECT 67.450000 19.150000 67.650000 19.350000 ;
        RECT 67.450000 19.580000 67.650000 19.780000 ;
        RECT 67.450000 20.010000 67.650000 20.210000 ;
        RECT 67.450000 20.440000 67.650000 20.640000 ;
        RECT 67.450000 20.870000 67.650000 21.070000 ;
        RECT 67.450000 21.300000 67.650000 21.500000 ;
        RECT 67.450000 21.730000 67.650000 21.930000 ;
        RECT 67.450000 22.160000 67.650000 22.360000 ;
        RECT 67.760000 82.855000 67.960000 83.055000 ;
        RECT 67.760000 83.265000 67.960000 83.465000 ;
        RECT 67.760000 83.675000 67.960000 83.875000 ;
        RECT 67.760000 84.085000 67.960000 84.285000 ;
        RECT 67.760000 84.495000 67.960000 84.695000 ;
        RECT 67.760000 84.905000 67.960000 85.105000 ;
        RECT 67.760000 85.315000 67.960000 85.515000 ;
        RECT 67.760000 85.725000 67.960000 85.925000 ;
        RECT 67.760000 86.135000 67.960000 86.335000 ;
        RECT 67.760000 86.545000 67.960000 86.745000 ;
        RECT 67.760000 86.955000 67.960000 87.155000 ;
        RECT 67.760000 87.365000 67.960000 87.565000 ;
        RECT 67.760000 87.775000 67.960000 87.975000 ;
        RECT 67.760000 88.185000 67.960000 88.385000 ;
        RECT 67.760000 88.595000 67.960000 88.795000 ;
        RECT 67.760000 89.005000 67.960000 89.205000 ;
        RECT 67.760000 89.415000 67.960000 89.615000 ;
        RECT 67.760000 89.825000 67.960000 90.025000 ;
        RECT 67.760000 90.235000 67.960000 90.435000 ;
        RECT 67.760000 90.645000 67.960000 90.845000 ;
        RECT 67.760000 91.055000 67.960000 91.255000 ;
        RECT 67.760000 91.465000 67.960000 91.665000 ;
        RECT 67.760000 91.875000 67.960000 92.075000 ;
        RECT 67.760000 92.285000 67.960000 92.485000 ;
        RECT 67.760000 92.695000 67.960000 92.895000 ;
        RECT 67.810000 68.125000 68.010000 68.325000 ;
        RECT 67.810000 68.535000 68.010000 68.735000 ;
        RECT 67.810000 68.945000 68.010000 69.145000 ;
        RECT 67.810000 69.355000 68.010000 69.555000 ;
        RECT 67.810000 69.765000 68.010000 69.965000 ;
        RECT 67.810000 70.175000 68.010000 70.375000 ;
        RECT 67.810000 70.585000 68.010000 70.785000 ;
        RECT 67.810000 70.995000 68.010000 71.195000 ;
        RECT 67.810000 71.405000 68.010000 71.605000 ;
        RECT 67.810000 71.815000 68.010000 72.015000 ;
        RECT 67.810000 72.225000 68.010000 72.425000 ;
        RECT 67.810000 72.635000 68.010000 72.835000 ;
        RECT 67.810000 73.045000 68.010000 73.245000 ;
        RECT 67.810000 73.450000 68.010000 73.650000 ;
        RECT 67.810000 73.855000 68.010000 74.055000 ;
        RECT 67.810000 74.260000 68.010000 74.460000 ;
        RECT 67.810000 74.665000 68.010000 74.865000 ;
        RECT 67.810000 75.070000 68.010000 75.270000 ;
        RECT 67.810000 75.475000 68.010000 75.675000 ;
        RECT 67.810000 75.880000 68.010000 76.080000 ;
        RECT 67.810000 76.285000 68.010000 76.485000 ;
        RECT 67.810000 76.690000 68.010000 76.890000 ;
        RECT 67.810000 77.095000 68.010000 77.295000 ;
        RECT 67.810000 77.500000 68.010000 77.700000 ;
        RECT 67.810000 77.905000 68.010000 78.105000 ;
        RECT 67.810000 78.310000 68.010000 78.510000 ;
        RECT 67.810000 78.715000 68.010000 78.915000 ;
        RECT 67.810000 79.120000 68.010000 79.320000 ;
        RECT 67.810000 79.525000 68.010000 79.725000 ;
        RECT 67.810000 79.930000 68.010000 80.130000 ;
        RECT 67.810000 80.335000 68.010000 80.535000 ;
        RECT 67.810000 80.740000 68.010000 80.940000 ;
        RECT 67.810000 81.145000 68.010000 81.345000 ;
        RECT 67.810000 81.550000 68.010000 81.750000 ;
        RECT 67.810000 81.955000 68.010000 82.155000 ;
        RECT 67.810000 82.360000 68.010000 82.560000 ;
        RECT 67.855000 17.860000 68.055000 18.060000 ;
        RECT 67.855000 18.290000 68.055000 18.490000 ;
        RECT 67.855000 18.720000 68.055000 18.920000 ;
        RECT 67.855000 19.150000 68.055000 19.350000 ;
        RECT 67.855000 19.580000 68.055000 19.780000 ;
        RECT 67.855000 20.010000 68.055000 20.210000 ;
        RECT 67.855000 20.440000 68.055000 20.640000 ;
        RECT 67.855000 20.870000 68.055000 21.070000 ;
        RECT 67.855000 21.300000 68.055000 21.500000 ;
        RECT 67.855000 21.730000 68.055000 21.930000 ;
        RECT 67.855000 22.160000 68.055000 22.360000 ;
        RECT 68.170000 82.855000 68.370000 83.055000 ;
        RECT 68.170000 83.265000 68.370000 83.465000 ;
        RECT 68.170000 83.675000 68.370000 83.875000 ;
        RECT 68.170000 84.085000 68.370000 84.285000 ;
        RECT 68.170000 84.495000 68.370000 84.695000 ;
        RECT 68.170000 84.905000 68.370000 85.105000 ;
        RECT 68.170000 85.315000 68.370000 85.515000 ;
        RECT 68.170000 85.725000 68.370000 85.925000 ;
        RECT 68.170000 86.135000 68.370000 86.335000 ;
        RECT 68.170000 86.545000 68.370000 86.745000 ;
        RECT 68.170000 86.955000 68.370000 87.155000 ;
        RECT 68.170000 87.365000 68.370000 87.565000 ;
        RECT 68.170000 87.775000 68.370000 87.975000 ;
        RECT 68.170000 88.185000 68.370000 88.385000 ;
        RECT 68.170000 88.595000 68.370000 88.795000 ;
        RECT 68.170000 89.005000 68.370000 89.205000 ;
        RECT 68.170000 89.415000 68.370000 89.615000 ;
        RECT 68.170000 89.825000 68.370000 90.025000 ;
        RECT 68.170000 90.235000 68.370000 90.435000 ;
        RECT 68.170000 90.645000 68.370000 90.845000 ;
        RECT 68.170000 91.055000 68.370000 91.255000 ;
        RECT 68.170000 91.465000 68.370000 91.665000 ;
        RECT 68.170000 91.875000 68.370000 92.075000 ;
        RECT 68.170000 92.285000 68.370000 92.485000 ;
        RECT 68.170000 92.695000 68.370000 92.895000 ;
        RECT 68.210000 68.125000 68.410000 68.325000 ;
        RECT 68.210000 68.535000 68.410000 68.735000 ;
        RECT 68.210000 68.945000 68.410000 69.145000 ;
        RECT 68.210000 69.355000 68.410000 69.555000 ;
        RECT 68.210000 69.765000 68.410000 69.965000 ;
        RECT 68.210000 70.175000 68.410000 70.375000 ;
        RECT 68.210000 70.585000 68.410000 70.785000 ;
        RECT 68.210000 70.995000 68.410000 71.195000 ;
        RECT 68.210000 71.405000 68.410000 71.605000 ;
        RECT 68.210000 71.815000 68.410000 72.015000 ;
        RECT 68.210000 72.225000 68.410000 72.425000 ;
        RECT 68.210000 72.635000 68.410000 72.835000 ;
        RECT 68.210000 73.045000 68.410000 73.245000 ;
        RECT 68.210000 73.450000 68.410000 73.650000 ;
        RECT 68.210000 73.855000 68.410000 74.055000 ;
        RECT 68.210000 74.260000 68.410000 74.460000 ;
        RECT 68.210000 74.665000 68.410000 74.865000 ;
        RECT 68.210000 75.070000 68.410000 75.270000 ;
        RECT 68.210000 75.475000 68.410000 75.675000 ;
        RECT 68.210000 75.880000 68.410000 76.080000 ;
        RECT 68.210000 76.285000 68.410000 76.485000 ;
        RECT 68.210000 76.690000 68.410000 76.890000 ;
        RECT 68.210000 77.095000 68.410000 77.295000 ;
        RECT 68.210000 77.500000 68.410000 77.700000 ;
        RECT 68.210000 77.905000 68.410000 78.105000 ;
        RECT 68.210000 78.310000 68.410000 78.510000 ;
        RECT 68.210000 78.715000 68.410000 78.915000 ;
        RECT 68.210000 79.120000 68.410000 79.320000 ;
        RECT 68.210000 79.525000 68.410000 79.725000 ;
        RECT 68.210000 79.930000 68.410000 80.130000 ;
        RECT 68.210000 80.335000 68.410000 80.535000 ;
        RECT 68.210000 80.740000 68.410000 80.940000 ;
        RECT 68.210000 81.145000 68.410000 81.345000 ;
        RECT 68.210000 81.550000 68.410000 81.750000 ;
        RECT 68.210000 81.955000 68.410000 82.155000 ;
        RECT 68.210000 82.360000 68.410000 82.560000 ;
        RECT 68.260000 17.860000 68.460000 18.060000 ;
        RECT 68.260000 18.290000 68.460000 18.490000 ;
        RECT 68.260000 18.720000 68.460000 18.920000 ;
        RECT 68.260000 19.150000 68.460000 19.350000 ;
        RECT 68.260000 19.580000 68.460000 19.780000 ;
        RECT 68.260000 20.010000 68.460000 20.210000 ;
        RECT 68.260000 20.440000 68.460000 20.640000 ;
        RECT 68.260000 20.870000 68.460000 21.070000 ;
        RECT 68.260000 21.300000 68.460000 21.500000 ;
        RECT 68.260000 21.730000 68.460000 21.930000 ;
        RECT 68.260000 22.160000 68.460000 22.360000 ;
        RECT 68.580000 82.855000 68.780000 83.055000 ;
        RECT 68.580000 83.265000 68.780000 83.465000 ;
        RECT 68.580000 83.675000 68.780000 83.875000 ;
        RECT 68.580000 84.085000 68.780000 84.285000 ;
        RECT 68.580000 84.495000 68.780000 84.695000 ;
        RECT 68.580000 84.905000 68.780000 85.105000 ;
        RECT 68.580000 85.315000 68.780000 85.515000 ;
        RECT 68.580000 85.725000 68.780000 85.925000 ;
        RECT 68.580000 86.135000 68.780000 86.335000 ;
        RECT 68.580000 86.545000 68.780000 86.745000 ;
        RECT 68.580000 86.955000 68.780000 87.155000 ;
        RECT 68.580000 87.365000 68.780000 87.565000 ;
        RECT 68.580000 87.775000 68.780000 87.975000 ;
        RECT 68.580000 88.185000 68.780000 88.385000 ;
        RECT 68.580000 88.595000 68.780000 88.795000 ;
        RECT 68.580000 89.005000 68.780000 89.205000 ;
        RECT 68.580000 89.415000 68.780000 89.615000 ;
        RECT 68.580000 89.825000 68.780000 90.025000 ;
        RECT 68.580000 90.235000 68.780000 90.435000 ;
        RECT 68.580000 90.645000 68.780000 90.845000 ;
        RECT 68.580000 91.055000 68.780000 91.255000 ;
        RECT 68.580000 91.465000 68.780000 91.665000 ;
        RECT 68.580000 91.875000 68.780000 92.075000 ;
        RECT 68.580000 92.285000 68.780000 92.485000 ;
        RECT 68.580000 92.695000 68.780000 92.895000 ;
        RECT 68.610000 68.125000 68.810000 68.325000 ;
        RECT 68.610000 68.535000 68.810000 68.735000 ;
        RECT 68.610000 68.945000 68.810000 69.145000 ;
        RECT 68.610000 69.355000 68.810000 69.555000 ;
        RECT 68.610000 69.765000 68.810000 69.965000 ;
        RECT 68.610000 70.175000 68.810000 70.375000 ;
        RECT 68.610000 70.585000 68.810000 70.785000 ;
        RECT 68.610000 70.995000 68.810000 71.195000 ;
        RECT 68.610000 71.405000 68.810000 71.605000 ;
        RECT 68.610000 71.815000 68.810000 72.015000 ;
        RECT 68.610000 72.225000 68.810000 72.425000 ;
        RECT 68.610000 72.635000 68.810000 72.835000 ;
        RECT 68.610000 73.045000 68.810000 73.245000 ;
        RECT 68.610000 73.450000 68.810000 73.650000 ;
        RECT 68.610000 73.855000 68.810000 74.055000 ;
        RECT 68.610000 74.260000 68.810000 74.460000 ;
        RECT 68.610000 74.665000 68.810000 74.865000 ;
        RECT 68.610000 75.070000 68.810000 75.270000 ;
        RECT 68.610000 75.475000 68.810000 75.675000 ;
        RECT 68.610000 75.880000 68.810000 76.080000 ;
        RECT 68.610000 76.285000 68.810000 76.485000 ;
        RECT 68.610000 76.690000 68.810000 76.890000 ;
        RECT 68.610000 77.095000 68.810000 77.295000 ;
        RECT 68.610000 77.500000 68.810000 77.700000 ;
        RECT 68.610000 77.905000 68.810000 78.105000 ;
        RECT 68.610000 78.310000 68.810000 78.510000 ;
        RECT 68.610000 78.715000 68.810000 78.915000 ;
        RECT 68.610000 79.120000 68.810000 79.320000 ;
        RECT 68.610000 79.525000 68.810000 79.725000 ;
        RECT 68.610000 79.930000 68.810000 80.130000 ;
        RECT 68.610000 80.335000 68.810000 80.535000 ;
        RECT 68.610000 80.740000 68.810000 80.940000 ;
        RECT 68.610000 81.145000 68.810000 81.345000 ;
        RECT 68.610000 81.550000 68.810000 81.750000 ;
        RECT 68.610000 81.955000 68.810000 82.155000 ;
        RECT 68.610000 82.360000 68.810000 82.560000 ;
        RECT 68.665000 17.860000 68.865000 18.060000 ;
        RECT 68.665000 18.290000 68.865000 18.490000 ;
        RECT 68.665000 18.720000 68.865000 18.920000 ;
        RECT 68.665000 19.150000 68.865000 19.350000 ;
        RECT 68.665000 19.580000 68.865000 19.780000 ;
        RECT 68.665000 20.010000 68.865000 20.210000 ;
        RECT 68.665000 20.440000 68.865000 20.640000 ;
        RECT 68.665000 20.870000 68.865000 21.070000 ;
        RECT 68.665000 21.300000 68.865000 21.500000 ;
        RECT 68.665000 21.730000 68.865000 21.930000 ;
        RECT 68.665000 22.160000 68.865000 22.360000 ;
        RECT 68.990000 82.855000 69.190000 83.055000 ;
        RECT 68.990000 83.265000 69.190000 83.465000 ;
        RECT 68.990000 83.675000 69.190000 83.875000 ;
        RECT 68.990000 84.085000 69.190000 84.285000 ;
        RECT 68.990000 84.495000 69.190000 84.695000 ;
        RECT 68.990000 84.905000 69.190000 85.105000 ;
        RECT 68.990000 85.315000 69.190000 85.515000 ;
        RECT 68.990000 85.725000 69.190000 85.925000 ;
        RECT 68.990000 86.135000 69.190000 86.335000 ;
        RECT 68.990000 86.545000 69.190000 86.745000 ;
        RECT 68.990000 86.955000 69.190000 87.155000 ;
        RECT 68.990000 87.365000 69.190000 87.565000 ;
        RECT 68.990000 87.775000 69.190000 87.975000 ;
        RECT 68.990000 88.185000 69.190000 88.385000 ;
        RECT 68.990000 88.595000 69.190000 88.795000 ;
        RECT 68.990000 89.005000 69.190000 89.205000 ;
        RECT 68.990000 89.415000 69.190000 89.615000 ;
        RECT 68.990000 89.825000 69.190000 90.025000 ;
        RECT 68.990000 90.235000 69.190000 90.435000 ;
        RECT 68.990000 90.645000 69.190000 90.845000 ;
        RECT 68.990000 91.055000 69.190000 91.255000 ;
        RECT 68.990000 91.465000 69.190000 91.665000 ;
        RECT 68.990000 91.875000 69.190000 92.075000 ;
        RECT 68.990000 92.285000 69.190000 92.485000 ;
        RECT 68.990000 92.695000 69.190000 92.895000 ;
        RECT 69.010000 68.125000 69.210000 68.325000 ;
        RECT 69.010000 68.535000 69.210000 68.735000 ;
        RECT 69.010000 68.945000 69.210000 69.145000 ;
        RECT 69.010000 69.355000 69.210000 69.555000 ;
        RECT 69.010000 69.765000 69.210000 69.965000 ;
        RECT 69.010000 70.175000 69.210000 70.375000 ;
        RECT 69.010000 70.585000 69.210000 70.785000 ;
        RECT 69.010000 70.995000 69.210000 71.195000 ;
        RECT 69.010000 71.405000 69.210000 71.605000 ;
        RECT 69.010000 71.815000 69.210000 72.015000 ;
        RECT 69.010000 72.225000 69.210000 72.425000 ;
        RECT 69.010000 72.635000 69.210000 72.835000 ;
        RECT 69.010000 73.045000 69.210000 73.245000 ;
        RECT 69.010000 73.450000 69.210000 73.650000 ;
        RECT 69.010000 73.855000 69.210000 74.055000 ;
        RECT 69.010000 74.260000 69.210000 74.460000 ;
        RECT 69.010000 74.665000 69.210000 74.865000 ;
        RECT 69.010000 75.070000 69.210000 75.270000 ;
        RECT 69.010000 75.475000 69.210000 75.675000 ;
        RECT 69.010000 75.880000 69.210000 76.080000 ;
        RECT 69.010000 76.285000 69.210000 76.485000 ;
        RECT 69.010000 76.690000 69.210000 76.890000 ;
        RECT 69.010000 77.095000 69.210000 77.295000 ;
        RECT 69.010000 77.500000 69.210000 77.700000 ;
        RECT 69.010000 77.905000 69.210000 78.105000 ;
        RECT 69.010000 78.310000 69.210000 78.510000 ;
        RECT 69.010000 78.715000 69.210000 78.915000 ;
        RECT 69.010000 79.120000 69.210000 79.320000 ;
        RECT 69.010000 79.525000 69.210000 79.725000 ;
        RECT 69.010000 79.930000 69.210000 80.130000 ;
        RECT 69.010000 80.335000 69.210000 80.535000 ;
        RECT 69.010000 80.740000 69.210000 80.940000 ;
        RECT 69.010000 81.145000 69.210000 81.345000 ;
        RECT 69.010000 81.550000 69.210000 81.750000 ;
        RECT 69.010000 81.955000 69.210000 82.155000 ;
        RECT 69.010000 82.360000 69.210000 82.560000 ;
        RECT 69.070000 17.860000 69.270000 18.060000 ;
        RECT 69.070000 18.290000 69.270000 18.490000 ;
        RECT 69.070000 18.720000 69.270000 18.920000 ;
        RECT 69.070000 19.150000 69.270000 19.350000 ;
        RECT 69.070000 19.580000 69.270000 19.780000 ;
        RECT 69.070000 20.010000 69.270000 20.210000 ;
        RECT 69.070000 20.440000 69.270000 20.640000 ;
        RECT 69.070000 20.870000 69.270000 21.070000 ;
        RECT 69.070000 21.300000 69.270000 21.500000 ;
        RECT 69.070000 21.730000 69.270000 21.930000 ;
        RECT 69.070000 22.160000 69.270000 22.360000 ;
        RECT 69.400000 82.855000 69.600000 83.055000 ;
        RECT 69.400000 83.265000 69.600000 83.465000 ;
        RECT 69.400000 83.675000 69.600000 83.875000 ;
        RECT 69.400000 84.085000 69.600000 84.285000 ;
        RECT 69.400000 84.495000 69.600000 84.695000 ;
        RECT 69.400000 84.905000 69.600000 85.105000 ;
        RECT 69.400000 85.315000 69.600000 85.515000 ;
        RECT 69.400000 85.725000 69.600000 85.925000 ;
        RECT 69.400000 86.135000 69.600000 86.335000 ;
        RECT 69.400000 86.545000 69.600000 86.745000 ;
        RECT 69.400000 86.955000 69.600000 87.155000 ;
        RECT 69.400000 87.365000 69.600000 87.565000 ;
        RECT 69.400000 87.775000 69.600000 87.975000 ;
        RECT 69.400000 88.185000 69.600000 88.385000 ;
        RECT 69.400000 88.595000 69.600000 88.795000 ;
        RECT 69.400000 89.005000 69.600000 89.205000 ;
        RECT 69.400000 89.415000 69.600000 89.615000 ;
        RECT 69.400000 89.825000 69.600000 90.025000 ;
        RECT 69.400000 90.235000 69.600000 90.435000 ;
        RECT 69.400000 90.645000 69.600000 90.845000 ;
        RECT 69.400000 91.055000 69.600000 91.255000 ;
        RECT 69.400000 91.465000 69.600000 91.665000 ;
        RECT 69.400000 91.875000 69.600000 92.075000 ;
        RECT 69.400000 92.285000 69.600000 92.485000 ;
        RECT 69.400000 92.695000 69.600000 92.895000 ;
        RECT 69.410000 68.125000 69.610000 68.325000 ;
        RECT 69.410000 68.535000 69.610000 68.735000 ;
        RECT 69.410000 68.945000 69.610000 69.145000 ;
        RECT 69.410000 69.355000 69.610000 69.555000 ;
        RECT 69.410000 69.765000 69.610000 69.965000 ;
        RECT 69.410000 70.175000 69.610000 70.375000 ;
        RECT 69.410000 70.585000 69.610000 70.785000 ;
        RECT 69.410000 70.995000 69.610000 71.195000 ;
        RECT 69.410000 71.405000 69.610000 71.605000 ;
        RECT 69.410000 71.815000 69.610000 72.015000 ;
        RECT 69.410000 72.225000 69.610000 72.425000 ;
        RECT 69.410000 72.635000 69.610000 72.835000 ;
        RECT 69.410000 73.045000 69.610000 73.245000 ;
        RECT 69.410000 73.450000 69.610000 73.650000 ;
        RECT 69.410000 73.855000 69.610000 74.055000 ;
        RECT 69.410000 74.260000 69.610000 74.460000 ;
        RECT 69.410000 74.665000 69.610000 74.865000 ;
        RECT 69.410000 75.070000 69.610000 75.270000 ;
        RECT 69.410000 75.475000 69.610000 75.675000 ;
        RECT 69.410000 75.880000 69.610000 76.080000 ;
        RECT 69.410000 76.285000 69.610000 76.485000 ;
        RECT 69.410000 76.690000 69.610000 76.890000 ;
        RECT 69.410000 77.095000 69.610000 77.295000 ;
        RECT 69.410000 77.500000 69.610000 77.700000 ;
        RECT 69.410000 77.905000 69.610000 78.105000 ;
        RECT 69.410000 78.310000 69.610000 78.510000 ;
        RECT 69.410000 78.715000 69.610000 78.915000 ;
        RECT 69.410000 79.120000 69.610000 79.320000 ;
        RECT 69.410000 79.525000 69.610000 79.725000 ;
        RECT 69.410000 79.930000 69.610000 80.130000 ;
        RECT 69.410000 80.335000 69.610000 80.535000 ;
        RECT 69.410000 80.740000 69.610000 80.940000 ;
        RECT 69.410000 81.145000 69.610000 81.345000 ;
        RECT 69.410000 81.550000 69.610000 81.750000 ;
        RECT 69.410000 81.955000 69.610000 82.155000 ;
        RECT 69.410000 82.360000 69.610000 82.560000 ;
        RECT 69.475000 17.860000 69.675000 18.060000 ;
        RECT 69.475000 18.290000 69.675000 18.490000 ;
        RECT 69.475000 18.720000 69.675000 18.920000 ;
        RECT 69.475000 19.150000 69.675000 19.350000 ;
        RECT 69.475000 19.580000 69.675000 19.780000 ;
        RECT 69.475000 20.010000 69.675000 20.210000 ;
        RECT 69.475000 20.440000 69.675000 20.640000 ;
        RECT 69.475000 20.870000 69.675000 21.070000 ;
        RECT 69.475000 21.300000 69.675000 21.500000 ;
        RECT 69.475000 21.730000 69.675000 21.930000 ;
        RECT 69.475000 22.160000 69.675000 22.360000 ;
        RECT 69.810000 68.125000 70.010000 68.325000 ;
        RECT 69.810000 68.535000 70.010000 68.735000 ;
        RECT 69.810000 68.945000 70.010000 69.145000 ;
        RECT 69.810000 69.355000 70.010000 69.555000 ;
        RECT 69.810000 69.765000 70.010000 69.965000 ;
        RECT 69.810000 70.175000 70.010000 70.375000 ;
        RECT 69.810000 70.585000 70.010000 70.785000 ;
        RECT 69.810000 70.995000 70.010000 71.195000 ;
        RECT 69.810000 71.405000 70.010000 71.605000 ;
        RECT 69.810000 71.815000 70.010000 72.015000 ;
        RECT 69.810000 72.225000 70.010000 72.425000 ;
        RECT 69.810000 72.635000 70.010000 72.835000 ;
        RECT 69.810000 73.045000 70.010000 73.245000 ;
        RECT 69.810000 73.450000 70.010000 73.650000 ;
        RECT 69.810000 73.855000 70.010000 74.055000 ;
        RECT 69.810000 74.260000 70.010000 74.460000 ;
        RECT 69.810000 74.665000 70.010000 74.865000 ;
        RECT 69.810000 75.070000 70.010000 75.270000 ;
        RECT 69.810000 75.475000 70.010000 75.675000 ;
        RECT 69.810000 75.880000 70.010000 76.080000 ;
        RECT 69.810000 76.285000 70.010000 76.485000 ;
        RECT 69.810000 76.690000 70.010000 76.890000 ;
        RECT 69.810000 77.095000 70.010000 77.295000 ;
        RECT 69.810000 77.500000 70.010000 77.700000 ;
        RECT 69.810000 77.905000 70.010000 78.105000 ;
        RECT 69.810000 78.310000 70.010000 78.510000 ;
        RECT 69.810000 78.715000 70.010000 78.915000 ;
        RECT 69.810000 79.120000 70.010000 79.320000 ;
        RECT 69.810000 79.525000 70.010000 79.725000 ;
        RECT 69.810000 79.930000 70.010000 80.130000 ;
        RECT 69.810000 80.335000 70.010000 80.535000 ;
        RECT 69.810000 80.740000 70.010000 80.940000 ;
        RECT 69.810000 81.145000 70.010000 81.345000 ;
        RECT 69.810000 81.550000 70.010000 81.750000 ;
        RECT 69.810000 81.955000 70.010000 82.155000 ;
        RECT 69.810000 82.360000 70.010000 82.560000 ;
        RECT 69.810000 82.855000 70.010000 83.055000 ;
        RECT 69.810000 83.265000 70.010000 83.465000 ;
        RECT 69.810000 83.675000 70.010000 83.875000 ;
        RECT 69.810000 84.085000 70.010000 84.285000 ;
        RECT 69.810000 84.495000 70.010000 84.695000 ;
        RECT 69.810000 84.905000 70.010000 85.105000 ;
        RECT 69.810000 85.315000 70.010000 85.515000 ;
        RECT 69.810000 85.725000 70.010000 85.925000 ;
        RECT 69.810000 86.135000 70.010000 86.335000 ;
        RECT 69.810000 86.545000 70.010000 86.745000 ;
        RECT 69.810000 86.955000 70.010000 87.155000 ;
        RECT 69.810000 87.365000 70.010000 87.565000 ;
        RECT 69.810000 87.775000 70.010000 87.975000 ;
        RECT 69.810000 88.185000 70.010000 88.385000 ;
        RECT 69.810000 88.595000 70.010000 88.795000 ;
        RECT 69.810000 89.005000 70.010000 89.205000 ;
        RECT 69.810000 89.415000 70.010000 89.615000 ;
        RECT 69.810000 89.825000 70.010000 90.025000 ;
        RECT 69.810000 90.235000 70.010000 90.435000 ;
        RECT 69.810000 90.645000 70.010000 90.845000 ;
        RECT 69.810000 91.055000 70.010000 91.255000 ;
        RECT 69.810000 91.465000 70.010000 91.665000 ;
        RECT 69.810000 91.875000 70.010000 92.075000 ;
        RECT 69.810000 92.285000 70.010000 92.485000 ;
        RECT 69.810000 92.695000 70.010000 92.895000 ;
        RECT 69.880000 17.860000 70.080000 18.060000 ;
        RECT 69.880000 18.290000 70.080000 18.490000 ;
        RECT 69.880000 18.720000 70.080000 18.920000 ;
        RECT 69.880000 19.150000 70.080000 19.350000 ;
        RECT 69.880000 19.580000 70.080000 19.780000 ;
        RECT 69.880000 20.010000 70.080000 20.210000 ;
        RECT 69.880000 20.440000 70.080000 20.640000 ;
        RECT 69.880000 20.870000 70.080000 21.070000 ;
        RECT 69.880000 21.300000 70.080000 21.500000 ;
        RECT 69.880000 21.730000 70.080000 21.930000 ;
        RECT 69.880000 22.160000 70.080000 22.360000 ;
        RECT 70.210000 68.125000 70.410000 68.325000 ;
        RECT 70.210000 68.535000 70.410000 68.735000 ;
        RECT 70.210000 68.945000 70.410000 69.145000 ;
        RECT 70.210000 69.355000 70.410000 69.555000 ;
        RECT 70.210000 69.765000 70.410000 69.965000 ;
        RECT 70.210000 70.175000 70.410000 70.375000 ;
        RECT 70.210000 70.585000 70.410000 70.785000 ;
        RECT 70.210000 70.995000 70.410000 71.195000 ;
        RECT 70.210000 71.405000 70.410000 71.605000 ;
        RECT 70.210000 71.815000 70.410000 72.015000 ;
        RECT 70.210000 72.225000 70.410000 72.425000 ;
        RECT 70.210000 72.635000 70.410000 72.835000 ;
        RECT 70.210000 73.045000 70.410000 73.245000 ;
        RECT 70.210000 73.450000 70.410000 73.650000 ;
        RECT 70.210000 73.855000 70.410000 74.055000 ;
        RECT 70.210000 74.260000 70.410000 74.460000 ;
        RECT 70.210000 74.665000 70.410000 74.865000 ;
        RECT 70.210000 75.070000 70.410000 75.270000 ;
        RECT 70.210000 75.475000 70.410000 75.675000 ;
        RECT 70.210000 75.880000 70.410000 76.080000 ;
        RECT 70.210000 76.285000 70.410000 76.485000 ;
        RECT 70.210000 76.690000 70.410000 76.890000 ;
        RECT 70.210000 77.095000 70.410000 77.295000 ;
        RECT 70.210000 77.500000 70.410000 77.700000 ;
        RECT 70.210000 77.905000 70.410000 78.105000 ;
        RECT 70.210000 78.310000 70.410000 78.510000 ;
        RECT 70.210000 78.715000 70.410000 78.915000 ;
        RECT 70.210000 79.120000 70.410000 79.320000 ;
        RECT 70.210000 79.525000 70.410000 79.725000 ;
        RECT 70.210000 79.930000 70.410000 80.130000 ;
        RECT 70.210000 80.335000 70.410000 80.535000 ;
        RECT 70.210000 80.740000 70.410000 80.940000 ;
        RECT 70.210000 81.145000 70.410000 81.345000 ;
        RECT 70.210000 81.550000 70.410000 81.750000 ;
        RECT 70.210000 81.955000 70.410000 82.155000 ;
        RECT 70.210000 82.360000 70.410000 82.560000 ;
        RECT 70.220000 82.855000 70.420000 83.055000 ;
        RECT 70.220000 83.265000 70.420000 83.465000 ;
        RECT 70.220000 83.675000 70.420000 83.875000 ;
        RECT 70.220000 84.085000 70.420000 84.285000 ;
        RECT 70.220000 84.495000 70.420000 84.695000 ;
        RECT 70.220000 84.905000 70.420000 85.105000 ;
        RECT 70.220000 85.315000 70.420000 85.515000 ;
        RECT 70.220000 85.725000 70.420000 85.925000 ;
        RECT 70.220000 86.135000 70.420000 86.335000 ;
        RECT 70.220000 86.545000 70.420000 86.745000 ;
        RECT 70.220000 86.955000 70.420000 87.155000 ;
        RECT 70.220000 87.365000 70.420000 87.565000 ;
        RECT 70.220000 87.775000 70.420000 87.975000 ;
        RECT 70.220000 88.185000 70.420000 88.385000 ;
        RECT 70.220000 88.595000 70.420000 88.795000 ;
        RECT 70.220000 89.005000 70.420000 89.205000 ;
        RECT 70.220000 89.415000 70.420000 89.615000 ;
        RECT 70.220000 89.825000 70.420000 90.025000 ;
        RECT 70.220000 90.235000 70.420000 90.435000 ;
        RECT 70.220000 90.645000 70.420000 90.845000 ;
        RECT 70.220000 91.055000 70.420000 91.255000 ;
        RECT 70.220000 91.465000 70.420000 91.665000 ;
        RECT 70.220000 91.875000 70.420000 92.075000 ;
        RECT 70.220000 92.285000 70.420000 92.485000 ;
        RECT 70.220000 92.695000 70.420000 92.895000 ;
        RECT 70.285000 17.860000 70.485000 18.060000 ;
        RECT 70.285000 18.290000 70.485000 18.490000 ;
        RECT 70.285000 18.720000 70.485000 18.920000 ;
        RECT 70.285000 19.150000 70.485000 19.350000 ;
        RECT 70.285000 19.580000 70.485000 19.780000 ;
        RECT 70.285000 20.010000 70.485000 20.210000 ;
        RECT 70.285000 20.440000 70.485000 20.640000 ;
        RECT 70.285000 20.870000 70.485000 21.070000 ;
        RECT 70.285000 21.300000 70.485000 21.500000 ;
        RECT 70.285000 21.730000 70.485000 21.930000 ;
        RECT 70.285000 22.160000 70.485000 22.360000 ;
        RECT 70.610000 68.125000 70.810000 68.325000 ;
        RECT 70.610000 68.535000 70.810000 68.735000 ;
        RECT 70.610000 68.945000 70.810000 69.145000 ;
        RECT 70.610000 69.355000 70.810000 69.555000 ;
        RECT 70.610000 69.765000 70.810000 69.965000 ;
        RECT 70.610000 70.175000 70.810000 70.375000 ;
        RECT 70.610000 70.585000 70.810000 70.785000 ;
        RECT 70.610000 70.995000 70.810000 71.195000 ;
        RECT 70.610000 71.405000 70.810000 71.605000 ;
        RECT 70.610000 71.815000 70.810000 72.015000 ;
        RECT 70.610000 72.225000 70.810000 72.425000 ;
        RECT 70.610000 72.635000 70.810000 72.835000 ;
        RECT 70.610000 73.045000 70.810000 73.245000 ;
        RECT 70.610000 73.450000 70.810000 73.650000 ;
        RECT 70.610000 73.855000 70.810000 74.055000 ;
        RECT 70.610000 74.260000 70.810000 74.460000 ;
        RECT 70.610000 74.665000 70.810000 74.865000 ;
        RECT 70.610000 75.070000 70.810000 75.270000 ;
        RECT 70.610000 75.475000 70.810000 75.675000 ;
        RECT 70.610000 75.880000 70.810000 76.080000 ;
        RECT 70.610000 76.285000 70.810000 76.485000 ;
        RECT 70.610000 76.690000 70.810000 76.890000 ;
        RECT 70.610000 77.095000 70.810000 77.295000 ;
        RECT 70.610000 77.500000 70.810000 77.700000 ;
        RECT 70.610000 77.905000 70.810000 78.105000 ;
        RECT 70.610000 78.310000 70.810000 78.510000 ;
        RECT 70.610000 78.715000 70.810000 78.915000 ;
        RECT 70.610000 79.120000 70.810000 79.320000 ;
        RECT 70.610000 79.525000 70.810000 79.725000 ;
        RECT 70.610000 79.930000 70.810000 80.130000 ;
        RECT 70.610000 80.335000 70.810000 80.535000 ;
        RECT 70.610000 80.740000 70.810000 80.940000 ;
        RECT 70.610000 81.145000 70.810000 81.345000 ;
        RECT 70.610000 81.550000 70.810000 81.750000 ;
        RECT 70.610000 81.955000 70.810000 82.155000 ;
        RECT 70.610000 82.360000 70.810000 82.560000 ;
        RECT 70.630000 82.855000 70.830000 83.055000 ;
        RECT 70.630000 83.265000 70.830000 83.465000 ;
        RECT 70.630000 83.675000 70.830000 83.875000 ;
        RECT 70.630000 84.085000 70.830000 84.285000 ;
        RECT 70.630000 84.495000 70.830000 84.695000 ;
        RECT 70.630000 84.905000 70.830000 85.105000 ;
        RECT 70.630000 85.315000 70.830000 85.515000 ;
        RECT 70.630000 85.725000 70.830000 85.925000 ;
        RECT 70.630000 86.135000 70.830000 86.335000 ;
        RECT 70.630000 86.545000 70.830000 86.745000 ;
        RECT 70.630000 86.955000 70.830000 87.155000 ;
        RECT 70.630000 87.365000 70.830000 87.565000 ;
        RECT 70.630000 87.775000 70.830000 87.975000 ;
        RECT 70.630000 88.185000 70.830000 88.385000 ;
        RECT 70.630000 88.595000 70.830000 88.795000 ;
        RECT 70.630000 89.005000 70.830000 89.205000 ;
        RECT 70.630000 89.415000 70.830000 89.615000 ;
        RECT 70.630000 89.825000 70.830000 90.025000 ;
        RECT 70.630000 90.235000 70.830000 90.435000 ;
        RECT 70.630000 90.645000 70.830000 90.845000 ;
        RECT 70.630000 91.055000 70.830000 91.255000 ;
        RECT 70.630000 91.465000 70.830000 91.665000 ;
        RECT 70.630000 91.875000 70.830000 92.075000 ;
        RECT 70.630000 92.285000 70.830000 92.485000 ;
        RECT 70.630000 92.695000 70.830000 92.895000 ;
        RECT 70.690000 17.860000 70.890000 18.060000 ;
        RECT 70.690000 18.290000 70.890000 18.490000 ;
        RECT 70.690000 18.720000 70.890000 18.920000 ;
        RECT 70.690000 19.150000 70.890000 19.350000 ;
        RECT 70.690000 19.580000 70.890000 19.780000 ;
        RECT 70.690000 20.010000 70.890000 20.210000 ;
        RECT 70.690000 20.440000 70.890000 20.640000 ;
        RECT 70.690000 20.870000 70.890000 21.070000 ;
        RECT 70.690000 21.300000 70.890000 21.500000 ;
        RECT 70.690000 21.730000 70.890000 21.930000 ;
        RECT 70.690000 22.160000 70.890000 22.360000 ;
        RECT 71.010000 68.125000 71.210000 68.325000 ;
        RECT 71.010000 68.535000 71.210000 68.735000 ;
        RECT 71.010000 68.945000 71.210000 69.145000 ;
        RECT 71.010000 69.355000 71.210000 69.555000 ;
        RECT 71.010000 69.765000 71.210000 69.965000 ;
        RECT 71.010000 70.175000 71.210000 70.375000 ;
        RECT 71.010000 70.585000 71.210000 70.785000 ;
        RECT 71.010000 70.995000 71.210000 71.195000 ;
        RECT 71.010000 71.405000 71.210000 71.605000 ;
        RECT 71.010000 71.815000 71.210000 72.015000 ;
        RECT 71.010000 72.225000 71.210000 72.425000 ;
        RECT 71.010000 72.635000 71.210000 72.835000 ;
        RECT 71.010000 73.045000 71.210000 73.245000 ;
        RECT 71.010000 73.450000 71.210000 73.650000 ;
        RECT 71.010000 73.855000 71.210000 74.055000 ;
        RECT 71.010000 74.260000 71.210000 74.460000 ;
        RECT 71.010000 74.665000 71.210000 74.865000 ;
        RECT 71.010000 75.070000 71.210000 75.270000 ;
        RECT 71.010000 75.475000 71.210000 75.675000 ;
        RECT 71.010000 75.880000 71.210000 76.080000 ;
        RECT 71.010000 76.285000 71.210000 76.485000 ;
        RECT 71.010000 76.690000 71.210000 76.890000 ;
        RECT 71.010000 77.095000 71.210000 77.295000 ;
        RECT 71.010000 77.500000 71.210000 77.700000 ;
        RECT 71.010000 77.905000 71.210000 78.105000 ;
        RECT 71.010000 78.310000 71.210000 78.510000 ;
        RECT 71.010000 78.715000 71.210000 78.915000 ;
        RECT 71.010000 79.120000 71.210000 79.320000 ;
        RECT 71.010000 79.525000 71.210000 79.725000 ;
        RECT 71.010000 79.930000 71.210000 80.130000 ;
        RECT 71.010000 80.335000 71.210000 80.535000 ;
        RECT 71.010000 80.740000 71.210000 80.940000 ;
        RECT 71.010000 81.145000 71.210000 81.345000 ;
        RECT 71.010000 81.550000 71.210000 81.750000 ;
        RECT 71.010000 81.955000 71.210000 82.155000 ;
        RECT 71.010000 82.360000 71.210000 82.560000 ;
        RECT 71.040000 82.855000 71.240000 83.055000 ;
        RECT 71.040000 83.265000 71.240000 83.465000 ;
        RECT 71.040000 83.675000 71.240000 83.875000 ;
        RECT 71.040000 84.085000 71.240000 84.285000 ;
        RECT 71.040000 84.495000 71.240000 84.695000 ;
        RECT 71.040000 84.905000 71.240000 85.105000 ;
        RECT 71.040000 85.315000 71.240000 85.515000 ;
        RECT 71.040000 85.725000 71.240000 85.925000 ;
        RECT 71.040000 86.135000 71.240000 86.335000 ;
        RECT 71.040000 86.545000 71.240000 86.745000 ;
        RECT 71.040000 86.955000 71.240000 87.155000 ;
        RECT 71.040000 87.365000 71.240000 87.565000 ;
        RECT 71.040000 87.775000 71.240000 87.975000 ;
        RECT 71.040000 88.185000 71.240000 88.385000 ;
        RECT 71.040000 88.595000 71.240000 88.795000 ;
        RECT 71.040000 89.005000 71.240000 89.205000 ;
        RECT 71.040000 89.415000 71.240000 89.615000 ;
        RECT 71.040000 89.825000 71.240000 90.025000 ;
        RECT 71.040000 90.235000 71.240000 90.435000 ;
        RECT 71.040000 90.645000 71.240000 90.845000 ;
        RECT 71.040000 91.055000 71.240000 91.255000 ;
        RECT 71.040000 91.465000 71.240000 91.665000 ;
        RECT 71.040000 91.875000 71.240000 92.075000 ;
        RECT 71.040000 92.285000 71.240000 92.485000 ;
        RECT 71.040000 92.695000 71.240000 92.895000 ;
        RECT 71.095000 17.860000 71.295000 18.060000 ;
        RECT 71.095000 18.290000 71.295000 18.490000 ;
        RECT 71.095000 18.720000 71.295000 18.920000 ;
        RECT 71.095000 19.150000 71.295000 19.350000 ;
        RECT 71.095000 19.580000 71.295000 19.780000 ;
        RECT 71.095000 20.010000 71.295000 20.210000 ;
        RECT 71.095000 20.440000 71.295000 20.640000 ;
        RECT 71.095000 20.870000 71.295000 21.070000 ;
        RECT 71.095000 21.300000 71.295000 21.500000 ;
        RECT 71.095000 21.730000 71.295000 21.930000 ;
        RECT 71.095000 22.160000 71.295000 22.360000 ;
        RECT 71.410000 68.125000 71.610000 68.325000 ;
        RECT 71.410000 68.535000 71.610000 68.735000 ;
        RECT 71.410000 68.945000 71.610000 69.145000 ;
        RECT 71.410000 69.355000 71.610000 69.555000 ;
        RECT 71.410000 69.765000 71.610000 69.965000 ;
        RECT 71.410000 70.175000 71.610000 70.375000 ;
        RECT 71.410000 70.585000 71.610000 70.785000 ;
        RECT 71.410000 70.995000 71.610000 71.195000 ;
        RECT 71.410000 71.405000 71.610000 71.605000 ;
        RECT 71.410000 71.815000 71.610000 72.015000 ;
        RECT 71.410000 72.225000 71.610000 72.425000 ;
        RECT 71.410000 72.635000 71.610000 72.835000 ;
        RECT 71.410000 73.045000 71.610000 73.245000 ;
        RECT 71.410000 73.450000 71.610000 73.650000 ;
        RECT 71.410000 73.855000 71.610000 74.055000 ;
        RECT 71.410000 74.260000 71.610000 74.460000 ;
        RECT 71.410000 74.665000 71.610000 74.865000 ;
        RECT 71.410000 75.070000 71.610000 75.270000 ;
        RECT 71.410000 75.475000 71.610000 75.675000 ;
        RECT 71.410000 75.880000 71.610000 76.080000 ;
        RECT 71.410000 76.285000 71.610000 76.485000 ;
        RECT 71.410000 76.690000 71.610000 76.890000 ;
        RECT 71.410000 77.095000 71.610000 77.295000 ;
        RECT 71.410000 77.500000 71.610000 77.700000 ;
        RECT 71.410000 77.905000 71.610000 78.105000 ;
        RECT 71.410000 78.310000 71.610000 78.510000 ;
        RECT 71.410000 78.715000 71.610000 78.915000 ;
        RECT 71.410000 79.120000 71.610000 79.320000 ;
        RECT 71.410000 79.525000 71.610000 79.725000 ;
        RECT 71.410000 79.930000 71.610000 80.130000 ;
        RECT 71.410000 80.335000 71.610000 80.535000 ;
        RECT 71.410000 80.740000 71.610000 80.940000 ;
        RECT 71.410000 81.145000 71.610000 81.345000 ;
        RECT 71.410000 81.550000 71.610000 81.750000 ;
        RECT 71.410000 81.955000 71.610000 82.155000 ;
        RECT 71.410000 82.360000 71.610000 82.560000 ;
        RECT 71.450000 82.855000 71.650000 83.055000 ;
        RECT 71.450000 83.265000 71.650000 83.465000 ;
        RECT 71.450000 83.675000 71.650000 83.875000 ;
        RECT 71.450000 84.085000 71.650000 84.285000 ;
        RECT 71.450000 84.495000 71.650000 84.695000 ;
        RECT 71.450000 84.905000 71.650000 85.105000 ;
        RECT 71.450000 85.315000 71.650000 85.515000 ;
        RECT 71.450000 85.725000 71.650000 85.925000 ;
        RECT 71.450000 86.135000 71.650000 86.335000 ;
        RECT 71.450000 86.545000 71.650000 86.745000 ;
        RECT 71.450000 86.955000 71.650000 87.155000 ;
        RECT 71.450000 87.365000 71.650000 87.565000 ;
        RECT 71.450000 87.775000 71.650000 87.975000 ;
        RECT 71.450000 88.185000 71.650000 88.385000 ;
        RECT 71.450000 88.595000 71.650000 88.795000 ;
        RECT 71.450000 89.005000 71.650000 89.205000 ;
        RECT 71.450000 89.415000 71.650000 89.615000 ;
        RECT 71.450000 89.825000 71.650000 90.025000 ;
        RECT 71.450000 90.235000 71.650000 90.435000 ;
        RECT 71.450000 90.645000 71.650000 90.845000 ;
        RECT 71.450000 91.055000 71.650000 91.255000 ;
        RECT 71.450000 91.465000 71.650000 91.665000 ;
        RECT 71.450000 91.875000 71.650000 92.075000 ;
        RECT 71.450000 92.285000 71.650000 92.485000 ;
        RECT 71.450000 92.695000 71.650000 92.895000 ;
        RECT 71.500000 17.860000 71.700000 18.060000 ;
        RECT 71.500000 18.290000 71.700000 18.490000 ;
        RECT 71.500000 18.720000 71.700000 18.920000 ;
        RECT 71.500000 19.150000 71.700000 19.350000 ;
        RECT 71.500000 19.580000 71.700000 19.780000 ;
        RECT 71.500000 20.010000 71.700000 20.210000 ;
        RECT 71.500000 20.440000 71.700000 20.640000 ;
        RECT 71.500000 20.870000 71.700000 21.070000 ;
        RECT 71.500000 21.300000 71.700000 21.500000 ;
        RECT 71.500000 21.730000 71.700000 21.930000 ;
        RECT 71.500000 22.160000 71.700000 22.360000 ;
        RECT 71.810000 68.125000 72.010000 68.325000 ;
        RECT 71.810000 68.535000 72.010000 68.735000 ;
        RECT 71.810000 68.945000 72.010000 69.145000 ;
        RECT 71.810000 69.355000 72.010000 69.555000 ;
        RECT 71.810000 69.765000 72.010000 69.965000 ;
        RECT 71.810000 70.175000 72.010000 70.375000 ;
        RECT 71.810000 70.585000 72.010000 70.785000 ;
        RECT 71.810000 70.995000 72.010000 71.195000 ;
        RECT 71.810000 71.405000 72.010000 71.605000 ;
        RECT 71.810000 71.815000 72.010000 72.015000 ;
        RECT 71.810000 72.225000 72.010000 72.425000 ;
        RECT 71.810000 72.635000 72.010000 72.835000 ;
        RECT 71.810000 73.045000 72.010000 73.245000 ;
        RECT 71.810000 73.450000 72.010000 73.650000 ;
        RECT 71.810000 73.855000 72.010000 74.055000 ;
        RECT 71.810000 74.260000 72.010000 74.460000 ;
        RECT 71.810000 74.665000 72.010000 74.865000 ;
        RECT 71.810000 75.070000 72.010000 75.270000 ;
        RECT 71.810000 75.475000 72.010000 75.675000 ;
        RECT 71.810000 75.880000 72.010000 76.080000 ;
        RECT 71.810000 76.285000 72.010000 76.485000 ;
        RECT 71.810000 76.690000 72.010000 76.890000 ;
        RECT 71.810000 77.095000 72.010000 77.295000 ;
        RECT 71.810000 77.500000 72.010000 77.700000 ;
        RECT 71.810000 77.905000 72.010000 78.105000 ;
        RECT 71.810000 78.310000 72.010000 78.510000 ;
        RECT 71.810000 78.715000 72.010000 78.915000 ;
        RECT 71.810000 79.120000 72.010000 79.320000 ;
        RECT 71.810000 79.525000 72.010000 79.725000 ;
        RECT 71.810000 79.930000 72.010000 80.130000 ;
        RECT 71.810000 80.335000 72.010000 80.535000 ;
        RECT 71.810000 80.740000 72.010000 80.940000 ;
        RECT 71.810000 81.145000 72.010000 81.345000 ;
        RECT 71.810000 81.550000 72.010000 81.750000 ;
        RECT 71.810000 81.955000 72.010000 82.155000 ;
        RECT 71.810000 82.360000 72.010000 82.560000 ;
        RECT 71.860000 82.855000 72.060000 83.055000 ;
        RECT 71.860000 83.265000 72.060000 83.465000 ;
        RECT 71.860000 83.675000 72.060000 83.875000 ;
        RECT 71.860000 84.085000 72.060000 84.285000 ;
        RECT 71.860000 84.495000 72.060000 84.695000 ;
        RECT 71.860000 84.905000 72.060000 85.105000 ;
        RECT 71.860000 85.315000 72.060000 85.515000 ;
        RECT 71.860000 85.725000 72.060000 85.925000 ;
        RECT 71.860000 86.135000 72.060000 86.335000 ;
        RECT 71.860000 86.545000 72.060000 86.745000 ;
        RECT 71.860000 86.955000 72.060000 87.155000 ;
        RECT 71.860000 87.365000 72.060000 87.565000 ;
        RECT 71.860000 87.775000 72.060000 87.975000 ;
        RECT 71.860000 88.185000 72.060000 88.385000 ;
        RECT 71.860000 88.595000 72.060000 88.795000 ;
        RECT 71.860000 89.005000 72.060000 89.205000 ;
        RECT 71.860000 89.415000 72.060000 89.615000 ;
        RECT 71.860000 89.825000 72.060000 90.025000 ;
        RECT 71.860000 90.235000 72.060000 90.435000 ;
        RECT 71.860000 90.645000 72.060000 90.845000 ;
        RECT 71.860000 91.055000 72.060000 91.255000 ;
        RECT 71.860000 91.465000 72.060000 91.665000 ;
        RECT 71.860000 91.875000 72.060000 92.075000 ;
        RECT 71.860000 92.285000 72.060000 92.485000 ;
        RECT 71.860000 92.695000 72.060000 92.895000 ;
        RECT 71.905000 17.860000 72.105000 18.060000 ;
        RECT 71.905000 18.290000 72.105000 18.490000 ;
        RECT 71.905000 18.720000 72.105000 18.920000 ;
        RECT 71.905000 19.150000 72.105000 19.350000 ;
        RECT 71.905000 19.580000 72.105000 19.780000 ;
        RECT 71.905000 20.010000 72.105000 20.210000 ;
        RECT 71.905000 20.440000 72.105000 20.640000 ;
        RECT 71.905000 20.870000 72.105000 21.070000 ;
        RECT 71.905000 21.300000 72.105000 21.500000 ;
        RECT 71.905000 21.730000 72.105000 21.930000 ;
        RECT 71.905000 22.160000 72.105000 22.360000 ;
        RECT 72.210000 68.125000 72.410000 68.325000 ;
        RECT 72.210000 68.535000 72.410000 68.735000 ;
        RECT 72.210000 68.945000 72.410000 69.145000 ;
        RECT 72.210000 69.355000 72.410000 69.555000 ;
        RECT 72.210000 69.765000 72.410000 69.965000 ;
        RECT 72.210000 70.175000 72.410000 70.375000 ;
        RECT 72.210000 70.585000 72.410000 70.785000 ;
        RECT 72.210000 70.995000 72.410000 71.195000 ;
        RECT 72.210000 71.405000 72.410000 71.605000 ;
        RECT 72.210000 71.815000 72.410000 72.015000 ;
        RECT 72.210000 72.225000 72.410000 72.425000 ;
        RECT 72.210000 72.635000 72.410000 72.835000 ;
        RECT 72.210000 73.045000 72.410000 73.245000 ;
        RECT 72.210000 73.450000 72.410000 73.650000 ;
        RECT 72.210000 73.855000 72.410000 74.055000 ;
        RECT 72.210000 74.260000 72.410000 74.460000 ;
        RECT 72.210000 74.665000 72.410000 74.865000 ;
        RECT 72.210000 75.070000 72.410000 75.270000 ;
        RECT 72.210000 75.475000 72.410000 75.675000 ;
        RECT 72.210000 75.880000 72.410000 76.080000 ;
        RECT 72.210000 76.285000 72.410000 76.485000 ;
        RECT 72.210000 76.690000 72.410000 76.890000 ;
        RECT 72.210000 77.095000 72.410000 77.295000 ;
        RECT 72.210000 77.500000 72.410000 77.700000 ;
        RECT 72.210000 77.905000 72.410000 78.105000 ;
        RECT 72.210000 78.310000 72.410000 78.510000 ;
        RECT 72.210000 78.715000 72.410000 78.915000 ;
        RECT 72.210000 79.120000 72.410000 79.320000 ;
        RECT 72.210000 79.525000 72.410000 79.725000 ;
        RECT 72.210000 79.930000 72.410000 80.130000 ;
        RECT 72.210000 80.335000 72.410000 80.535000 ;
        RECT 72.210000 80.740000 72.410000 80.940000 ;
        RECT 72.210000 81.145000 72.410000 81.345000 ;
        RECT 72.210000 81.550000 72.410000 81.750000 ;
        RECT 72.210000 81.955000 72.410000 82.155000 ;
        RECT 72.210000 82.360000 72.410000 82.560000 ;
        RECT 72.270000 82.855000 72.470000 83.055000 ;
        RECT 72.270000 83.265000 72.470000 83.465000 ;
        RECT 72.270000 83.675000 72.470000 83.875000 ;
        RECT 72.270000 84.085000 72.470000 84.285000 ;
        RECT 72.270000 84.495000 72.470000 84.695000 ;
        RECT 72.270000 84.905000 72.470000 85.105000 ;
        RECT 72.270000 85.315000 72.470000 85.515000 ;
        RECT 72.270000 85.725000 72.470000 85.925000 ;
        RECT 72.270000 86.135000 72.470000 86.335000 ;
        RECT 72.270000 86.545000 72.470000 86.745000 ;
        RECT 72.270000 86.955000 72.470000 87.155000 ;
        RECT 72.270000 87.365000 72.470000 87.565000 ;
        RECT 72.270000 87.775000 72.470000 87.975000 ;
        RECT 72.270000 88.185000 72.470000 88.385000 ;
        RECT 72.270000 88.595000 72.470000 88.795000 ;
        RECT 72.270000 89.005000 72.470000 89.205000 ;
        RECT 72.270000 89.415000 72.470000 89.615000 ;
        RECT 72.270000 89.825000 72.470000 90.025000 ;
        RECT 72.270000 90.235000 72.470000 90.435000 ;
        RECT 72.270000 90.645000 72.470000 90.845000 ;
        RECT 72.270000 91.055000 72.470000 91.255000 ;
        RECT 72.270000 91.465000 72.470000 91.665000 ;
        RECT 72.270000 91.875000 72.470000 92.075000 ;
        RECT 72.270000 92.285000 72.470000 92.485000 ;
        RECT 72.270000 92.695000 72.470000 92.895000 ;
        RECT 72.315000 17.860000 72.515000 18.060000 ;
        RECT 72.315000 18.290000 72.515000 18.490000 ;
        RECT 72.315000 18.720000 72.515000 18.920000 ;
        RECT 72.315000 19.150000 72.515000 19.350000 ;
        RECT 72.315000 19.580000 72.515000 19.780000 ;
        RECT 72.315000 20.010000 72.515000 20.210000 ;
        RECT 72.315000 20.440000 72.515000 20.640000 ;
        RECT 72.315000 20.870000 72.515000 21.070000 ;
        RECT 72.315000 21.300000 72.515000 21.500000 ;
        RECT 72.315000 21.730000 72.515000 21.930000 ;
        RECT 72.315000 22.160000 72.515000 22.360000 ;
        RECT 72.610000 68.125000 72.810000 68.325000 ;
        RECT 72.610000 68.535000 72.810000 68.735000 ;
        RECT 72.610000 68.945000 72.810000 69.145000 ;
        RECT 72.610000 69.355000 72.810000 69.555000 ;
        RECT 72.610000 69.765000 72.810000 69.965000 ;
        RECT 72.610000 70.175000 72.810000 70.375000 ;
        RECT 72.610000 70.585000 72.810000 70.785000 ;
        RECT 72.610000 70.995000 72.810000 71.195000 ;
        RECT 72.610000 71.405000 72.810000 71.605000 ;
        RECT 72.610000 71.815000 72.810000 72.015000 ;
        RECT 72.610000 72.225000 72.810000 72.425000 ;
        RECT 72.610000 72.635000 72.810000 72.835000 ;
        RECT 72.610000 73.045000 72.810000 73.245000 ;
        RECT 72.610000 73.450000 72.810000 73.650000 ;
        RECT 72.610000 73.855000 72.810000 74.055000 ;
        RECT 72.610000 74.260000 72.810000 74.460000 ;
        RECT 72.610000 74.665000 72.810000 74.865000 ;
        RECT 72.610000 75.070000 72.810000 75.270000 ;
        RECT 72.610000 75.475000 72.810000 75.675000 ;
        RECT 72.610000 75.880000 72.810000 76.080000 ;
        RECT 72.610000 76.285000 72.810000 76.485000 ;
        RECT 72.610000 76.690000 72.810000 76.890000 ;
        RECT 72.610000 77.095000 72.810000 77.295000 ;
        RECT 72.610000 77.500000 72.810000 77.700000 ;
        RECT 72.610000 77.905000 72.810000 78.105000 ;
        RECT 72.610000 78.310000 72.810000 78.510000 ;
        RECT 72.610000 78.715000 72.810000 78.915000 ;
        RECT 72.610000 79.120000 72.810000 79.320000 ;
        RECT 72.610000 79.525000 72.810000 79.725000 ;
        RECT 72.610000 79.930000 72.810000 80.130000 ;
        RECT 72.610000 80.335000 72.810000 80.535000 ;
        RECT 72.610000 80.740000 72.810000 80.940000 ;
        RECT 72.610000 81.145000 72.810000 81.345000 ;
        RECT 72.610000 81.550000 72.810000 81.750000 ;
        RECT 72.610000 81.955000 72.810000 82.155000 ;
        RECT 72.610000 82.360000 72.810000 82.560000 ;
        RECT 72.680000 82.855000 72.880000 83.055000 ;
        RECT 72.680000 83.265000 72.880000 83.465000 ;
        RECT 72.680000 83.675000 72.880000 83.875000 ;
        RECT 72.680000 84.085000 72.880000 84.285000 ;
        RECT 72.680000 84.495000 72.880000 84.695000 ;
        RECT 72.680000 84.905000 72.880000 85.105000 ;
        RECT 72.680000 85.315000 72.880000 85.515000 ;
        RECT 72.680000 85.725000 72.880000 85.925000 ;
        RECT 72.680000 86.135000 72.880000 86.335000 ;
        RECT 72.680000 86.545000 72.880000 86.745000 ;
        RECT 72.680000 86.955000 72.880000 87.155000 ;
        RECT 72.680000 87.365000 72.880000 87.565000 ;
        RECT 72.680000 87.775000 72.880000 87.975000 ;
        RECT 72.680000 88.185000 72.880000 88.385000 ;
        RECT 72.680000 88.595000 72.880000 88.795000 ;
        RECT 72.680000 89.005000 72.880000 89.205000 ;
        RECT 72.680000 89.415000 72.880000 89.615000 ;
        RECT 72.680000 89.825000 72.880000 90.025000 ;
        RECT 72.680000 90.235000 72.880000 90.435000 ;
        RECT 72.680000 90.645000 72.880000 90.845000 ;
        RECT 72.680000 91.055000 72.880000 91.255000 ;
        RECT 72.680000 91.465000 72.880000 91.665000 ;
        RECT 72.680000 91.875000 72.880000 92.075000 ;
        RECT 72.680000 92.285000 72.880000 92.485000 ;
        RECT 72.680000 92.695000 72.880000 92.895000 ;
        RECT 72.725000 17.860000 72.925000 18.060000 ;
        RECT 72.725000 18.290000 72.925000 18.490000 ;
        RECT 72.725000 18.720000 72.925000 18.920000 ;
        RECT 72.725000 19.150000 72.925000 19.350000 ;
        RECT 72.725000 19.580000 72.925000 19.780000 ;
        RECT 72.725000 20.010000 72.925000 20.210000 ;
        RECT 72.725000 20.440000 72.925000 20.640000 ;
        RECT 72.725000 20.870000 72.925000 21.070000 ;
        RECT 72.725000 21.300000 72.925000 21.500000 ;
        RECT 72.725000 21.730000 72.925000 21.930000 ;
        RECT 72.725000 22.160000 72.925000 22.360000 ;
        RECT 73.010000 68.125000 73.210000 68.325000 ;
        RECT 73.010000 68.535000 73.210000 68.735000 ;
        RECT 73.010000 68.945000 73.210000 69.145000 ;
        RECT 73.010000 69.355000 73.210000 69.555000 ;
        RECT 73.010000 69.765000 73.210000 69.965000 ;
        RECT 73.010000 70.175000 73.210000 70.375000 ;
        RECT 73.010000 70.585000 73.210000 70.785000 ;
        RECT 73.010000 70.995000 73.210000 71.195000 ;
        RECT 73.010000 71.405000 73.210000 71.605000 ;
        RECT 73.010000 71.815000 73.210000 72.015000 ;
        RECT 73.010000 72.225000 73.210000 72.425000 ;
        RECT 73.010000 72.635000 73.210000 72.835000 ;
        RECT 73.010000 73.045000 73.210000 73.245000 ;
        RECT 73.010000 73.450000 73.210000 73.650000 ;
        RECT 73.010000 73.855000 73.210000 74.055000 ;
        RECT 73.010000 74.260000 73.210000 74.460000 ;
        RECT 73.010000 74.665000 73.210000 74.865000 ;
        RECT 73.010000 75.070000 73.210000 75.270000 ;
        RECT 73.010000 75.475000 73.210000 75.675000 ;
        RECT 73.010000 75.880000 73.210000 76.080000 ;
        RECT 73.010000 76.285000 73.210000 76.485000 ;
        RECT 73.010000 76.690000 73.210000 76.890000 ;
        RECT 73.010000 77.095000 73.210000 77.295000 ;
        RECT 73.010000 77.500000 73.210000 77.700000 ;
        RECT 73.010000 77.905000 73.210000 78.105000 ;
        RECT 73.010000 78.310000 73.210000 78.510000 ;
        RECT 73.010000 78.715000 73.210000 78.915000 ;
        RECT 73.010000 79.120000 73.210000 79.320000 ;
        RECT 73.010000 79.525000 73.210000 79.725000 ;
        RECT 73.010000 79.930000 73.210000 80.130000 ;
        RECT 73.010000 80.335000 73.210000 80.535000 ;
        RECT 73.010000 80.740000 73.210000 80.940000 ;
        RECT 73.010000 81.145000 73.210000 81.345000 ;
        RECT 73.010000 81.550000 73.210000 81.750000 ;
        RECT 73.010000 81.955000 73.210000 82.155000 ;
        RECT 73.010000 82.360000 73.210000 82.560000 ;
        RECT 73.090000 82.855000 73.290000 83.055000 ;
        RECT 73.090000 83.265000 73.290000 83.465000 ;
        RECT 73.090000 83.675000 73.290000 83.875000 ;
        RECT 73.090000 84.085000 73.290000 84.285000 ;
        RECT 73.090000 84.495000 73.290000 84.695000 ;
        RECT 73.090000 84.905000 73.290000 85.105000 ;
        RECT 73.090000 85.315000 73.290000 85.515000 ;
        RECT 73.090000 85.725000 73.290000 85.925000 ;
        RECT 73.090000 86.135000 73.290000 86.335000 ;
        RECT 73.090000 86.545000 73.290000 86.745000 ;
        RECT 73.090000 86.955000 73.290000 87.155000 ;
        RECT 73.090000 87.365000 73.290000 87.565000 ;
        RECT 73.090000 87.775000 73.290000 87.975000 ;
        RECT 73.090000 88.185000 73.290000 88.385000 ;
        RECT 73.090000 88.595000 73.290000 88.795000 ;
        RECT 73.090000 89.005000 73.290000 89.205000 ;
        RECT 73.090000 89.415000 73.290000 89.615000 ;
        RECT 73.090000 89.825000 73.290000 90.025000 ;
        RECT 73.090000 90.235000 73.290000 90.435000 ;
        RECT 73.090000 90.645000 73.290000 90.845000 ;
        RECT 73.090000 91.055000 73.290000 91.255000 ;
        RECT 73.090000 91.465000 73.290000 91.665000 ;
        RECT 73.090000 91.875000 73.290000 92.075000 ;
        RECT 73.090000 92.285000 73.290000 92.485000 ;
        RECT 73.090000 92.695000 73.290000 92.895000 ;
        RECT 73.135000 17.860000 73.335000 18.060000 ;
        RECT 73.135000 18.290000 73.335000 18.490000 ;
        RECT 73.135000 18.720000 73.335000 18.920000 ;
        RECT 73.135000 19.150000 73.335000 19.350000 ;
        RECT 73.135000 19.580000 73.335000 19.780000 ;
        RECT 73.135000 20.010000 73.335000 20.210000 ;
        RECT 73.135000 20.440000 73.335000 20.640000 ;
        RECT 73.135000 20.870000 73.335000 21.070000 ;
        RECT 73.135000 21.300000 73.335000 21.500000 ;
        RECT 73.135000 21.730000 73.335000 21.930000 ;
        RECT 73.135000 22.160000 73.335000 22.360000 ;
        RECT 73.410000 68.125000 73.610000 68.325000 ;
        RECT 73.410000 68.535000 73.610000 68.735000 ;
        RECT 73.410000 68.945000 73.610000 69.145000 ;
        RECT 73.410000 69.355000 73.610000 69.555000 ;
        RECT 73.410000 69.765000 73.610000 69.965000 ;
        RECT 73.410000 70.175000 73.610000 70.375000 ;
        RECT 73.410000 70.585000 73.610000 70.785000 ;
        RECT 73.410000 70.995000 73.610000 71.195000 ;
        RECT 73.410000 71.405000 73.610000 71.605000 ;
        RECT 73.410000 71.815000 73.610000 72.015000 ;
        RECT 73.410000 72.225000 73.610000 72.425000 ;
        RECT 73.410000 72.635000 73.610000 72.835000 ;
        RECT 73.410000 73.045000 73.610000 73.245000 ;
        RECT 73.410000 73.450000 73.610000 73.650000 ;
        RECT 73.410000 73.855000 73.610000 74.055000 ;
        RECT 73.410000 74.260000 73.610000 74.460000 ;
        RECT 73.410000 74.665000 73.610000 74.865000 ;
        RECT 73.410000 75.070000 73.610000 75.270000 ;
        RECT 73.410000 75.475000 73.610000 75.675000 ;
        RECT 73.410000 75.880000 73.610000 76.080000 ;
        RECT 73.410000 76.285000 73.610000 76.485000 ;
        RECT 73.410000 76.690000 73.610000 76.890000 ;
        RECT 73.410000 77.095000 73.610000 77.295000 ;
        RECT 73.410000 77.500000 73.610000 77.700000 ;
        RECT 73.410000 77.905000 73.610000 78.105000 ;
        RECT 73.410000 78.310000 73.610000 78.510000 ;
        RECT 73.410000 78.715000 73.610000 78.915000 ;
        RECT 73.410000 79.120000 73.610000 79.320000 ;
        RECT 73.410000 79.525000 73.610000 79.725000 ;
        RECT 73.410000 79.930000 73.610000 80.130000 ;
        RECT 73.410000 80.335000 73.610000 80.535000 ;
        RECT 73.410000 80.740000 73.610000 80.940000 ;
        RECT 73.410000 81.145000 73.610000 81.345000 ;
        RECT 73.410000 81.550000 73.610000 81.750000 ;
        RECT 73.410000 81.955000 73.610000 82.155000 ;
        RECT 73.410000 82.360000 73.610000 82.560000 ;
        RECT 73.500000 82.855000 73.700000 83.055000 ;
        RECT 73.500000 83.265000 73.700000 83.465000 ;
        RECT 73.500000 83.675000 73.700000 83.875000 ;
        RECT 73.500000 84.085000 73.700000 84.285000 ;
        RECT 73.500000 84.495000 73.700000 84.695000 ;
        RECT 73.500000 84.905000 73.700000 85.105000 ;
        RECT 73.500000 85.315000 73.700000 85.515000 ;
        RECT 73.500000 85.725000 73.700000 85.925000 ;
        RECT 73.500000 86.135000 73.700000 86.335000 ;
        RECT 73.500000 86.545000 73.700000 86.745000 ;
        RECT 73.500000 86.955000 73.700000 87.155000 ;
        RECT 73.500000 87.365000 73.700000 87.565000 ;
        RECT 73.500000 87.775000 73.700000 87.975000 ;
        RECT 73.500000 88.185000 73.700000 88.385000 ;
        RECT 73.500000 88.595000 73.700000 88.795000 ;
        RECT 73.500000 89.005000 73.700000 89.205000 ;
        RECT 73.500000 89.415000 73.700000 89.615000 ;
        RECT 73.500000 89.825000 73.700000 90.025000 ;
        RECT 73.500000 90.235000 73.700000 90.435000 ;
        RECT 73.500000 90.645000 73.700000 90.845000 ;
        RECT 73.500000 91.055000 73.700000 91.255000 ;
        RECT 73.500000 91.465000 73.700000 91.665000 ;
        RECT 73.500000 91.875000 73.700000 92.075000 ;
        RECT 73.500000 92.285000 73.700000 92.485000 ;
        RECT 73.500000 92.695000 73.700000 92.895000 ;
        RECT 73.545000 17.860000 73.745000 18.060000 ;
        RECT 73.545000 18.290000 73.745000 18.490000 ;
        RECT 73.545000 18.720000 73.745000 18.920000 ;
        RECT 73.545000 19.150000 73.745000 19.350000 ;
        RECT 73.545000 19.580000 73.745000 19.780000 ;
        RECT 73.545000 20.010000 73.745000 20.210000 ;
        RECT 73.545000 20.440000 73.745000 20.640000 ;
        RECT 73.545000 20.870000 73.745000 21.070000 ;
        RECT 73.545000 21.300000 73.745000 21.500000 ;
        RECT 73.545000 21.730000 73.745000 21.930000 ;
        RECT 73.545000 22.160000 73.745000 22.360000 ;
        RECT 73.810000 68.125000 74.010000 68.325000 ;
        RECT 73.810000 68.535000 74.010000 68.735000 ;
        RECT 73.810000 68.945000 74.010000 69.145000 ;
        RECT 73.810000 69.355000 74.010000 69.555000 ;
        RECT 73.810000 69.765000 74.010000 69.965000 ;
        RECT 73.810000 70.175000 74.010000 70.375000 ;
        RECT 73.810000 70.585000 74.010000 70.785000 ;
        RECT 73.810000 70.995000 74.010000 71.195000 ;
        RECT 73.810000 71.405000 74.010000 71.605000 ;
        RECT 73.810000 71.815000 74.010000 72.015000 ;
        RECT 73.810000 72.225000 74.010000 72.425000 ;
        RECT 73.810000 72.635000 74.010000 72.835000 ;
        RECT 73.810000 73.045000 74.010000 73.245000 ;
        RECT 73.810000 73.450000 74.010000 73.650000 ;
        RECT 73.810000 73.855000 74.010000 74.055000 ;
        RECT 73.810000 74.260000 74.010000 74.460000 ;
        RECT 73.810000 74.665000 74.010000 74.865000 ;
        RECT 73.810000 75.070000 74.010000 75.270000 ;
        RECT 73.810000 75.475000 74.010000 75.675000 ;
        RECT 73.810000 75.880000 74.010000 76.080000 ;
        RECT 73.810000 76.285000 74.010000 76.485000 ;
        RECT 73.810000 76.690000 74.010000 76.890000 ;
        RECT 73.810000 77.095000 74.010000 77.295000 ;
        RECT 73.810000 77.500000 74.010000 77.700000 ;
        RECT 73.810000 77.905000 74.010000 78.105000 ;
        RECT 73.810000 78.310000 74.010000 78.510000 ;
        RECT 73.810000 78.715000 74.010000 78.915000 ;
        RECT 73.810000 79.120000 74.010000 79.320000 ;
        RECT 73.810000 79.525000 74.010000 79.725000 ;
        RECT 73.810000 79.930000 74.010000 80.130000 ;
        RECT 73.810000 80.335000 74.010000 80.535000 ;
        RECT 73.810000 80.740000 74.010000 80.940000 ;
        RECT 73.810000 81.145000 74.010000 81.345000 ;
        RECT 73.810000 81.550000 74.010000 81.750000 ;
        RECT 73.810000 81.955000 74.010000 82.155000 ;
        RECT 73.810000 82.360000 74.010000 82.560000 ;
        RECT 73.910000 82.855000 74.110000 83.055000 ;
        RECT 73.910000 83.265000 74.110000 83.465000 ;
        RECT 73.910000 83.675000 74.110000 83.875000 ;
        RECT 73.910000 84.085000 74.110000 84.285000 ;
        RECT 73.910000 84.495000 74.110000 84.695000 ;
        RECT 73.910000 84.905000 74.110000 85.105000 ;
        RECT 73.910000 85.315000 74.110000 85.515000 ;
        RECT 73.910000 85.725000 74.110000 85.925000 ;
        RECT 73.910000 86.135000 74.110000 86.335000 ;
        RECT 73.910000 86.545000 74.110000 86.745000 ;
        RECT 73.910000 86.955000 74.110000 87.155000 ;
        RECT 73.910000 87.365000 74.110000 87.565000 ;
        RECT 73.910000 87.775000 74.110000 87.975000 ;
        RECT 73.910000 88.185000 74.110000 88.385000 ;
        RECT 73.910000 88.595000 74.110000 88.795000 ;
        RECT 73.910000 89.005000 74.110000 89.205000 ;
        RECT 73.910000 89.415000 74.110000 89.615000 ;
        RECT 73.910000 89.825000 74.110000 90.025000 ;
        RECT 73.910000 90.235000 74.110000 90.435000 ;
        RECT 73.910000 90.645000 74.110000 90.845000 ;
        RECT 73.910000 91.055000 74.110000 91.255000 ;
        RECT 73.910000 91.465000 74.110000 91.665000 ;
        RECT 73.910000 91.875000 74.110000 92.075000 ;
        RECT 73.910000 92.285000 74.110000 92.485000 ;
        RECT 73.910000 92.695000 74.110000 92.895000 ;
        RECT 73.955000 17.860000 74.155000 18.060000 ;
        RECT 73.955000 18.290000 74.155000 18.490000 ;
        RECT 73.955000 18.720000 74.155000 18.920000 ;
        RECT 73.955000 19.150000 74.155000 19.350000 ;
        RECT 73.955000 19.580000 74.155000 19.780000 ;
        RECT 73.955000 20.010000 74.155000 20.210000 ;
        RECT 73.955000 20.440000 74.155000 20.640000 ;
        RECT 73.955000 20.870000 74.155000 21.070000 ;
        RECT 73.955000 21.300000 74.155000 21.500000 ;
        RECT 73.955000 21.730000 74.155000 21.930000 ;
        RECT 73.955000 22.160000 74.155000 22.360000 ;
        RECT 74.210000 68.125000 74.410000 68.325000 ;
        RECT 74.210000 68.535000 74.410000 68.735000 ;
        RECT 74.210000 68.945000 74.410000 69.145000 ;
        RECT 74.210000 69.355000 74.410000 69.555000 ;
        RECT 74.210000 69.765000 74.410000 69.965000 ;
        RECT 74.210000 70.175000 74.410000 70.375000 ;
        RECT 74.210000 70.585000 74.410000 70.785000 ;
        RECT 74.210000 70.995000 74.410000 71.195000 ;
        RECT 74.210000 71.405000 74.410000 71.605000 ;
        RECT 74.210000 71.815000 74.410000 72.015000 ;
        RECT 74.210000 72.225000 74.410000 72.425000 ;
        RECT 74.210000 72.635000 74.410000 72.835000 ;
        RECT 74.210000 73.045000 74.410000 73.245000 ;
        RECT 74.210000 73.450000 74.410000 73.650000 ;
        RECT 74.210000 73.855000 74.410000 74.055000 ;
        RECT 74.210000 74.260000 74.410000 74.460000 ;
        RECT 74.210000 74.665000 74.410000 74.865000 ;
        RECT 74.210000 75.070000 74.410000 75.270000 ;
        RECT 74.210000 75.475000 74.410000 75.675000 ;
        RECT 74.210000 75.880000 74.410000 76.080000 ;
        RECT 74.210000 76.285000 74.410000 76.485000 ;
        RECT 74.210000 76.690000 74.410000 76.890000 ;
        RECT 74.210000 77.095000 74.410000 77.295000 ;
        RECT 74.210000 77.500000 74.410000 77.700000 ;
        RECT 74.210000 77.905000 74.410000 78.105000 ;
        RECT 74.210000 78.310000 74.410000 78.510000 ;
        RECT 74.210000 78.715000 74.410000 78.915000 ;
        RECT 74.210000 79.120000 74.410000 79.320000 ;
        RECT 74.210000 79.525000 74.410000 79.725000 ;
        RECT 74.210000 79.930000 74.410000 80.130000 ;
        RECT 74.210000 80.335000 74.410000 80.535000 ;
        RECT 74.210000 80.740000 74.410000 80.940000 ;
        RECT 74.210000 81.145000 74.410000 81.345000 ;
        RECT 74.210000 81.550000 74.410000 81.750000 ;
        RECT 74.210000 81.955000 74.410000 82.155000 ;
        RECT 74.210000 82.360000 74.410000 82.560000 ;
        RECT 74.320000 82.855000 74.520000 83.055000 ;
        RECT 74.320000 83.265000 74.520000 83.465000 ;
        RECT 74.320000 83.675000 74.520000 83.875000 ;
        RECT 74.320000 84.085000 74.520000 84.285000 ;
        RECT 74.320000 84.495000 74.520000 84.695000 ;
        RECT 74.320000 84.905000 74.520000 85.105000 ;
        RECT 74.320000 85.315000 74.520000 85.515000 ;
        RECT 74.320000 85.725000 74.520000 85.925000 ;
        RECT 74.320000 86.135000 74.520000 86.335000 ;
        RECT 74.320000 86.545000 74.520000 86.745000 ;
        RECT 74.320000 86.955000 74.520000 87.155000 ;
        RECT 74.320000 87.365000 74.520000 87.565000 ;
        RECT 74.320000 87.775000 74.520000 87.975000 ;
        RECT 74.320000 88.185000 74.520000 88.385000 ;
        RECT 74.320000 88.595000 74.520000 88.795000 ;
        RECT 74.320000 89.005000 74.520000 89.205000 ;
        RECT 74.320000 89.415000 74.520000 89.615000 ;
        RECT 74.320000 89.825000 74.520000 90.025000 ;
        RECT 74.320000 90.235000 74.520000 90.435000 ;
        RECT 74.320000 90.645000 74.520000 90.845000 ;
        RECT 74.320000 91.055000 74.520000 91.255000 ;
        RECT 74.320000 91.465000 74.520000 91.665000 ;
        RECT 74.320000 91.875000 74.520000 92.075000 ;
        RECT 74.320000 92.285000 74.520000 92.485000 ;
        RECT 74.320000 92.695000 74.520000 92.895000 ;
        RECT 74.365000 17.860000 74.565000 18.060000 ;
        RECT 74.365000 18.290000 74.565000 18.490000 ;
        RECT 74.365000 18.720000 74.565000 18.920000 ;
        RECT 74.365000 19.150000 74.565000 19.350000 ;
        RECT 74.365000 19.580000 74.565000 19.780000 ;
        RECT 74.365000 20.010000 74.565000 20.210000 ;
        RECT 74.365000 20.440000 74.565000 20.640000 ;
        RECT 74.365000 20.870000 74.565000 21.070000 ;
        RECT 74.365000 21.300000 74.565000 21.500000 ;
        RECT 74.365000 21.730000 74.565000 21.930000 ;
        RECT 74.365000 22.160000 74.565000 22.360000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.600000 62.090000 24.500000 66.530000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 62.090000 74.655000 66.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 24.475000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.690000 62.160000  0.890000 62.360000 ;
        RECT  0.690000 62.570000  0.890000 62.770000 ;
        RECT  0.690000 62.980000  0.890000 63.180000 ;
        RECT  0.690000 63.390000  0.890000 63.590000 ;
        RECT  0.690000 63.800000  0.890000 64.000000 ;
        RECT  0.690000 64.210000  0.890000 64.410000 ;
        RECT  0.690000 64.620000  0.890000 64.820000 ;
        RECT  0.690000 65.030000  0.890000 65.230000 ;
        RECT  0.690000 65.440000  0.890000 65.640000 ;
        RECT  0.690000 65.850000  0.890000 66.050000 ;
        RECT  0.690000 66.260000  0.890000 66.460000 ;
        RECT  1.095000 62.160000  1.295000 62.360000 ;
        RECT  1.095000 62.570000  1.295000 62.770000 ;
        RECT  1.095000 62.980000  1.295000 63.180000 ;
        RECT  1.095000 63.390000  1.295000 63.590000 ;
        RECT  1.095000 63.800000  1.295000 64.000000 ;
        RECT  1.095000 64.210000  1.295000 64.410000 ;
        RECT  1.095000 64.620000  1.295000 64.820000 ;
        RECT  1.095000 65.030000  1.295000 65.230000 ;
        RECT  1.095000 65.440000  1.295000 65.640000 ;
        RECT  1.095000 65.850000  1.295000 66.050000 ;
        RECT  1.095000 66.260000  1.295000 66.460000 ;
        RECT  1.500000 62.160000  1.700000 62.360000 ;
        RECT  1.500000 62.570000  1.700000 62.770000 ;
        RECT  1.500000 62.980000  1.700000 63.180000 ;
        RECT  1.500000 63.390000  1.700000 63.590000 ;
        RECT  1.500000 63.800000  1.700000 64.000000 ;
        RECT  1.500000 64.210000  1.700000 64.410000 ;
        RECT  1.500000 64.620000  1.700000 64.820000 ;
        RECT  1.500000 65.030000  1.700000 65.230000 ;
        RECT  1.500000 65.440000  1.700000 65.640000 ;
        RECT  1.500000 65.850000  1.700000 66.050000 ;
        RECT  1.500000 66.260000  1.700000 66.460000 ;
        RECT  1.905000 62.160000  2.105000 62.360000 ;
        RECT  1.905000 62.570000  2.105000 62.770000 ;
        RECT  1.905000 62.980000  2.105000 63.180000 ;
        RECT  1.905000 63.390000  2.105000 63.590000 ;
        RECT  1.905000 63.800000  2.105000 64.000000 ;
        RECT  1.905000 64.210000  2.105000 64.410000 ;
        RECT  1.905000 64.620000  2.105000 64.820000 ;
        RECT  1.905000 65.030000  2.105000 65.230000 ;
        RECT  1.905000 65.440000  2.105000 65.640000 ;
        RECT  1.905000 65.850000  2.105000 66.050000 ;
        RECT  1.905000 66.260000  2.105000 66.460000 ;
        RECT  2.310000 62.160000  2.510000 62.360000 ;
        RECT  2.310000 62.570000  2.510000 62.770000 ;
        RECT  2.310000 62.980000  2.510000 63.180000 ;
        RECT  2.310000 63.390000  2.510000 63.590000 ;
        RECT  2.310000 63.800000  2.510000 64.000000 ;
        RECT  2.310000 64.210000  2.510000 64.410000 ;
        RECT  2.310000 64.620000  2.510000 64.820000 ;
        RECT  2.310000 65.030000  2.510000 65.230000 ;
        RECT  2.310000 65.440000  2.510000 65.640000 ;
        RECT  2.310000 65.850000  2.510000 66.050000 ;
        RECT  2.310000 66.260000  2.510000 66.460000 ;
        RECT  2.715000 62.160000  2.915000 62.360000 ;
        RECT  2.715000 62.570000  2.915000 62.770000 ;
        RECT  2.715000 62.980000  2.915000 63.180000 ;
        RECT  2.715000 63.390000  2.915000 63.590000 ;
        RECT  2.715000 63.800000  2.915000 64.000000 ;
        RECT  2.715000 64.210000  2.915000 64.410000 ;
        RECT  2.715000 64.620000  2.915000 64.820000 ;
        RECT  2.715000 65.030000  2.915000 65.230000 ;
        RECT  2.715000 65.440000  2.915000 65.640000 ;
        RECT  2.715000 65.850000  2.915000 66.050000 ;
        RECT  2.715000 66.260000  2.915000 66.460000 ;
        RECT  3.120000 62.160000  3.320000 62.360000 ;
        RECT  3.120000 62.570000  3.320000 62.770000 ;
        RECT  3.120000 62.980000  3.320000 63.180000 ;
        RECT  3.120000 63.390000  3.320000 63.590000 ;
        RECT  3.120000 63.800000  3.320000 64.000000 ;
        RECT  3.120000 64.210000  3.320000 64.410000 ;
        RECT  3.120000 64.620000  3.320000 64.820000 ;
        RECT  3.120000 65.030000  3.320000 65.230000 ;
        RECT  3.120000 65.440000  3.320000 65.640000 ;
        RECT  3.120000 65.850000  3.320000 66.050000 ;
        RECT  3.120000 66.260000  3.320000 66.460000 ;
        RECT  3.525000 62.160000  3.725000 62.360000 ;
        RECT  3.525000 62.570000  3.725000 62.770000 ;
        RECT  3.525000 62.980000  3.725000 63.180000 ;
        RECT  3.525000 63.390000  3.725000 63.590000 ;
        RECT  3.525000 63.800000  3.725000 64.000000 ;
        RECT  3.525000 64.210000  3.725000 64.410000 ;
        RECT  3.525000 64.620000  3.725000 64.820000 ;
        RECT  3.525000 65.030000  3.725000 65.230000 ;
        RECT  3.525000 65.440000  3.725000 65.640000 ;
        RECT  3.525000 65.850000  3.725000 66.050000 ;
        RECT  3.525000 66.260000  3.725000 66.460000 ;
        RECT  3.930000 62.160000  4.130000 62.360000 ;
        RECT  3.930000 62.570000  4.130000 62.770000 ;
        RECT  3.930000 62.980000  4.130000 63.180000 ;
        RECT  3.930000 63.390000  4.130000 63.590000 ;
        RECT  3.930000 63.800000  4.130000 64.000000 ;
        RECT  3.930000 64.210000  4.130000 64.410000 ;
        RECT  3.930000 64.620000  4.130000 64.820000 ;
        RECT  3.930000 65.030000  4.130000 65.230000 ;
        RECT  3.930000 65.440000  4.130000 65.640000 ;
        RECT  3.930000 65.850000  4.130000 66.050000 ;
        RECT  3.930000 66.260000  4.130000 66.460000 ;
        RECT  4.335000 62.160000  4.535000 62.360000 ;
        RECT  4.335000 62.570000  4.535000 62.770000 ;
        RECT  4.335000 62.980000  4.535000 63.180000 ;
        RECT  4.335000 63.390000  4.535000 63.590000 ;
        RECT  4.335000 63.800000  4.535000 64.000000 ;
        RECT  4.335000 64.210000  4.535000 64.410000 ;
        RECT  4.335000 64.620000  4.535000 64.820000 ;
        RECT  4.335000 65.030000  4.535000 65.230000 ;
        RECT  4.335000 65.440000  4.535000 65.640000 ;
        RECT  4.335000 65.850000  4.535000 66.050000 ;
        RECT  4.335000 66.260000  4.535000 66.460000 ;
        RECT  4.740000 62.160000  4.940000 62.360000 ;
        RECT  4.740000 62.570000  4.940000 62.770000 ;
        RECT  4.740000 62.980000  4.940000 63.180000 ;
        RECT  4.740000 63.390000  4.940000 63.590000 ;
        RECT  4.740000 63.800000  4.940000 64.000000 ;
        RECT  4.740000 64.210000  4.940000 64.410000 ;
        RECT  4.740000 64.620000  4.940000 64.820000 ;
        RECT  4.740000 65.030000  4.940000 65.230000 ;
        RECT  4.740000 65.440000  4.940000 65.640000 ;
        RECT  4.740000 65.850000  4.940000 66.050000 ;
        RECT  4.740000 66.260000  4.940000 66.460000 ;
        RECT  5.145000 62.160000  5.345000 62.360000 ;
        RECT  5.145000 62.570000  5.345000 62.770000 ;
        RECT  5.145000 62.980000  5.345000 63.180000 ;
        RECT  5.145000 63.390000  5.345000 63.590000 ;
        RECT  5.145000 63.800000  5.345000 64.000000 ;
        RECT  5.145000 64.210000  5.345000 64.410000 ;
        RECT  5.145000 64.620000  5.345000 64.820000 ;
        RECT  5.145000 65.030000  5.345000 65.230000 ;
        RECT  5.145000 65.440000  5.345000 65.640000 ;
        RECT  5.145000 65.850000  5.345000 66.050000 ;
        RECT  5.145000 66.260000  5.345000 66.460000 ;
        RECT  5.550000 62.160000  5.750000 62.360000 ;
        RECT  5.550000 62.570000  5.750000 62.770000 ;
        RECT  5.550000 62.980000  5.750000 63.180000 ;
        RECT  5.550000 63.390000  5.750000 63.590000 ;
        RECT  5.550000 63.800000  5.750000 64.000000 ;
        RECT  5.550000 64.210000  5.750000 64.410000 ;
        RECT  5.550000 64.620000  5.750000 64.820000 ;
        RECT  5.550000 65.030000  5.750000 65.230000 ;
        RECT  5.550000 65.440000  5.750000 65.640000 ;
        RECT  5.550000 65.850000  5.750000 66.050000 ;
        RECT  5.550000 66.260000  5.750000 66.460000 ;
        RECT  5.955000 62.160000  6.155000 62.360000 ;
        RECT  5.955000 62.570000  6.155000 62.770000 ;
        RECT  5.955000 62.980000  6.155000 63.180000 ;
        RECT  5.955000 63.390000  6.155000 63.590000 ;
        RECT  5.955000 63.800000  6.155000 64.000000 ;
        RECT  5.955000 64.210000  6.155000 64.410000 ;
        RECT  5.955000 64.620000  6.155000 64.820000 ;
        RECT  5.955000 65.030000  6.155000 65.230000 ;
        RECT  5.955000 65.440000  6.155000 65.640000 ;
        RECT  5.955000 65.850000  6.155000 66.050000 ;
        RECT  5.955000 66.260000  6.155000 66.460000 ;
        RECT  6.360000 62.160000  6.560000 62.360000 ;
        RECT  6.360000 62.570000  6.560000 62.770000 ;
        RECT  6.360000 62.980000  6.560000 63.180000 ;
        RECT  6.360000 63.390000  6.560000 63.590000 ;
        RECT  6.360000 63.800000  6.560000 64.000000 ;
        RECT  6.360000 64.210000  6.560000 64.410000 ;
        RECT  6.360000 64.620000  6.560000 64.820000 ;
        RECT  6.360000 65.030000  6.560000 65.230000 ;
        RECT  6.360000 65.440000  6.560000 65.640000 ;
        RECT  6.360000 65.850000  6.560000 66.050000 ;
        RECT  6.360000 66.260000  6.560000 66.460000 ;
        RECT  6.765000 62.160000  6.965000 62.360000 ;
        RECT  6.765000 62.570000  6.965000 62.770000 ;
        RECT  6.765000 62.980000  6.965000 63.180000 ;
        RECT  6.765000 63.390000  6.965000 63.590000 ;
        RECT  6.765000 63.800000  6.965000 64.000000 ;
        RECT  6.765000 64.210000  6.965000 64.410000 ;
        RECT  6.765000 64.620000  6.965000 64.820000 ;
        RECT  6.765000 65.030000  6.965000 65.230000 ;
        RECT  6.765000 65.440000  6.965000 65.640000 ;
        RECT  6.765000 65.850000  6.965000 66.050000 ;
        RECT  6.765000 66.260000  6.965000 66.460000 ;
        RECT  7.170000 62.160000  7.370000 62.360000 ;
        RECT  7.170000 62.570000  7.370000 62.770000 ;
        RECT  7.170000 62.980000  7.370000 63.180000 ;
        RECT  7.170000 63.390000  7.370000 63.590000 ;
        RECT  7.170000 63.800000  7.370000 64.000000 ;
        RECT  7.170000 64.210000  7.370000 64.410000 ;
        RECT  7.170000 64.620000  7.370000 64.820000 ;
        RECT  7.170000 65.030000  7.370000 65.230000 ;
        RECT  7.170000 65.440000  7.370000 65.640000 ;
        RECT  7.170000 65.850000  7.370000 66.050000 ;
        RECT  7.170000 66.260000  7.370000 66.460000 ;
        RECT  7.575000 62.160000  7.775000 62.360000 ;
        RECT  7.575000 62.570000  7.775000 62.770000 ;
        RECT  7.575000 62.980000  7.775000 63.180000 ;
        RECT  7.575000 63.390000  7.775000 63.590000 ;
        RECT  7.575000 63.800000  7.775000 64.000000 ;
        RECT  7.575000 64.210000  7.775000 64.410000 ;
        RECT  7.575000 64.620000  7.775000 64.820000 ;
        RECT  7.575000 65.030000  7.775000 65.230000 ;
        RECT  7.575000 65.440000  7.775000 65.640000 ;
        RECT  7.575000 65.850000  7.775000 66.050000 ;
        RECT  7.575000 66.260000  7.775000 66.460000 ;
        RECT  7.980000 62.160000  8.180000 62.360000 ;
        RECT  7.980000 62.570000  8.180000 62.770000 ;
        RECT  7.980000 62.980000  8.180000 63.180000 ;
        RECT  7.980000 63.390000  8.180000 63.590000 ;
        RECT  7.980000 63.800000  8.180000 64.000000 ;
        RECT  7.980000 64.210000  8.180000 64.410000 ;
        RECT  7.980000 64.620000  8.180000 64.820000 ;
        RECT  7.980000 65.030000  8.180000 65.230000 ;
        RECT  7.980000 65.440000  8.180000 65.640000 ;
        RECT  7.980000 65.850000  8.180000 66.050000 ;
        RECT  7.980000 66.260000  8.180000 66.460000 ;
        RECT  8.385000 62.160000  8.585000 62.360000 ;
        RECT  8.385000 62.570000  8.585000 62.770000 ;
        RECT  8.385000 62.980000  8.585000 63.180000 ;
        RECT  8.385000 63.390000  8.585000 63.590000 ;
        RECT  8.385000 63.800000  8.585000 64.000000 ;
        RECT  8.385000 64.210000  8.585000 64.410000 ;
        RECT  8.385000 64.620000  8.585000 64.820000 ;
        RECT  8.385000 65.030000  8.585000 65.230000 ;
        RECT  8.385000 65.440000  8.585000 65.640000 ;
        RECT  8.385000 65.850000  8.585000 66.050000 ;
        RECT  8.385000 66.260000  8.585000 66.460000 ;
        RECT  8.790000 62.160000  8.990000 62.360000 ;
        RECT  8.790000 62.570000  8.990000 62.770000 ;
        RECT  8.790000 62.980000  8.990000 63.180000 ;
        RECT  8.790000 63.390000  8.990000 63.590000 ;
        RECT  8.790000 63.800000  8.990000 64.000000 ;
        RECT  8.790000 64.210000  8.990000 64.410000 ;
        RECT  8.790000 64.620000  8.990000 64.820000 ;
        RECT  8.790000 65.030000  8.990000 65.230000 ;
        RECT  8.790000 65.440000  8.990000 65.640000 ;
        RECT  8.790000 65.850000  8.990000 66.050000 ;
        RECT  8.790000 66.260000  8.990000 66.460000 ;
        RECT  9.195000 62.160000  9.395000 62.360000 ;
        RECT  9.195000 62.570000  9.395000 62.770000 ;
        RECT  9.195000 62.980000  9.395000 63.180000 ;
        RECT  9.195000 63.390000  9.395000 63.590000 ;
        RECT  9.195000 63.800000  9.395000 64.000000 ;
        RECT  9.195000 64.210000  9.395000 64.410000 ;
        RECT  9.195000 64.620000  9.395000 64.820000 ;
        RECT  9.195000 65.030000  9.395000 65.230000 ;
        RECT  9.195000 65.440000  9.395000 65.640000 ;
        RECT  9.195000 65.850000  9.395000 66.050000 ;
        RECT  9.195000 66.260000  9.395000 66.460000 ;
        RECT  9.600000 62.160000  9.800000 62.360000 ;
        RECT  9.600000 62.570000  9.800000 62.770000 ;
        RECT  9.600000 62.980000  9.800000 63.180000 ;
        RECT  9.600000 63.390000  9.800000 63.590000 ;
        RECT  9.600000 63.800000  9.800000 64.000000 ;
        RECT  9.600000 64.210000  9.800000 64.410000 ;
        RECT  9.600000 64.620000  9.800000 64.820000 ;
        RECT  9.600000 65.030000  9.800000 65.230000 ;
        RECT  9.600000 65.440000  9.800000 65.640000 ;
        RECT  9.600000 65.850000  9.800000 66.050000 ;
        RECT  9.600000 66.260000  9.800000 66.460000 ;
        RECT 10.005000 62.160000 10.205000 62.360000 ;
        RECT 10.005000 62.570000 10.205000 62.770000 ;
        RECT 10.005000 62.980000 10.205000 63.180000 ;
        RECT 10.005000 63.390000 10.205000 63.590000 ;
        RECT 10.005000 63.800000 10.205000 64.000000 ;
        RECT 10.005000 64.210000 10.205000 64.410000 ;
        RECT 10.005000 64.620000 10.205000 64.820000 ;
        RECT 10.005000 65.030000 10.205000 65.230000 ;
        RECT 10.005000 65.440000 10.205000 65.640000 ;
        RECT 10.005000 65.850000 10.205000 66.050000 ;
        RECT 10.005000 66.260000 10.205000 66.460000 ;
        RECT 10.410000 62.160000 10.610000 62.360000 ;
        RECT 10.410000 62.570000 10.610000 62.770000 ;
        RECT 10.410000 62.980000 10.610000 63.180000 ;
        RECT 10.410000 63.390000 10.610000 63.590000 ;
        RECT 10.410000 63.800000 10.610000 64.000000 ;
        RECT 10.410000 64.210000 10.610000 64.410000 ;
        RECT 10.410000 64.620000 10.610000 64.820000 ;
        RECT 10.410000 65.030000 10.610000 65.230000 ;
        RECT 10.410000 65.440000 10.610000 65.640000 ;
        RECT 10.410000 65.850000 10.610000 66.050000 ;
        RECT 10.410000 66.260000 10.610000 66.460000 ;
        RECT 10.815000 62.160000 11.015000 62.360000 ;
        RECT 10.815000 62.570000 11.015000 62.770000 ;
        RECT 10.815000 62.980000 11.015000 63.180000 ;
        RECT 10.815000 63.390000 11.015000 63.590000 ;
        RECT 10.815000 63.800000 11.015000 64.000000 ;
        RECT 10.815000 64.210000 11.015000 64.410000 ;
        RECT 10.815000 64.620000 11.015000 64.820000 ;
        RECT 10.815000 65.030000 11.015000 65.230000 ;
        RECT 10.815000 65.440000 11.015000 65.640000 ;
        RECT 10.815000 65.850000 11.015000 66.050000 ;
        RECT 10.815000 66.260000 11.015000 66.460000 ;
        RECT 11.220000 62.160000 11.420000 62.360000 ;
        RECT 11.220000 62.570000 11.420000 62.770000 ;
        RECT 11.220000 62.980000 11.420000 63.180000 ;
        RECT 11.220000 63.390000 11.420000 63.590000 ;
        RECT 11.220000 63.800000 11.420000 64.000000 ;
        RECT 11.220000 64.210000 11.420000 64.410000 ;
        RECT 11.220000 64.620000 11.420000 64.820000 ;
        RECT 11.220000 65.030000 11.420000 65.230000 ;
        RECT 11.220000 65.440000 11.420000 65.640000 ;
        RECT 11.220000 65.850000 11.420000 66.050000 ;
        RECT 11.220000 66.260000 11.420000 66.460000 ;
        RECT 11.625000 62.160000 11.825000 62.360000 ;
        RECT 11.625000 62.570000 11.825000 62.770000 ;
        RECT 11.625000 62.980000 11.825000 63.180000 ;
        RECT 11.625000 63.390000 11.825000 63.590000 ;
        RECT 11.625000 63.800000 11.825000 64.000000 ;
        RECT 11.625000 64.210000 11.825000 64.410000 ;
        RECT 11.625000 64.620000 11.825000 64.820000 ;
        RECT 11.625000 65.030000 11.825000 65.230000 ;
        RECT 11.625000 65.440000 11.825000 65.640000 ;
        RECT 11.625000 65.850000 11.825000 66.050000 ;
        RECT 11.625000 66.260000 11.825000 66.460000 ;
        RECT 12.030000 62.160000 12.230000 62.360000 ;
        RECT 12.030000 62.570000 12.230000 62.770000 ;
        RECT 12.030000 62.980000 12.230000 63.180000 ;
        RECT 12.030000 63.390000 12.230000 63.590000 ;
        RECT 12.030000 63.800000 12.230000 64.000000 ;
        RECT 12.030000 64.210000 12.230000 64.410000 ;
        RECT 12.030000 64.620000 12.230000 64.820000 ;
        RECT 12.030000 65.030000 12.230000 65.230000 ;
        RECT 12.030000 65.440000 12.230000 65.640000 ;
        RECT 12.030000 65.850000 12.230000 66.050000 ;
        RECT 12.030000 66.260000 12.230000 66.460000 ;
        RECT 12.435000 62.160000 12.635000 62.360000 ;
        RECT 12.435000 62.570000 12.635000 62.770000 ;
        RECT 12.435000 62.980000 12.635000 63.180000 ;
        RECT 12.435000 63.390000 12.635000 63.590000 ;
        RECT 12.435000 63.800000 12.635000 64.000000 ;
        RECT 12.435000 64.210000 12.635000 64.410000 ;
        RECT 12.435000 64.620000 12.635000 64.820000 ;
        RECT 12.435000 65.030000 12.635000 65.230000 ;
        RECT 12.435000 65.440000 12.635000 65.640000 ;
        RECT 12.435000 65.850000 12.635000 66.050000 ;
        RECT 12.435000 66.260000 12.635000 66.460000 ;
        RECT 12.840000 62.160000 13.040000 62.360000 ;
        RECT 12.840000 62.570000 13.040000 62.770000 ;
        RECT 12.840000 62.980000 13.040000 63.180000 ;
        RECT 12.840000 63.390000 13.040000 63.590000 ;
        RECT 12.840000 63.800000 13.040000 64.000000 ;
        RECT 12.840000 64.210000 13.040000 64.410000 ;
        RECT 12.840000 64.620000 13.040000 64.820000 ;
        RECT 12.840000 65.030000 13.040000 65.230000 ;
        RECT 12.840000 65.440000 13.040000 65.640000 ;
        RECT 12.840000 65.850000 13.040000 66.050000 ;
        RECT 12.840000 66.260000 13.040000 66.460000 ;
        RECT 13.245000 62.160000 13.445000 62.360000 ;
        RECT 13.245000 62.570000 13.445000 62.770000 ;
        RECT 13.245000 62.980000 13.445000 63.180000 ;
        RECT 13.245000 63.390000 13.445000 63.590000 ;
        RECT 13.245000 63.800000 13.445000 64.000000 ;
        RECT 13.245000 64.210000 13.445000 64.410000 ;
        RECT 13.245000 64.620000 13.445000 64.820000 ;
        RECT 13.245000 65.030000 13.445000 65.230000 ;
        RECT 13.245000 65.440000 13.445000 65.640000 ;
        RECT 13.245000 65.850000 13.445000 66.050000 ;
        RECT 13.245000 66.260000 13.445000 66.460000 ;
        RECT 13.650000 62.160000 13.850000 62.360000 ;
        RECT 13.650000 62.570000 13.850000 62.770000 ;
        RECT 13.650000 62.980000 13.850000 63.180000 ;
        RECT 13.650000 63.390000 13.850000 63.590000 ;
        RECT 13.650000 63.800000 13.850000 64.000000 ;
        RECT 13.650000 64.210000 13.850000 64.410000 ;
        RECT 13.650000 64.620000 13.850000 64.820000 ;
        RECT 13.650000 65.030000 13.850000 65.230000 ;
        RECT 13.650000 65.440000 13.850000 65.640000 ;
        RECT 13.650000 65.850000 13.850000 66.050000 ;
        RECT 13.650000 66.260000 13.850000 66.460000 ;
        RECT 14.055000 62.160000 14.255000 62.360000 ;
        RECT 14.055000 62.570000 14.255000 62.770000 ;
        RECT 14.055000 62.980000 14.255000 63.180000 ;
        RECT 14.055000 63.390000 14.255000 63.590000 ;
        RECT 14.055000 63.800000 14.255000 64.000000 ;
        RECT 14.055000 64.210000 14.255000 64.410000 ;
        RECT 14.055000 64.620000 14.255000 64.820000 ;
        RECT 14.055000 65.030000 14.255000 65.230000 ;
        RECT 14.055000 65.440000 14.255000 65.640000 ;
        RECT 14.055000 65.850000 14.255000 66.050000 ;
        RECT 14.055000 66.260000 14.255000 66.460000 ;
        RECT 14.460000 62.160000 14.660000 62.360000 ;
        RECT 14.460000 62.570000 14.660000 62.770000 ;
        RECT 14.460000 62.980000 14.660000 63.180000 ;
        RECT 14.460000 63.390000 14.660000 63.590000 ;
        RECT 14.460000 63.800000 14.660000 64.000000 ;
        RECT 14.460000 64.210000 14.660000 64.410000 ;
        RECT 14.460000 64.620000 14.660000 64.820000 ;
        RECT 14.460000 65.030000 14.660000 65.230000 ;
        RECT 14.460000 65.440000 14.660000 65.640000 ;
        RECT 14.460000 65.850000 14.660000 66.050000 ;
        RECT 14.460000 66.260000 14.660000 66.460000 ;
        RECT 14.865000 62.160000 15.065000 62.360000 ;
        RECT 14.865000 62.570000 15.065000 62.770000 ;
        RECT 14.865000 62.980000 15.065000 63.180000 ;
        RECT 14.865000 63.390000 15.065000 63.590000 ;
        RECT 14.865000 63.800000 15.065000 64.000000 ;
        RECT 14.865000 64.210000 15.065000 64.410000 ;
        RECT 14.865000 64.620000 15.065000 64.820000 ;
        RECT 14.865000 65.030000 15.065000 65.230000 ;
        RECT 14.865000 65.440000 15.065000 65.640000 ;
        RECT 14.865000 65.850000 15.065000 66.050000 ;
        RECT 14.865000 66.260000 15.065000 66.460000 ;
        RECT 15.270000 62.160000 15.470000 62.360000 ;
        RECT 15.270000 62.570000 15.470000 62.770000 ;
        RECT 15.270000 62.980000 15.470000 63.180000 ;
        RECT 15.270000 63.390000 15.470000 63.590000 ;
        RECT 15.270000 63.800000 15.470000 64.000000 ;
        RECT 15.270000 64.210000 15.470000 64.410000 ;
        RECT 15.270000 64.620000 15.470000 64.820000 ;
        RECT 15.270000 65.030000 15.470000 65.230000 ;
        RECT 15.270000 65.440000 15.470000 65.640000 ;
        RECT 15.270000 65.850000 15.470000 66.050000 ;
        RECT 15.270000 66.260000 15.470000 66.460000 ;
        RECT 15.675000 62.160000 15.875000 62.360000 ;
        RECT 15.675000 62.570000 15.875000 62.770000 ;
        RECT 15.675000 62.980000 15.875000 63.180000 ;
        RECT 15.675000 63.390000 15.875000 63.590000 ;
        RECT 15.675000 63.800000 15.875000 64.000000 ;
        RECT 15.675000 64.210000 15.875000 64.410000 ;
        RECT 15.675000 64.620000 15.875000 64.820000 ;
        RECT 15.675000 65.030000 15.875000 65.230000 ;
        RECT 15.675000 65.440000 15.875000 65.640000 ;
        RECT 15.675000 65.850000 15.875000 66.050000 ;
        RECT 15.675000 66.260000 15.875000 66.460000 ;
        RECT 16.080000 62.160000 16.280000 62.360000 ;
        RECT 16.080000 62.570000 16.280000 62.770000 ;
        RECT 16.080000 62.980000 16.280000 63.180000 ;
        RECT 16.080000 63.390000 16.280000 63.590000 ;
        RECT 16.080000 63.800000 16.280000 64.000000 ;
        RECT 16.080000 64.210000 16.280000 64.410000 ;
        RECT 16.080000 64.620000 16.280000 64.820000 ;
        RECT 16.080000 65.030000 16.280000 65.230000 ;
        RECT 16.080000 65.440000 16.280000 65.640000 ;
        RECT 16.080000 65.850000 16.280000 66.050000 ;
        RECT 16.080000 66.260000 16.280000 66.460000 ;
        RECT 16.485000 62.160000 16.685000 62.360000 ;
        RECT 16.485000 62.570000 16.685000 62.770000 ;
        RECT 16.485000 62.980000 16.685000 63.180000 ;
        RECT 16.485000 63.390000 16.685000 63.590000 ;
        RECT 16.485000 63.800000 16.685000 64.000000 ;
        RECT 16.485000 64.210000 16.685000 64.410000 ;
        RECT 16.485000 64.620000 16.685000 64.820000 ;
        RECT 16.485000 65.030000 16.685000 65.230000 ;
        RECT 16.485000 65.440000 16.685000 65.640000 ;
        RECT 16.485000 65.850000 16.685000 66.050000 ;
        RECT 16.485000 66.260000 16.685000 66.460000 ;
        RECT 16.890000 62.160000 17.090000 62.360000 ;
        RECT 16.890000 62.570000 17.090000 62.770000 ;
        RECT 16.890000 62.980000 17.090000 63.180000 ;
        RECT 16.890000 63.390000 17.090000 63.590000 ;
        RECT 16.890000 63.800000 17.090000 64.000000 ;
        RECT 16.890000 64.210000 17.090000 64.410000 ;
        RECT 16.890000 64.620000 17.090000 64.820000 ;
        RECT 16.890000 65.030000 17.090000 65.230000 ;
        RECT 16.890000 65.440000 17.090000 65.640000 ;
        RECT 16.890000 65.850000 17.090000 66.050000 ;
        RECT 16.890000 66.260000 17.090000 66.460000 ;
        RECT 17.295000 62.160000 17.495000 62.360000 ;
        RECT 17.295000 62.570000 17.495000 62.770000 ;
        RECT 17.295000 62.980000 17.495000 63.180000 ;
        RECT 17.295000 63.390000 17.495000 63.590000 ;
        RECT 17.295000 63.800000 17.495000 64.000000 ;
        RECT 17.295000 64.210000 17.495000 64.410000 ;
        RECT 17.295000 64.620000 17.495000 64.820000 ;
        RECT 17.295000 65.030000 17.495000 65.230000 ;
        RECT 17.295000 65.440000 17.495000 65.640000 ;
        RECT 17.295000 65.850000 17.495000 66.050000 ;
        RECT 17.295000 66.260000 17.495000 66.460000 ;
        RECT 17.700000 62.160000 17.900000 62.360000 ;
        RECT 17.700000 62.570000 17.900000 62.770000 ;
        RECT 17.700000 62.980000 17.900000 63.180000 ;
        RECT 17.700000 63.390000 17.900000 63.590000 ;
        RECT 17.700000 63.800000 17.900000 64.000000 ;
        RECT 17.700000 64.210000 17.900000 64.410000 ;
        RECT 17.700000 64.620000 17.900000 64.820000 ;
        RECT 17.700000 65.030000 17.900000 65.230000 ;
        RECT 17.700000 65.440000 17.900000 65.640000 ;
        RECT 17.700000 65.850000 17.900000 66.050000 ;
        RECT 17.700000 66.260000 17.900000 66.460000 ;
        RECT 18.105000 62.160000 18.305000 62.360000 ;
        RECT 18.105000 62.570000 18.305000 62.770000 ;
        RECT 18.105000 62.980000 18.305000 63.180000 ;
        RECT 18.105000 63.390000 18.305000 63.590000 ;
        RECT 18.105000 63.800000 18.305000 64.000000 ;
        RECT 18.105000 64.210000 18.305000 64.410000 ;
        RECT 18.105000 64.620000 18.305000 64.820000 ;
        RECT 18.105000 65.030000 18.305000 65.230000 ;
        RECT 18.105000 65.440000 18.305000 65.640000 ;
        RECT 18.105000 65.850000 18.305000 66.050000 ;
        RECT 18.105000 66.260000 18.305000 66.460000 ;
        RECT 18.510000 62.160000 18.710000 62.360000 ;
        RECT 18.510000 62.570000 18.710000 62.770000 ;
        RECT 18.510000 62.980000 18.710000 63.180000 ;
        RECT 18.510000 63.390000 18.710000 63.590000 ;
        RECT 18.510000 63.800000 18.710000 64.000000 ;
        RECT 18.510000 64.210000 18.710000 64.410000 ;
        RECT 18.510000 64.620000 18.710000 64.820000 ;
        RECT 18.510000 65.030000 18.710000 65.230000 ;
        RECT 18.510000 65.440000 18.710000 65.640000 ;
        RECT 18.510000 65.850000 18.710000 66.050000 ;
        RECT 18.510000 66.260000 18.710000 66.460000 ;
        RECT 18.915000 62.160000 19.115000 62.360000 ;
        RECT 18.915000 62.570000 19.115000 62.770000 ;
        RECT 18.915000 62.980000 19.115000 63.180000 ;
        RECT 18.915000 63.390000 19.115000 63.590000 ;
        RECT 18.915000 63.800000 19.115000 64.000000 ;
        RECT 18.915000 64.210000 19.115000 64.410000 ;
        RECT 18.915000 64.620000 19.115000 64.820000 ;
        RECT 18.915000 65.030000 19.115000 65.230000 ;
        RECT 18.915000 65.440000 19.115000 65.640000 ;
        RECT 18.915000 65.850000 19.115000 66.050000 ;
        RECT 18.915000 66.260000 19.115000 66.460000 ;
        RECT 19.320000 62.160000 19.520000 62.360000 ;
        RECT 19.320000 62.570000 19.520000 62.770000 ;
        RECT 19.320000 62.980000 19.520000 63.180000 ;
        RECT 19.320000 63.390000 19.520000 63.590000 ;
        RECT 19.320000 63.800000 19.520000 64.000000 ;
        RECT 19.320000 64.210000 19.520000 64.410000 ;
        RECT 19.320000 64.620000 19.520000 64.820000 ;
        RECT 19.320000 65.030000 19.520000 65.230000 ;
        RECT 19.320000 65.440000 19.520000 65.640000 ;
        RECT 19.320000 65.850000 19.520000 66.050000 ;
        RECT 19.320000 66.260000 19.520000 66.460000 ;
        RECT 19.725000 62.160000 19.925000 62.360000 ;
        RECT 19.725000 62.570000 19.925000 62.770000 ;
        RECT 19.725000 62.980000 19.925000 63.180000 ;
        RECT 19.725000 63.390000 19.925000 63.590000 ;
        RECT 19.725000 63.800000 19.925000 64.000000 ;
        RECT 19.725000 64.210000 19.925000 64.410000 ;
        RECT 19.725000 64.620000 19.925000 64.820000 ;
        RECT 19.725000 65.030000 19.925000 65.230000 ;
        RECT 19.725000 65.440000 19.925000 65.640000 ;
        RECT 19.725000 65.850000 19.925000 66.050000 ;
        RECT 19.725000 66.260000 19.925000 66.460000 ;
        RECT 20.130000 62.160000 20.330000 62.360000 ;
        RECT 20.130000 62.570000 20.330000 62.770000 ;
        RECT 20.130000 62.980000 20.330000 63.180000 ;
        RECT 20.130000 63.390000 20.330000 63.590000 ;
        RECT 20.130000 63.800000 20.330000 64.000000 ;
        RECT 20.130000 64.210000 20.330000 64.410000 ;
        RECT 20.130000 64.620000 20.330000 64.820000 ;
        RECT 20.130000 65.030000 20.330000 65.230000 ;
        RECT 20.130000 65.440000 20.330000 65.640000 ;
        RECT 20.130000 65.850000 20.330000 66.050000 ;
        RECT 20.130000 66.260000 20.330000 66.460000 ;
        RECT 20.535000 62.160000 20.735000 62.360000 ;
        RECT 20.535000 62.570000 20.735000 62.770000 ;
        RECT 20.535000 62.980000 20.735000 63.180000 ;
        RECT 20.535000 63.390000 20.735000 63.590000 ;
        RECT 20.535000 63.800000 20.735000 64.000000 ;
        RECT 20.535000 64.210000 20.735000 64.410000 ;
        RECT 20.535000 64.620000 20.735000 64.820000 ;
        RECT 20.535000 65.030000 20.735000 65.230000 ;
        RECT 20.535000 65.440000 20.735000 65.640000 ;
        RECT 20.535000 65.850000 20.735000 66.050000 ;
        RECT 20.535000 66.260000 20.735000 66.460000 ;
        RECT 20.940000 62.160000 21.140000 62.360000 ;
        RECT 20.940000 62.570000 21.140000 62.770000 ;
        RECT 20.940000 62.980000 21.140000 63.180000 ;
        RECT 20.940000 63.390000 21.140000 63.590000 ;
        RECT 20.940000 63.800000 21.140000 64.000000 ;
        RECT 20.940000 64.210000 21.140000 64.410000 ;
        RECT 20.940000 64.620000 21.140000 64.820000 ;
        RECT 20.940000 65.030000 21.140000 65.230000 ;
        RECT 20.940000 65.440000 21.140000 65.640000 ;
        RECT 20.940000 65.850000 21.140000 66.050000 ;
        RECT 20.940000 66.260000 21.140000 66.460000 ;
        RECT 21.345000 62.160000 21.545000 62.360000 ;
        RECT 21.345000 62.570000 21.545000 62.770000 ;
        RECT 21.345000 62.980000 21.545000 63.180000 ;
        RECT 21.345000 63.390000 21.545000 63.590000 ;
        RECT 21.345000 63.800000 21.545000 64.000000 ;
        RECT 21.345000 64.210000 21.545000 64.410000 ;
        RECT 21.345000 64.620000 21.545000 64.820000 ;
        RECT 21.345000 65.030000 21.545000 65.230000 ;
        RECT 21.345000 65.440000 21.545000 65.640000 ;
        RECT 21.345000 65.850000 21.545000 66.050000 ;
        RECT 21.345000 66.260000 21.545000 66.460000 ;
        RECT 21.750000 62.160000 21.950000 62.360000 ;
        RECT 21.750000 62.570000 21.950000 62.770000 ;
        RECT 21.750000 62.980000 21.950000 63.180000 ;
        RECT 21.750000 63.390000 21.950000 63.590000 ;
        RECT 21.750000 63.800000 21.950000 64.000000 ;
        RECT 21.750000 64.210000 21.950000 64.410000 ;
        RECT 21.750000 64.620000 21.950000 64.820000 ;
        RECT 21.750000 65.030000 21.950000 65.230000 ;
        RECT 21.750000 65.440000 21.950000 65.640000 ;
        RECT 21.750000 65.850000 21.950000 66.050000 ;
        RECT 21.750000 66.260000 21.950000 66.460000 ;
        RECT 22.160000 62.160000 22.360000 62.360000 ;
        RECT 22.160000 62.570000 22.360000 62.770000 ;
        RECT 22.160000 62.980000 22.360000 63.180000 ;
        RECT 22.160000 63.390000 22.360000 63.590000 ;
        RECT 22.160000 63.800000 22.360000 64.000000 ;
        RECT 22.160000 64.210000 22.360000 64.410000 ;
        RECT 22.160000 64.620000 22.360000 64.820000 ;
        RECT 22.160000 65.030000 22.360000 65.230000 ;
        RECT 22.160000 65.440000 22.360000 65.640000 ;
        RECT 22.160000 65.850000 22.360000 66.050000 ;
        RECT 22.160000 66.260000 22.360000 66.460000 ;
        RECT 22.570000 62.160000 22.770000 62.360000 ;
        RECT 22.570000 62.570000 22.770000 62.770000 ;
        RECT 22.570000 62.980000 22.770000 63.180000 ;
        RECT 22.570000 63.390000 22.770000 63.590000 ;
        RECT 22.570000 63.800000 22.770000 64.000000 ;
        RECT 22.570000 64.210000 22.770000 64.410000 ;
        RECT 22.570000 64.620000 22.770000 64.820000 ;
        RECT 22.570000 65.030000 22.770000 65.230000 ;
        RECT 22.570000 65.440000 22.770000 65.640000 ;
        RECT 22.570000 65.850000 22.770000 66.050000 ;
        RECT 22.570000 66.260000 22.770000 66.460000 ;
        RECT 22.980000 62.160000 23.180000 62.360000 ;
        RECT 22.980000 62.570000 23.180000 62.770000 ;
        RECT 22.980000 62.980000 23.180000 63.180000 ;
        RECT 22.980000 63.390000 23.180000 63.590000 ;
        RECT 22.980000 63.800000 23.180000 64.000000 ;
        RECT 22.980000 64.210000 23.180000 64.410000 ;
        RECT 22.980000 64.620000 23.180000 64.820000 ;
        RECT 22.980000 65.030000 23.180000 65.230000 ;
        RECT 22.980000 65.440000 23.180000 65.640000 ;
        RECT 22.980000 65.850000 23.180000 66.050000 ;
        RECT 22.980000 66.260000 23.180000 66.460000 ;
        RECT 23.390000 62.160000 23.590000 62.360000 ;
        RECT 23.390000 62.570000 23.590000 62.770000 ;
        RECT 23.390000 62.980000 23.590000 63.180000 ;
        RECT 23.390000 63.390000 23.590000 63.590000 ;
        RECT 23.390000 63.800000 23.590000 64.000000 ;
        RECT 23.390000 64.210000 23.590000 64.410000 ;
        RECT 23.390000 64.620000 23.590000 64.820000 ;
        RECT 23.390000 65.030000 23.590000 65.230000 ;
        RECT 23.390000 65.440000 23.590000 65.640000 ;
        RECT 23.390000 65.850000 23.590000 66.050000 ;
        RECT 23.390000 66.260000 23.590000 66.460000 ;
        RECT 23.800000 62.160000 24.000000 62.360000 ;
        RECT 23.800000 62.570000 24.000000 62.770000 ;
        RECT 23.800000 62.980000 24.000000 63.180000 ;
        RECT 23.800000 63.390000 24.000000 63.590000 ;
        RECT 23.800000 63.800000 24.000000 64.000000 ;
        RECT 23.800000 64.210000 24.000000 64.410000 ;
        RECT 23.800000 64.620000 24.000000 64.820000 ;
        RECT 23.800000 65.030000 24.000000 65.230000 ;
        RECT 23.800000 65.440000 24.000000 65.640000 ;
        RECT 23.800000 65.850000 24.000000 66.050000 ;
        RECT 23.800000 66.260000 24.000000 66.460000 ;
        RECT 24.210000 62.160000 24.410000 62.360000 ;
        RECT 24.210000 62.570000 24.410000 62.770000 ;
        RECT 24.210000 62.980000 24.410000 63.180000 ;
        RECT 24.210000 63.390000 24.410000 63.590000 ;
        RECT 24.210000 63.800000 24.410000 64.000000 ;
        RECT 24.210000 64.210000 24.410000 64.410000 ;
        RECT 24.210000 64.620000 24.410000 64.820000 ;
        RECT 24.210000 65.030000 24.410000 65.230000 ;
        RECT 24.210000 65.440000 24.410000 65.640000 ;
        RECT 24.210000 65.850000 24.410000 66.050000 ;
        RECT 24.210000 66.260000 24.410000 66.460000 ;
        RECT 50.845000 62.160000 51.045000 62.360000 ;
        RECT 50.845000 62.570000 51.045000 62.770000 ;
        RECT 50.845000 62.980000 51.045000 63.180000 ;
        RECT 50.845000 63.390000 51.045000 63.590000 ;
        RECT 50.845000 63.800000 51.045000 64.000000 ;
        RECT 50.845000 64.210000 51.045000 64.410000 ;
        RECT 50.845000 64.620000 51.045000 64.820000 ;
        RECT 50.845000 65.030000 51.045000 65.230000 ;
        RECT 50.845000 65.440000 51.045000 65.640000 ;
        RECT 50.845000 65.850000 51.045000 66.050000 ;
        RECT 50.845000 66.260000 51.045000 66.460000 ;
        RECT 51.250000 62.160000 51.450000 62.360000 ;
        RECT 51.250000 62.570000 51.450000 62.770000 ;
        RECT 51.250000 62.980000 51.450000 63.180000 ;
        RECT 51.250000 63.390000 51.450000 63.590000 ;
        RECT 51.250000 63.800000 51.450000 64.000000 ;
        RECT 51.250000 64.210000 51.450000 64.410000 ;
        RECT 51.250000 64.620000 51.450000 64.820000 ;
        RECT 51.250000 65.030000 51.450000 65.230000 ;
        RECT 51.250000 65.440000 51.450000 65.640000 ;
        RECT 51.250000 65.850000 51.450000 66.050000 ;
        RECT 51.250000 66.260000 51.450000 66.460000 ;
        RECT 51.655000 62.160000 51.855000 62.360000 ;
        RECT 51.655000 62.570000 51.855000 62.770000 ;
        RECT 51.655000 62.980000 51.855000 63.180000 ;
        RECT 51.655000 63.390000 51.855000 63.590000 ;
        RECT 51.655000 63.800000 51.855000 64.000000 ;
        RECT 51.655000 64.210000 51.855000 64.410000 ;
        RECT 51.655000 64.620000 51.855000 64.820000 ;
        RECT 51.655000 65.030000 51.855000 65.230000 ;
        RECT 51.655000 65.440000 51.855000 65.640000 ;
        RECT 51.655000 65.850000 51.855000 66.050000 ;
        RECT 51.655000 66.260000 51.855000 66.460000 ;
        RECT 52.060000 62.160000 52.260000 62.360000 ;
        RECT 52.060000 62.570000 52.260000 62.770000 ;
        RECT 52.060000 62.980000 52.260000 63.180000 ;
        RECT 52.060000 63.390000 52.260000 63.590000 ;
        RECT 52.060000 63.800000 52.260000 64.000000 ;
        RECT 52.060000 64.210000 52.260000 64.410000 ;
        RECT 52.060000 64.620000 52.260000 64.820000 ;
        RECT 52.060000 65.030000 52.260000 65.230000 ;
        RECT 52.060000 65.440000 52.260000 65.640000 ;
        RECT 52.060000 65.850000 52.260000 66.050000 ;
        RECT 52.060000 66.260000 52.260000 66.460000 ;
        RECT 52.465000 62.160000 52.665000 62.360000 ;
        RECT 52.465000 62.570000 52.665000 62.770000 ;
        RECT 52.465000 62.980000 52.665000 63.180000 ;
        RECT 52.465000 63.390000 52.665000 63.590000 ;
        RECT 52.465000 63.800000 52.665000 64.000000 ;
        RECT 52.465000 64.210000 52.665000 64.410000 ;
        RECT 52.465000 64.620000 52.665000 64.820000 ;
        RECT 52.465000 65.030000 52.665000 65.230000 ;
        RECT 52.465000 65.440000 52.665000 65.640000 ;
        RECT 52.465000 65.850000 52.665000 66.050000 ;
        RECT 52.465000 66.260000 52.665000 66.460000 ;
        RECT 52.870000 62.160000 53.070000 62.360000 ;
        RECT 52.870000 62.570000 53.070000 62.770000 ;
        RECT 52.870000 62.980000 53.070000 63.180000 ;
        RECT 52.870000 63.390000 53.070000 63.590000 ;
        RECT 52.870000 63.800000 53.070000 64.000000 ;
        RECT 52.870000 64.210000 53.070000 64.410000 ;
        RECT 52.870000 64.620000 53.070000 64.820000 ;
        RECT 52.870000 65.030000 53.070000 65.230000 ;
        RECT 52.870000 65.440000 53.070000 65.640000 ;
        RECT 52.870000 65.850000 53.070000 66.050000 ;
        RECT 52.870000 66.260000 53.070000 66.460000 ;
        RECT 53.275000 62.160000 53.475000 62.360000 ;
        RECT 53.275000 62.570000 53.475000 62.770000 ;
        RECT 53.275000 62.980000 53.475000 63.180000 ;
        RECT 53.275000 63.390000 53.475000 63.590000 ;
        RECT 53.275000 63.800000 53.475000 64.000000 ;
        RECT 53.275000 64.210000 53.475000 64.410000 ;
        RECT 53.275000 64.620000 53.475000 64.820000 ;
        RECT 53.275000 65.030000 53.475000 65.230000 ;
        RECT 53.275000 65.440000 53.475000 65.640000 ;
        RECT 53.275000 65.850000 53.475000 66.050000 ;
        RECT 53.275000 66.260000 53.475000 66.460000 ;
        RECT 53.680000 62.160000 53.880000 62.360000 ;
        RECT 53.680000 62.570000 53.880000 62.770000 ;
        RECT 53.680000 62.980000 53.880000 63.180000 ;
        RECT 53.680000 63.390000 53.880000 63.590000 ;
        RECT 53.680000 63.800000 53.880000 64.000000 ;
        RECT 53.680000 64.210000 53.880000 64.410000 ;
        RECT 53.680000 64.620000 53.880000 64.820000 ;
        RECT 53.680000 65.030000 53.880000 65.230000 ;
        RECT 53.680000 65.440000 53.880000 65.640000 ;
        RECT 53.680000 65.850000 53.880000 66.050000 ;
        RECT 53.680000 66.260000 53.880000 66.460000 ;
        RECT 54.085000 62.160000 54.285000 62.360000 ;
        RECT 54.085000 62.570000 54.285000 62.770000 ;
        RECT 54.085000 62.980000 54.285000 63.180000 ;
        RECT 54.085000 63.390000 54.285000 63.590000 ;
        RECT 54.085000 63.800000 54.285000 64.000000 ;
        RECT 54.085000 64.210000 54.285000 64.410000 ;
        RECT 54.085000 64.620000 54.285000 64.820000 ;
        RECT 54.085000 65.030000 54.285000 65.230000 ;
        RECT 54.085000 65.440000 54.285000 65.640000 ;
        RECT 54.085000 65.850000 54.285000 66.050000 ;
        RECT 54.085000 66.260000 54.285000 66.460000 ;
        RECT 54.490000 62.160000 54.690000 62.360000 ;
        RECT 54.490000 62.570000 54.690000 62.770000 ;
        RECT 54.490000 62.980000 54.690000 63.180000 ;
        RECT 54.490000 63.390000 54.690000 63.590000 ;
        RECT 54.490000 63.800000 54.690000 64.000000 ;
        RECT 54.490000 64.210000 54.690000 64.410000 ;
        RECT 54.490000 64.620000 54.690000 64.820000 ;
        RECT 54.490000 65.030000 54.690000 65.230000 ;
        RECT 54.490000 65.440000 54.690000 65.640000 ;
        RECT 54.490000 65.850000 54.690000 66.050000 ;
        RECT 54.490000 66.260000 54.690000 66.460000 ;
        RECT 54.895000 62.160000 55.095000 62.360000 ;
        RECT 54.895000 62.570000 55.095000 62.770000 ;
        RECT 54.895000 62.980000 55.095000 63.180000 ;
        RECT 54.895000 63.390000 55.095000 63.590000 ;
        RECT 54.895000 63.800000 55.095000 64.000000 ;
        RECT 54.895000 64.210000 55.095000 64.410000 ;
        RECT 54.895000 64.620000 55.095000 64.820000 ;
        RECT 54.895000 65.030000 55.095000 65.230000 ;
        RECT 54.895000 65.440000 55.095000 65.640000 ;
        RECT 54.895000 65.850000 55.095000 66.050000 ;
        RECT 54.895000 66.260000 55.095000 66.460000 ;
        RECT 55.300000 62.160000 55.500000 62.360000 ;
        RECT 55.300000 62.570000 55.500000 62.770000 ;
        RECT 55.300000 62.980000 55.500000 63.180000 ;
        RECT 55.300000 63.390000 55.500000 63.590000 ;
        RECT 55.300000 63.800000 55.500000 64.000000 ;
        RECT 55.300000 64.210000 55.500000 64.410000 ;
        RECT 55.300000 64.620000 55.500000 64.820000 ;
        RECT 55.300000 65.030000 55.500000 65.230000 ;
        RECT 55.300000 65.440000 55.500000 65.640000 ;
        RECT 55.300000 65.850000 55.500000 66.050000 ;
        RECT 55.300000 66.260000 55.500000 66.460000 ;
        RECT 55.705000 62.160000 55.905000 62.360000 ;
        RECT 55.705000 62.570000 55.905000 62.770000 ;
        RECT 55.705000 62.980000 55.905000 63.180000 ;
        RECT 55.705000 63.390000 55.905000 63.590000 ;
        RECT 55.705000 63.800000 55.905000 64.000000 ;
        RECT 55.705000 64.210000 55.905000 64.410000 ;
        RECT 55.705000 64.620000 55.905000 64.820000 ;
        RECT 55.705000 65.030000 55.905000 65.230000 ;
        RECT 55.705000 65.440000 55.905000 65.640000 ;
        RECT 55.705000 65.850000 55.905000 66.050000 ;
        RECT 55.705000 66.260000 55.905000 66.460000 ;
        RECT 56.110000 62.160000 56.310000 62.360000 ;
        RECT 56.110000 62.570000 56.310000 62.770000 ;
        RECT 56.110000 62.980000 56.310000 63.180000 ;
        RECT 56.110000 63.390000 56.310000 63.590000 ;
        RECT 56.110000 63.800000 56.310000 64.000000 ;
        RECT 56.110000 64.210000 56.310000 64.410000 ;
        RECT 56.110000 64.620000 56.310000 64.820000 ;
        RECT 56.110000 65.030000 56.310000 65.230000 ;
        RECT 56.110000 65.440000 56.310000 65.640000 ;
        RECT 56.110000 65.850000 56.310000 66.050000 ;
        RECT 56.110000 66.260000 56.310000 66.460000 ;
        RECT 56.515000 62.160000 56.715000 62.360000 ;
        RECT 56.515000 62.570000 56.715000 62.770000 ;
        RECT 56.515000 62.980000 56.715000 63.180000 ;
        RECT 56.515000 63.390000 56.715000 63.590000 ;
        RECT 56.515000 63.800000 56.715000 64.000000 ;
        RECT 56.515000 64.210000 56.715000 64.410000 ;
        RECT 56.515000 64.620000 56.715000 64.820000 ;
        RECT 56.515000 65.030000 56.715000 65.230000 ;
        RECT 56.515000 65.440000 56.715000 65.640000 ;
        RECT 56.515000 65.850000 56.715000 66.050000 ;
        RECT 56.515000 66.260000 56.715000 66.460000 ;
        RECT 56.920000 62.160000 57.120000 62.360000 ;
        RECT 56.920000 62.570000 57.120000 62.770000 ;
        RECT 56.920000 62.980000 57.120000 63.180000 ;
        RECT 56.920000 63.390000 57.120000 63.590000 ;
        RECT 56.920000 63.800000 57.120000 64.000000 ;
        RECT 56.920000 64.210000 57.120000 64.410000 ;
        RECT 56.920000 64.620000 57.120000 64.820000 ;
        RECT 56.920000 65.030000 57.120000 65.230000 ;
        RECT 56.920000 65.440000 57.120000 65.640000 ;
        RECT 56.920000 65.850000 57.120000 66.050000 ;
        RECT 56.920000 66.260000 57.120000 66.460000 ;
        RECT 57.325000 62.160000 57.525000 62.360000 ;
        RECT 57.325000 62.570000 57.525000 62.770000 ;
        RECT 57.325000 62.980000 57.525000 63.180000 ;
        RECT 57.325000 63.390000 57.525000 63.590000 ;
        RECT 57.325000 63.800000 57.525000 64.000000 ;
        RECT 57.325000 64.210000 57.525000 64.410000 ;
        RECT 57.325000 64.620000 57.525000 64.820000 ;
        RECT 57.325000 65.030000 57.525000 65.230000 ;
        RECT 57.325000 65.440000 57.525000 65.640000 ;
        RECT 57.325000 65.850000 57.525000 66.050000 ;
        RECT 57.325000 66.260000 57.525000 66.460000 ;
        RECT 57.730000 62.160000 57.930000 62.360000 ;
        RECT 57.730000 62.570000 57.930000 62.770000 ;
        RECT 57.730000 62.980000 57.930000 63.180000 ;
        RECT 57.730000 63.390000 57.930000 63.590000 ;
        RECT 57.730000 63.800000 57.930000 64.000000 ;
        RECT 57.730000 64.210000 57.930000 64.410000 ;
        RECT 57.730000 64.620000 57.930000 64.820000 ;
        RECT 57.730000 65.030000 57.930000 65.230000 ;
        RECT 57.730000 65.440000 57.930000 65.640000 ;
        RECT 57.730000 65.850000 57.930000 66.050000 ;
        RECT 57.730000 66.260000 57.930000 66.460000 ;
        RECT 58.135000 62.160000 58.335000 62.360000 ;
        RECT 58.135000 62.570000 58.335000 62.770000 ;
        RECT 58.135000 62.980000 58.335000 63.180000 ;
        RECT 58.135000 63.390000 58.335000 63.590000 ;
        RECT 58.135000 63.800000 58.335000 64.000000 ;
        RECT 58.135000 64.210000 58.335000 64.410000 ;
        RECT 58.135000 64.620000 58.335000 64.820000 ;
        RECT 58.135000 65.030000 58.335000 65.230000 ;
        RECT 58.135000 65.440000 58.335000 65.640000 ;
        RECT 58.135000 65.850000 58.335000 66.050000 ;
        RECT 58.135000 66.260000 58.335000 66.460000 ;
        RECT 58.540000 62.160000 58.740000 62.360000 ;
        RECT 58.540000 62.570000 58.740000 62.770000 ;
        RECT 58.540000 62.980000 58.740000 63.180000 ;
        RECT 58.540000 63.390000 58.740000 63.590000 ;
        RECT 58.540000 63.800000 58.740000 64.000000 ;
        RECT 58.540000 64.210000 58.740000 64.410000 ;
        RECT 58.540000 64.620000 58.740000 64.820000 ;
        RECT 58.540000 65.030000 58.740000 65.230000 ;
        RECT 58.540000 65.440000 58.740000 65.640000 ;
        RECT 58.540000 65.850000 58.740000 66.050000 ;
        RECT 58.540000 66.260000 58.740000 66.460000 ;
        RECT 58.945000 62.160000 59.145000 62.360000 ;
        RECT 58.945000 62.570000 59.145000 62.770000 ;
        RECT 58.945000 62.980000 59.145000 63.180000 ;
        RECT 58.945000 63.390000 59.145000 63.590000 ;
        RECT 58.945000 63.800000 59.145000 64.000000 ;
        RECT 58.945000 64.210000 59.145000 64.410000 ;
        RECT 58.945000 64.620000 59.145000 64.820000 ;
        RECT 58.945000 65.030000 59.145000 65.230000 ;
        RECT 58.945000 65.440000 59.145000 65.640000 ;
        RECT 58.945000 65.850000 59.145000 66.050000 ;
        RECT 58.945000 66.260000 59.145000 66.460000 ;
        RECT 59.350000 62.160000 59.550000 62.360000 ;
        RECT 59.350000 62.570000 59.550000 62.770000 ;
        RECT 59.350000 62.980000 59.550000 63.180000 ;
        RECT 59.350000 63.390000 59.550000 63.590000 ;
        RECT 59.350000 63.800000 59.550000 64.000000 ;
        RECT 59.350000 64.210000 59.550000 64.410000 ;
        RECT 59.350000 64.620000 59.550000 64.820000 ;
        RECT 59.350000 65.030000 59.550000 65.230000 ;
        RECT 59.350000 65.440000 59.550000 65.640000 ;
        RECT 59.350000 65.850000 59.550000 66.050000 ;
        RECT 59.350000 66.260000 59.550000 66.460000 ;
        RECT 59.755000 62.160000 59.955000 62.360000 ;
        RECT 59.755000 62.570000 59.955000 62.770000 ;
        RECT 59.755000 62.980000 59.955000 63.180000 ;
        RECT 59.755000 63.390000 59.955000 63.590000 ;
        RECT 59.755000 63.800000 59.955000 64.000000 ;
        RECT 59.755000 64.210000 59.955000 64.410000 ;
        RECT 59.755000 64.620000 59.955000 64.820000 ;
        RECT 59.755000 65.030000 59.955000 65.230000 ;
        RECT 59.755000 65.440000 59.955000 65.640000 ;
        RECT 59.755000 65.850000 59.955000 66.050000 ;
        RECT 59.755000 66.260000 59.955000 66.460000 ;
        RECT 60.160000 62.160000 60.360000 62.360000 ;
        RECT 60.160000 62.570000 60.360000 62.770000 ;
        RECT 60.160000 62.980000 60.360000 63.180000 ;
        RECT 60.160000 63.390000 60.360000 63.590000 ;
        RECT 60.160000 63.800000 60.360000 64.000000 ;
        RECT 60.160000 64.210000 60.360000 64.410000 ;
        RECT 60.160000 64.620000 60.360000 64.820000 ;
        RECT 60.160000 65.030000 60.360000 65.230000 ;
        RECT 60.160000 65.440000 60.360000 65.640000 ;
        RECT 60.160000 65.850000 60.360000 66.050000 ;
        RECT 60.160000 66.260000 60.360000 66.460000 ;
        RECT 60.565000 62.160000 60.765000 62.360000 ;
        RECT 60.565000 62.570000 60.765000 62.770000 ;
        RECT 60.565000 62.980000 60.765000 63.180000 ;
        RECT 60.565000 63.390000 60.765000 63.590000 ;
        RECT 60.565000 63.800000 60.765000 64.000000 ;
        RECT 60.565000 64.210000 60.765000 64.410000 ;
        RECT 60.565000 64.620000 60.765000 64.820000 ;
        RECT 60.565000 65.030000 60.765000 65.230000 ;
        RECT 60.565000 65.440000 60.765000 65.640000 ;
        RECT 60.565000 65.850000 60.765000 66.050000 ;
        RECT 60.565000 66.260000 60.765000 66.460000 ;
        RECT 60.970000 62.160000 61.170000 62.360000 ;
        RECT 60.970000 62.570000 61.170000 62.770000 ;
        RECT 60.970000 62.980000 61.170000 63.180000 ;
        RECT 60.970000 63.390000 61.170000 63.590000 ;
        RECT 60.970000 63.800000 61.170000 64.000000 ;
        RECT 60.970000 64.210000 61.170000 64.410000 ;
        RECT 60.970000 64.620000 61.170000 64.820000 ;
        RECT 60.970000 65.030000 61.170000 65.230000 ;
        RECT 60.970000 65.440000 61.170000 65.640000 ;
        RECT 60.970000 65.850000 61.170000 66.050000 ;
        RECT 60.970000 66.260000 61.170000 66.460000 ;
        RECT 61.375000 62.160000 61.575000 62.360000 ;
        RECT 61.375000 62.570000 61.575000 62.770000 ;
        RECT 61.375000 62.980000 61.575000 63.180000 ;
        RECT 61.375000 63.390000 61.575000 63.590000 ;
        RECT 61.375000 63.800000 61.575000 64.000000 ;
        RECT 61.375000 64.210000 61.575000 64.410000 ;
        RECT 61.375000 64.620000 61.575000 64.820000 ;
        RECT 61.375000 65.030000 61.575000 65.230000 ;
        RECT 61.375000 65.440000 61.575000 65.640000 ;
        RECT 61.375000 65.850000 61.575000 66.050000 ;
        RECT 61.375000 66.260000 61.575000 66.460000 ;
        RECT 61.780000 62.160000 61.980000 62.360000 ;
        RECT 61.780000 62.570000 61.980000 62.770000 ;
        RECT 61.780000 62.980000 61.980000 63.180000 ;
        RECT 61.780000 63.390000 61.980000 63.590000 ;
        RECT 61.780000 63.800000 61.980000 64.000000 ;
        RECT 61.780000 64.210000 61.980000 64.410000 ;
        RECT 61.780000 64.620000 61.980000 64.820000 ;
        RECT 61.780000 65.030000 61.980000 65.230000 ;
        RECT 61.780000 65.440000 61.980000 65.640000 ;
        RECT 61.780000 65.850000 61.980000 66.050000 ;
        RECT 61.780000 66.260000 61.980000 66.460000 ;
        RECT 62.185000 62.160000 62.385000 62.360000 ;
        RECT 62.185000 62.570000 62.385000 62.770000 ;
        RECT 62.185000 62.980000 62.385000 63.180000 ;
        RECT 62.185000 63.390000 62.385000 63.590000 ;
        RECT 62.185000 63.800000 62.385000 64.000000 ;
        RECT 62.185000 64.210000 62.385000 64.410000 ;
        RECT 62.185000 64.620000 62.385000 64.820000 ;
        RECT 62.185000 65.030000 62.385000 65.230000 ;
        RECT 62.185000 65.440000 62.385000 65.640000 ;
        RECT 62.185000 65.850000 62.385000 66.050000 ;
        RECT 62.185000 66.260000 62.385000 66.460000 ;
        RECT 62.590000 62.160000 62.790000 62.360000 ;
        RECT 62.590000 62.570000 62.790000 62.770000 ;
        RECT 62.590000 62.980000 62.790000 63.180000 ;
        RECT 62.590000 63.390000 62.790000 63.590000 ;
        RECT 62.590000 63.800000 62.790000 64.000000 ;
        RECT 62.590000 64.210000 62.790000 64.410000 ;
        RECT 62.590000 64.620000 62.790000 64.820000 ;
        RECT 62.590000 65.030000 62.790000 65.230000 ;
        RECT 62.590000 65.440000 62.790000 65.640000 ;
        RECT 62.590000 65.850000 62.790000 66.050000 ;
        RECT 62.590000 66.260000 62.790000 66.460000 ;
        RECT 62.995000 62.160000 63.195000 62.360000 ;
        RECT 62.995000 62.570000 63.195000 62.770000 ;
        RECT 62.995000 62.980000 63.195000 63.180000 ;
        RECT 62.995000 63.390000 63.195000 63.590000 ;
        RECT 62.995000 63.800000 63.195000 64.000000 ;
        RECT 62.995000 64.210000 63.195000 64.410000 ;
        RECT 62.995000 64.620000 63.195000 64.820000 ;
        RECT 62.995000 65.030000 63.195000 65.230000 ;
        RECT 62.995000 65.440000 63.195000 65.640000 ;
        RECT 62.995000 65.850000 63.195000 66.050000 ;
        RECT 62.995000 66.260000 63.195000 66.460000 ;
        RECT 63.400000 62.160000 63.600000 62.360000 ;
        RECT 63.400000 62.570000 63.600000 62.770000 ;
        RECT 63.400000 62.980000 63.600000 63.180000 ;
        RECT 63.400000 63.390000 63.600000 63.590000 ;
        RECT 63.400000 63.800000 63.600000 64.000000 ;
        RECT 63.400000 64.210000 63.600000 64.410000 ;
        RECT 63.400000 64.620000 63.600000 64.820000 ;
        RECT 63.400000 65.030000 63.600000 65.230000 ;
        RECT 63.400000 65.440000 63.600000 65.640000 ;
        RECT 63.400000 65.850000 63.600000 66.050000 ;
        RECT 63.400000 66.260000 63.600000 66.460000 ;
        RECT 63.805000 62.160000 64.005000 62.360000 ;
        RECT 63.805000 62.570000 64.005000 62.770000 ;
        RECT 63.805000 62.980000 64.005000 63.180000 ;
        RECT 63.805000 63.390000 64.005000 63.590000 ;
        RECT 63.805000 63.800000 64.005000 64.000000 ;
        RECT 63.805000 64.210000 64.005000 64.410000 ;
        RECT 63.805000 64.620000 64.005000 64.820000 ;
        RECT 63.805000 65.030000 64.005000 65.230000 ;
        RECT 63.805000 65.440000 64.005000 65.640000 ;
        RECT 63.805000 65.850000 64.005000 66.050000 ;
        RECT 63.805000 66.260000 64.005000 66.460000 ;
        RECT 64.210000 62.160000 64.410000 62.360000 ;
        RECT 64.210000 62.570000 64.410000 62.770000 ;
        RECT 64.210000 62.980000 64.410000 63.180000 ;
        RECT 64.210000 63.390000 64.410000 63.590000 ;
        RECT 64.210000 63.800000 64.410000 64.000000 ;
        RECT 64.210000 64.210000 64.410000 64.410000 ;
        RECT 64.210000 64.620000 64.410000 64.820000 ;
        RECT 64.210000 65.030000 64.410000 65.230000 ;
        RECT 64.210000 65.440000 64.410000 65.640000 ;
        RECT 64.210000 65.850000 64.410000 66.050000 ;
        RECT 64.210000 66.260000 64.410000 66.460000 ;
        RECT 64.615000 62.160000 64.815000 62.360000 ;
        RECT 64.615000 62.570000 64.815000 62.770000 ;
        RECT 64.615000 62.980000 64.815000 63.180000 ;
        RECT 64.615000 63.390000 64.815000 63.590000 ;
        RECT 64.615000 63.800000 64.815000 64.000000 ;
        RECT 64.615000 64.210000 64.815000 64.410000 ;
        RECT 64.615000 64.620000 64.815000 64.820000 ;
        RECT 64.615000 65.030000 64.815000 65.230000 ;
        RECT 64.615000 65.440000 64.815000 65.640000 ;
        RECT 64.615000 65.850000 64.815000 66.050000 ;
        RECT 64.615000 66.260000 64.815000 66.460000 ;
        RECT 65.020000 62.160000 65.220000 62.360000 ;
        RECT 65.020000 62.570000 65.220000 62.770000 ;
        RECT 65.020000 62.980000 65.220000 63.180000 ;
        RECT 65.020000 63.390000 65.220000 63.590000 ;
        RECT 65.020000 63.800000 65.220000 64.000000 ;
        RECT 65.020000 64.210000 65.220000 64.410000 ;
        RECT 65.020000 64.620000 65.220000 64.820000 ;
        RECT 65.020000 65.030000 65.220000 65.230000 ;
        RECT 65.020000 65.440000 65.220000 65.640000 ;
        RECT 65.020000 65.850000 65.220000 66.050000 ;
        RECT 65.020000 66.260000 65.220000 66.460000 ;
        RECT 65.425000 62.160000 65.625000 62.360000 ;
        RECT 65.425000 62.570000 65.625000 62.770000 ;
        RECT 65.425000 62.980000 65.625000 63.180000 ;
        RECT 65.425000 63.390000 65.625000 63.590000 ;
        RECT 65.425000 63.800000 65.625000 64.000000 ;
        RECT 65.425000 64.210000 65.625000 64.410000 ;
        RECT 65.425000 64.620000 65.625000 64.820000 ;
        RECT 65.425000 65.030000 65.625000 65.230000 ;
        RECT 65.425000 65.440000 65.625000 65.640000 ;
        RECT 65.425000 65.850000 65.625000 66.050000 ;
        RECT 65.425000 66.260000 65.625000 66.460000 ;
        RECT 65.830000 62.160000 66.030000 62.360000 ;
        RECT 65.830000 62.570000 66.030000 62.770000 ;
        RECT 65.830000 62.980000 66.030000 63.180000 ;
        RECT 65.830000 63.390000 66.030000 63.590000 ;
        RECT 65.830000 63.800000 66.030000 64.000000 ;
        RECT 65.830000 64.210000 66.030000 64.410000 ;
        RECT 65.830000 64.620000 66.030000 64.820000 ;
        RECT 65.830000 65.030000 66.030000 65.230000 ;
        RECT 65.830000 65.440000 66.030000 65.640000 ;
        RECT 65.830000 65.850000 66.030000 66.050000 ;
        RECT 65.830000 66.260000 66.030000 66.460000 ;
        RECT 66.235000 62.160000 66.435000 62.360000 ;
        RECT 66.235000 62.570000 66.435000 62.770000 ;
        RECT 66.235000 62.980000 66.435000 63.180000 ;
        RECT 66.235000 63.390000 66.435000 63.590000 ;
        RECT 66.235000 63.800000 66.435000 64.000000 ;
        RECT 66.235000 64.210000 66.435000 64.410000 ;
        RECT 66.235000 64.620000 66.435000 64.820000 ;
        RECT 66.235000 65.030000 66.435000 65.230000 ;
        RECT 66.235000 65.440000 66.435000 65.640000 ;
        RECT 66.235000 65.850000 66.435000 66.050000 ;
        RECT 66.235000 66.260000 66.435000 66.460000 ;
        RECT 66.640000 62.160000 66.840000 62.360000 ;
        RECT 66.640000 62.570000 66.840000 62.770000 ;
        RECT 66.640000 62.980000 66.840000 63.180000 ;
        RECT 66.640000 63.390000 66.840000 63.590000 ;
        RECT 66.640000 63.800000 66.840000 64.000000 ;
        RECT 66.640000 64.210000 66.840000 64.410000 ;
        RECT 66.640000 64.620000 66.840000 64.820000 ;
        RECT 66.640000 65.030000 66.840000 65.230000 ;
        RECT 66.640000 65.440000 66.840000 65.640000 ;
        RECT 66.640000 65.850000 66.840000 66.050000 ;
        RECT 66.640000 66.260000 66.840000 66.460000 ;
        RECT 67.045000 62.160000 67.245000 62.360000 ;
        RECT 67.045000 62.570000 67.245000 62.770000 ;
        RECT 67.045000 62.980000 67.245000 63.180000 ;
        RECT 67.045000 63.390000 67.245000 63.590000 ;
        RECT 67.045000 63.800000 67.245000 64.000000 ;
        RECT 67.045000 64.210000 67.245000 64.410000 ;
        RECT 67.045000 64.620000 67.245000 64.820000 ;
        RECT 67.045000 65.030000 67.245000 65.230000 ;
        RECT 67.045000 65.440000 67.245000 65.640000 ;
        RECT 67.045000 65.850000 67.245000 66.050000 ;
        RECT 67.045000 66.260000 67.245000 66.460000 ;
        RECT 67.450000 62.160000 67.650000 62.360000 ;
        RECT 67.450000 62.570000 67.650000 62.770000 ;
        RECT 67.450000 62.980000 67.650000 63.180000 ;
        RECT 67.450000 63.390000 67.650000 63.590000 ;
        RECT 67.450000 63.800000 67.650000 64.000000 ;
        RECT 67.450000 64.210000 67.650000 64.410000 ;
        RECT 67.450000 64.620000 67.650000 64.820000 ;
        RECT 67.450000 65.030000 67.650000 65.230000 ;
        RECT 67.450000 65.440000 67.650000 65.640000 ;
        RECT 67.450000 65.850000 67.650000 66.050000 ;
        RECT 67.450000 66.260000 67.650000 66.460000 ;
        RECT 67.855000 62.160000 68.055000 62.360000 ;
        RECT 67.855000 62.570000 68.055000 62.770000 ;
        RECT 67.855000 62.980000 68.055000 63.180000 ;
        RECT 67.855000 63.390000 68.055000 63.590000 ;
        RECT 67.855000 63.800000 68.055000 64.000000 ;
        RECT 67.855000 64.210000 68.055000 64.410000 ;
        RECT 67.855000 64.620000 68.055000 64.820000 ;
        RECT 67.855000 65.030000 68.055000 65.230000 ;
        RECT 67.855000 65.440000 68.055000 65.640000 ;
        RECT 67.855000 65.850000 68.055000 66.050000 ;
        RECT 67.855000 66.260000 68.055000 66.460000 ;
        RECT 68.260000 62.160000 68.460000 62.360000 ;
        RECT 68.260000 62.570000 68.460000 62.770000 ;
        RECT 68.260000 62.980000 68.460000 63.180000 ;
        RECT 68.260000 63.390000 68.460000 63.590000 ;
        RECT 68.260000 63.800000 68.460000 64.000000 ;
        RECT 68.260000 64.210000 68.460000 64.410000 ;
        RECT 68.260000 64.620000 68.460000 64.820000 ;
        RECT 68.260000 65.030000 68.460000 65.230000 ;
        RECT 68.260000 65.440000 68.460000 65.640000 ;
        RECT 68.260000 65.850000 68.460000 66.050000 ;
        RECT 68.260000 66.260000 68.460000 66.460000 ;
        RECT 68.665000 62.160000 68.865000 62.360000 ;
        RECT 68.665000 62.570000 68.865000 62.770000 ;
        RECT 68.665000 62.980000 68.865000 63.180000 ;
        RECT 68.665000 63.390000 68.865000 63.590000 ;
        RECT 68.665000 63.800000 68.865000 64.000000 ;
        RECT 68.665000 64.210000 68.865000 64.410000 ;
        RECT 68.665000 64.620000 68.865000 64.820000 ;
        RECT 68.665000 65.030000 68.865000 65.230000 ;
        RECT 68.665000 65.440000 68.865000 65.640000 ;
        RECT 68.665000 65.850000 68.865000 66.050000 ;
        RECT 68.665000 66.260000 68.865000 66.460000 ;
        RECT 69.070000 62.160000 69.270000 62.360000 ;
        RECT 69.070000 62.570000 69.270000 62.770000 ;
        RECT 69.070000 62.980000 69.270000 63.180000 ;
        RECT 69.070000 63.390000 69.270000 63.590000 ;
        RECT 69.070000 63.800000 69.270000 64.000000 ;
        RECT 69.070000 64.210000 69.270000 64.410000 ;
        RECT 69.070000 64.620000 69.270000 64.820000 ;
        RECT 69.070000 65.030000 69.270000 65.230000 ;
        RECT 69.070000 65.440000 69.270000 65.640000 ;
        RECT 69.070000 65.850000 69.270000 66.050000 ;
        RECT 69.070000 66.260000 69.270000 66.460000 ;
        RECT 69.475000 62.160000 69.675000 62.360000 ;
        RECT 69.475000 62.570000 69.675000 62.770000 ;
        RECT 69.475000 62.980000 69.675000 63.180000 ;
        RECT 69.475000 63.390000 69.675000 63.590000 ;
        RECT 69.475000 63.800000 69.675000 64.000000 ;
        RECT 69.475000 64.210000 69.675000 64.410000 ;
        RECT 69.475000 64.620000 69.675000 64.820000 ;
        RECT 69.475000 65.030000 69.675000 65.230000 ;
        RECT 69.475000 65.440000 69.675000 65.640000 ;
        RECT 69.475000 65.850000 69.675000 66.050000 ;
        RECT 69.475000 66.260000 69.675000 66.460000 ;
        RECT 69.880000 62.160000 70.080000 62.360000 ;
        RECT 69.880000 62.570000 70.080000 62.770000 ;
        RECT 69.880000 62.980000 70.080000 63.180000 ;
        RECT 69.880000 63.390000 70.080000 63.590000 ;
        RECT 69.880000 63.800000 70.080000 64.000000 ;
        RECT 69.880000 64.210000 70.080000 64.410000 ;
        RECT 69.880000 64.620000 70.080000 64.820000 ;
        RECT 69.880000 65.030000 70.080000 65.230000 ;
        RECT 69.880000 65.440000 70.080000 65.640000 ;
        RECT 69.880000 65.850000 70.080000 66.050000 ;
        RECT 69.880000 66.260000 70.080000 66.460000 ;
        RECT 70.285000 62.160000 70.485000 62.360000 ;
        RECT 70.285000 62.570000 70.485000 62.770000 ;
        RECT 70.285000 62.980000 70.485000 63.180000 ;
        RECT 70.285000 63.390000 70.485000 63.590000 ;
        RECT 70.285000 63.800000 70.485000 64.000000 ;
        RECT 70.285000 64.210000 70.485000 64.410000 ;
        RECT 70.285000 64.620000 70.485000 64.820000 ;
        RECT 70.285000 65.030000 70.485000 65.230000 ;
        RECT 70.285000 65.440000 70.485000 65.640000 ;
        RECT 70.285000 65.850000 70.485000 66.050000 ;
        RECT 70.285000 66.260000 70.485000 66.460000 ;
        RECT 70.690000 62.160000 70.890000 62.360000 ;
        RECT 70.690000 62.570000 70.890000 62.770000 ;
        RECT 70.690000 62.980000 70.890000 63.180000 ;
        RECT 70.690000 63.390000 70.890000 63.590000 ;
        RECT 70.690000 63.800000 70.890000 64.000000 ;
        RECT 70.690000 64.210000 70.890000 64.410000 ;
        RECT 70.690000 64.620000 70.890000 64.820000 ;
        RECT 70.690000 65.030000 70.890000 65.230000 ;
        RECT 70.690000 65.440000 70.890000 65.640000 ;
        RECT 70.690000 65.850000 70.890000 66.050000 ;
        RECT 70.690000 66.260000 70.890000 66.460000 ;
        RECT 71.095000 62.160000 71.295000 62.360000 ;
        RECT 71.095000 62.570000 71.295000 62.770000 ;
        RECT 71.095000 62.980000 71.295000 63.180000 ;
        RECT 71.095000 63.390000 71.295000 63.590000 ;
        RECT 71.095000 63.800000 71.295000 64.000000 ;
        RECT 71.095000 64.210000 71.295000 64.410000 ;
        RECT 71.095000 64.620000 71.295000 64.820000 ;
        RECT 71.095000 65.030000 71.295000 65.230000 ;
        RECT 71.095000 65.440000 71.295000 65.640000 ;
        RECT 71.095000 65.850000 71.295000 66.050000 ;
        RECT 71.095000 66.260000 71.295000 66.460000 ;
        RECT 71.500000 62.160000 71.700000 62.360000 ;
        RECT 71.500000 62.570000 71.700000 62.770000 ;
        RECT 71.500000 62.980000 71.700000 63.180000 ;
        RECT 71.500000 63.390000 71.700000 63.590000 ;
        RECT 71.500000 63.800000 71.700000 64.000000 ;
        RECT 71.500000 64.210000 71.700000 64.410000 ;
        RECT 71.500000 64.620000 71.700000 64.820000 ;
        RECT 71.500000 65.030000 71.700000 65.230000 ;
        RECT 71.500000 65.440000 71.700000 65.640000 ;
        RECT 71.500000 65.850000 71.700000 66.050000 ;
        RECT 71.500000 66.260000 71.700000 66.460000 ;
        RECT 71.905000 62.160000 72.105000 62.360000 ;
        RECT 71.905000 62.570000 72.105000 62.770000 ;
        RECT 71.905000 62.980000 72.105000 63.180000 ;
        RECT 71.905000 63.390000 72.105000 63.590000 ;
        RECT 71.905000 63.800000 72.105000 64.000000 ;
        RECT 71.905000 64.210000 72.105000 64.410000 ;
        RECT 71.905000 64.620000 72.105000 64.820000 ;
        RECT 71.905000 65.030000 72.105000 65.230000 ;
        RECT 71.905000 65.440000 72.105000 65.640000 ;
        RECT 71.905000 65.850000 72.105000 66.050000 ;
        RECT 71.905000 66.260000 72.105000 66.460000 ;
        RECT 72.315000 62.160000 72.515000 62.360000 ;
        RECT 72.315000 62.570000 72.515000 62.770000 ;
        RECT 72.315000 62.980000 72.515000 63.180000 ;
        RECT 72.315000 63.390000 72.515000 63.590000 ;
        RECT 72.315000 63.800000 72.515000 64.000000 ;
        RECT 72.315000 64.210000 72.515000 64.410000 ;
        RECT 72.315000 64.620000 72.515000 64.820000 ;
        RECT 72.315000 65.030000 72.515000 65.230000 ;
        RECT 72.315000 65.440000 72.515000 65.640000 ;
        RECT 72.315000 65.850000 72.515000 66.050000 ;
        RECT 72.315000 66.260000 72.515000 66.460000 ;
        RECT 72.725000 62.160000 72.925000 62.360000 ;
        RECT 72.725000 62.570000 72.925000 62.770000 ;
        RECT 72.725000 62.980000 72.925000 63.180000 ;
        RECT 72.725000 63.390000 72.925000 63.590000 ;
        RECT 72.725000 63.800000 72.925000 64.000000 ;
        RECT 72.725000 64.210000 72.925000 64.410000 ;
        RECT 72.725000 64.620000 72.925000 64.820000 ;
        RECT 72.725000 65.030000 72.925000 65.230000 ;
        RECT 72.725000 65.440000 72.925000 65.640000 ;
        RECT 72.725000 65.850000 72.925000 66.050000 ;
        RECT 72.725000 66.260000 72.925000 66.460000 ;
        RECT 73.135000 62.160000 73.335000 62.360000 ;
        RECT 73.135000 62.570000 73.335000 62.770000 ;
        RECT 73.135000 62.980000 73.335000 63.180000 ;
        RECT 73.135000 63.390000 73.335000 63.590000 ;
        RECT 73.135000 63.800000 73.335000 64.000000 ;
        RECT 73.135000 64.210000 73.335000 64.410000 ;
        RECT 73.135000 64.620000 73.335000 64.820000 ;
        RECT 73.135000 65.030000 73.335000 65.230000 ;
        RECT 73.135000 65.440000 73.335000 65.640000 ;
        RECT 73.135000 65.850000 73.335000 66.050000 ;
        RECT 73.135000 66.260000 73.335000 66.460000 ;
        RECT 73.545000 62.160000 73.745000 62.360000 ;
        RECT 73.545000 62.570000 73.745000 62.770000 ;
        RECT 73.545000 62.980000 73.745000 63.180000 ;
        RECT 73.545000 63.390000 73.745000 63.590000 ;
        RECT 73.545000 63.800000 73.745000 64.000000 ;
        RECT 73.545000 64.210000 73.745000 64.410000 ;
        RECT 73.545000 64.620000 73.745000 64.820000 ;
        RECT 73.545000 65.030000 73.745000 65.230000 ;
        RECT 73.545000 65.440000 73.745000 65.640000 ;
        RECT 73.545000 65.850000 73.745000 66.050000 ;
        RECT 73.545000 66.260000 73.745000 66.460000 ;
        RECT 73.955000 62.160000 74.155000 62.360000 ;
        RECT 73.955000 62.570000 74.155000 62.770000 ;
        RECT 73.955000 62.980000 74.155000 63.180000 ;
        RECT 73.955000 63.390000 74.155000 63.590000 ;
        RECT 73.955000 63.800000 74.155000 64.000000 ;
        RECT 73.955000 64.210000 74.155000 64.410000 ;
        RECT 73.955000 64.620000 74.155000 64.820000 ;
        RECT 73.955000 65.030000 74.155000 65.230000 ;
        RECT 73.955000 65.440000 74.155000 65.640000 ;
        RECT 73.955000 65.850000 74.155000 66.050000 ;
        RECT 73.955000 66.260000 74.155000 66.460000 ;
        RECT 74.365000 62.160000 74.565000 62.360000 ;
        RECT 74.365000 62.570000 74.565000 62.770000 ;
        RECT 74.365000 62.980000 74.565000 63.180000 ;
        RECT 74.365000 63.390000 74.565000 63.590000 ;
        RECT 74.365000 63.800000 74.565000 64.000000 ;
        RECT 74.365000 64.210000 74.565000 64.410000 ;
        RECT 74.365000 64.620000 74.565000 64.820000 ;
        RECT 74.365000 65.030000 74.565000 65.230000 ;
        RECT 74.365000 65.440000 74.565000 65.640000 ;
        RECT 74.365000 65.850000 74.565000 66.050000 ;
        RECT 74.365000 66.260000 74.565000 66.460000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000 24.900000   3.005000 ;
      RECT  0.000000   3.005000  3.005000  14.385000 ;
      RECT  0.000000  14.385000 24.900000  17.390000 ;
      RECT  0.000000  22.830000 24.900000  25.835000 ;
      RECT  0.000000  25.835000  3.005000  58.685000 ;
      RECT  0.000000  58.685000 24.900000  61.690000 ;
      RECT  0.000000  66.930000 24.895000  67.635000 ;
      RECT  0.000000  93.355000 60.885000  93.360000 ;
      RECT  0.000000  93.360000 18.610000  96.365000 ;
      RECT  0.000000  96.365000  3.005000 194.995000 ;
      RECT  0.000000 194.995000 24.895000 198.000000 ;
      RECT  3.000000   3.002000 72.000000  14.390000 ;
      RECT  3.000000  25.830000 72.000000  58.690000 ;
      RECT  3.000000  96.355000 59.640000  96.360000 ;
      RECT  3.000000  96.355000 59.640000  96.360000 ;
      RECT  3.000000  96.360000 72.000000 195.000000 ;
      RECT 14.395000  93.330000 60.860000  93.355000 ;
      RECT 14.545000  93.180000 60.710000  93.330000 ;
      RECT 14.695000  93.030000 60.560000  93.180000 ;
      RECT 14.845000  92.880000 60.410000  93.030000 ;
      RECT 14.995000  92.730000 60.260000  92.880000 ;
      RECT 15.145000  92.580000 60.110000  92.730000 ;
      RECT 15.295000  92.430000 59.960000  92.580000 ;
      RECT 15.445000  92.280000 59.810000  92.430000 ;
      RECT 15.595000  92.130000 59.660000  92.280000 ;
      RECT 15.745000  91.980000 59.510000  92.130000 ;
      RECT 15.745000  96.225000 59.510000  96.355000 ;
      RECT 15.745000  96.225000 59.510000  96.355000 ;
      RECT 15.895000  91.830000 59.360000  91.980000 ;
      RECT 15.895000  96.075000 59.360000  96.225000 ;
      RECT 15.895000  96.075000 59.360000  96.225000 ;
      RECT 16.045000  91.680000 59.210000  91.830000 ;
      RECT 16.045000  95.925000 59.210000  96.075000 ;
      RECT 16.045000  95.925000 59.210000  96.075000 ;
      RECT 16.195000  91.530000 59.060000  91.680000 ;
      RECT 16.195000  95.775000 59.060000  95.925000 ;
      RECT 16.195000  95.775000 59.060000  95.925000 ;
      RECT 16.345000  91.380000 58.910000  91.530000 ;
      RECT 16.345000  95.625000 58.910000  95.775000 ;
      RECT 16.345000  95.625000 58.910000  95.775000 ;
      RECT 16.495000  91.230000 58.760000  91.380000 ;
      RECT 16.495000  95.475000 58.760000  95.625000 ;
      RECT 16.495000  95.475000 58.760000  95.625000 ;
      RECT 16.645000  91.080000 58.610000  91.230000 ;
      RECT 16.645000  95.325000 58.610000  95.475000 ;
      RECT 16.645000  95.325000 58.610000  95.475000 ;
      RECT 16.795000  90.930000 58.460000  91.080000 ;
      RECT 16.795000  95.175000 58.460000  95.325000 ;
      RECT 16.795000  95.175000 58.460000  95.325000 ;
      RECT 16.945000  90.780000 58.310000  90.930000 ;
      RECT 16.945000  95.025000 58.310000  95.175000 ;
      RECT 16.945000  95.025000 58.310000  95.175000 ;
      RECT 17.095000  90.630000 58.160000  90.780000 ;
      RECT 17.095000  94.875000 58.160000  95.025000 ;
      RECT 17.095000  94.875000 58.160000  95.025000 ;
      RECT 17.245000  90.480000 58.010000  90.630000 ;
      RECT 17.245000  94.725000 58.010000  94.875000 ;
      RECT 17.245000  94.725000 58.010000  94.875000 ;
      RECT 17.395000  90.330000 57.860000  90.480000 ;
      RECT 17.395000  94.575000 57.860000  94.725000 ;
      RECT 17.395000  94.575000 57.860000  94.725000 ;
      RECT 17.545000  90.180000 57.710000  90.330000 ;
      RECT 17.545000  94.425000 57.710000  94.575000 ;
      RECT 17.545000  94.425000 57.710000  94.575000 ;
      RECT 17.695000  90.030000 57.560000  90.180000 ;
      RECT 17.695000  94.275000 57.560000  94.425000 ;
      RECT 17.695000  94.275000 57.560000  94.425000 ;
      RECT 17.845000  89.880000 57.410000  90.030000 ;
      RECT 17.845000  94.125000 57.410000  94.275000 ;
      RECT 17.845000  94.125000 57.410000  94.275000 ;
      RECT 17.995000  89.730000 57.260000  89.880000 ;
      RECT 17.995000  93.975000 57.260000  94.125000 ;
      RECT 17.995000  93.975000 57.260000  94.125000 ;
      RECT 18.145000  89.580000 57.110000  89.730000 ;
      RECT 18.145000  93.825000 57.110000  93.975000 ;
      RECT 18.145000  93.825000 57.110000  93.975000 ;
      RECT 18.295000  89.430000 56.960000  89.580000 ;
      RECT 18.295000  93.675000 56.960000  93.825000 ;
      RECT 18.295000  93.675000 56.960000  93.825000 ;
      RECT 18.445000  89.280000 56.810000  89.430000 ;
      RECT 18.445000  93.525000 56.810000  93.675000 ;
      RECT 18.445000  93.525000 56.810000  93.675000 ;
      RECT 18.595000  89.130000 56.660000  89.280000 ;
      RECT 18.595000  93.375000 56.660000  93.525000 ;
      RECT 18.595000  93.375000 56.660000  93.525000 ;
      RECT 18.745000  88.980000 56.510000  89.130000 ;
      RECT 18.745000  93.225000 56.510000  93.375000 ;
      RECT 18.745000  93.225000 56.510000  93.375000 ;
      RECT 18.895000  88.830000 56.360000  88.980000 ;
      RECT 18.895000  93.075000 56.360000  93.225000 ;
      RECT 18.895000  93.075000 56.360000  93.225000 ;
      RECT 19.045000  88.680000 56.210000  88.830000 ;
      RECT 19.045000  92.925000 56.210000  93.075000 ;
      RECT 19.045000  92.925000 56.210000  93.075000 ;
      RECT 19.195000  88.530000 56.060000  88.680000 ;
      RECT 19.195000  92.775000 56.060000  92.925000 ;
      RECT 19.195000  92.775000 56.060000  92.925000 ;
      RECT 19.345000  88.380000 55.910000  88.530000 ;
      RECT 19.345000  92.625000 55.910000  92.775000 ;
      RECT 19.345000  92.625000 55.910000  92.775000 ;
      RECT 19.495000  88.230000 55.760000  88.380000 ;
      RECT 19.495000  92.475000 55.760000  92.625000 ;
      RECT 19.495000  92.475000 55.760000  92.625000 ;
      RECT 19.645000  88.080000 55.610000  88.230000 ;
      RECT 19.645000  92.325000 55.610000  92.475000 ;
      RECT 19.645000  92.325000 55.610000  92.475000 ;
      RECT 19.795000  87.930000 55.460000  88.080000 ;
      RECT 19.795000  92.175000 55.460000  92.325000 ;
      RECT 19.795000  92.175000 55.460000  92.325000 ;
      RECT 19.945000  87.780000 55.310000  87.930000 ;
      RECT 19.945000  92.025000 55.310000  92.175000 ;
      RECT 19.945000  92.025000 55.310000  92.175000 ;
      RECT 20.095000  87.630000 55.160000  87.780000 ;
      RECT 20.095000  91.875000 55.160000  92.025000 ;
      RECT 20.095000  91.875000 55.160000  92.025000 ;
      RECT 20.245000  87.480000 55.010000  87.630000 ;
      RECT 20.245000  91.725000 55.010000  91.875000 ;
      RECT 20.245000  91.725000 55.010000  91.875000 ;
      RECT 20.395000  87.330000 54.860000  87.480000 ;
      RECT 20.395000  91.575000 54.860000  91.725000 ;
      RECT 20.395000  91.575000 54.860000  91.725000 ;
      RECT 20.545000  87.180000 54.710000  87.330000 ;
      RECT 20.545000  91.425000 54.710000  91.575000 ;
      RECT 20.545000  91.425000 54.710000  91.575000 ;
      RECT 20.695000  87.030000 54.560000  87.180000 ;
      RECT 20.695000  91.275000 54.560000  91.425000 ;
      RECT 20.695000  91.275000 54.560000  91.425000 ;
      RECT 20.845000  86.880000 54.410000  87.030000 ;
      RECT 20.845000  91.125000 54.410000  91.275000 ;
      RECT 20.845000  91.125000 54.410000  91.275000 ;
      RECT 20.995000  86.730000 54.260000  86.880000 ;
      RECT 20.995000  90.975000 54.260000  91.125000 ;
      RECT 20.995000  90.975000 54.260000  91.125000 ;
      RECT 21.145000  86.580000 54.110000  86.730000 ;
      RECT 21.145000  90.825000 54.110000  90.975000 ;
      RECT 21.145000  90.825000 54.110000  90.975000 ;
      RECT 21.295000  86.430000 53.960000  86.580000 ;
      RECT 21.295000  90.675000 53.960000  90.825000 ;
      RECT 21.295000  90.675000 53.960000  90.825000 ;
      RECT 21.445000  86.280000 53.810000  86.430000 ;
      RECT 21.445000  90.525000 53.810000  90.675000 ;
      RECT 21.445000  90.525000 53.810000  90.675000 ;
      RECT 21.595000  86.130000 53.660000  86.280000 ;
      RECT 21.595000  90.375000 53.660000  90.525000 ;
      RECT 21.595000  90.375000 53.660000  90.525000 ;
      RECT 21.745000  85.980000 53.510000  86.130000 ;
      RECT 21.745000  90.225000 53.510000  90.375000 ;
      RECT 21.745000  90.225000 53.510000  90.375000 ;
      RECT 21.895000  85.830000 53.360000  85.980000 ;
      RECT 21.895000  90.075000 53.360000  90.225000 ;
      RECT 21.895000  90.075000 53.360000  90.225000 ;
      RECT 22.045000  85.680000 53.210000  85.830000 ;
      RECT 22.045000  89.925000 53.210000  90.075000 ;
      RECT 22.045000  89.925000 53.210000  90.075000 ;
      RECT 22.195000  85.530000 53.060000  85.680000 ;
      RECT 22.195000  89.775000 53.060000  89.925000 ;
      RECT 22.195000  89.775000 53.060000  89.925000 ;
      RECT 22.345000  85.380000 52.910000  85.530000 ;
      RECT 22.345000  89.625000 52.910000  89.775000 ;
      RECT 22.345000  89.625000 52.910000  89.775000 ;
      RECT 22.495000  85.230000 52.760000  85.380000 ;
      RECT 22.495000  89.475000 52.760000  89.625000 ;
      RECT 22.495000  89.475000 52.760000  89.625000 ;
      RECT 22.645000  85.080000 52.610000  85.230000 ;
      RECT 22.645000  89.325000 52.610000  89.475000 ;
      RECT 22.645000  89.325000 52.610000  89.475000 ;
      RECT 22.795000  84.930000 52.460000  85.080000 ;
      RECT 22.795000  89.175000 52.460000  89.325000 ;
      RECT 22.795000  89.175000 52.460000  89.325000 ;
      RECT 22.945000  84.780000 52.310000  84.930000 ;
      RECT 22.945000  89.025000 52.310000  89.175000 ;
      RECT 22.945000  89.025000 52.310000  89.175000 ;
      RECT 23.095000  84.630000 52.160000  84.780000 ;
      RECT 23.095000  88.875000 52.160000  89.025000 ;
      RECT 23.095000  88.875000 52.160000  89.025000 ;
      RECT 23.245000  84.480000 52.010000  84.630000 ;
      RECT 23.245000  88.725000 52.010000  88.875000 ;
      RECT 23.245000  88.725000 52.010000  88.875000 ;
      RECT 23.395000  84.330000 51.860000  84.480000 ;
      RECT 23.395000  88.575000 51.860000  88.725000 ;
      RECT 23.395000  88.575000 51.860000  88.725000 ;
      RECT 23.545000  84.180000 51.710000  84.330000 ;
      RECT 23.545000  88.425000 51.710000  88.575000 ;
      RECT 23.545000  88.425000 51.710000  88.575000 ;
      RECT 23.695000  84.030000 51.560000  84.180000 ;
      RECT 23.695000  88.275000 51.560000  88.425000 ;
      RECT 23.695000  88.275000 51.560000  88.425000 ;
      RECT 23.845000  83.880000 51.410000  84.030000 ;
      RECT 23.845000  88.125000 51.410000  88.275000 ;
      RECT 23.845000  88.125000 51.410000  88.275000 ;
      RECT 23.995000  83.730000 51.260000  83.880000 ;
      RECT 23.995000  87.975000 51.260000  88.125000 ;
      RECT 23.995000  87.975000 51.260000  88.125000 ;
      RECT 24.145000  83.580000 51.110000  83.730000 ;
      RECT 24.145000  87.825000 51.110000  87.975000 ;
      RECT 24.145000  87.825000 51.110000  87.975000 ;
      RECT 24.295000  83.430000 50.960000  83.580000 ;
      RECT 24.295000  87.675000 50.960000  87.825000 ;
      RECT 24.295000  87.675000 50.960000  87.825000 ;
      RECT 24.445000  83.280000 50.810000  83.430000 ;
      RECT 24.445000  87.525000 50.810000  87.675000 ;
      RECT 24.445000  87.525000 50.810000  87.675000 ;
      RECT 24.595000  83.130000 50.660000  83.280000 ;
      RECT 24.595000  87.375000 50.660000  87.525000 ;
      RECT 24.595000  87.375000 50.660000  87.525000 ;
      RECT 24.745000  82.980000 50.510000  83.130000 ;
      RECT 24.745000  87.225000 50.510000  87.375000 ;
      RECT 24.745000  87.225000 50.510000  87.375000 ;
      RECT 24.895000  66.930000 50.360000 198.000000 ;
      RECT 24.895000  82.830000 50.360000  82.980000 ;
      RECT 24.895000  87.075000 50.360000  87.225000 ;
      RECT 24.895000  87.075000 50.360000  87.225000 ;
      RECT 24.900000   0.000000 50.355000 198.000000 ;
      RECT 24.900000   0.000000 50.355000 198.000000 ;
      RECT 25.045000  86.925000 50.210000  87.075000 ;
      RECT 25.045000  86.925000 50.210000  87.075000 ;
      RECT 25.195000  86.775000 50.060000  86.925000 ;
      RECT 25.195000  86.775000 50.060000  86.925000 ;
      RECT 25.345000  86.625000 49.910000  86.775000 ;
      RECT 25.345000  86.625000 49.910000  86.775000 ;
      RECT 25.495000  86.475000 49.760000  86.625000 ;
      RECT 25.495000  86.475000 49.760000  86.625000 ;
      RECT 25.645000  86.325000 49.610000  86.475000 ;
      RECT 25.645000  86.325000 49.610000  86.475000 ;
      RECT 25.795000  86.175000 49.460000  86.325000 ;
      RECT 25.795000  86.175000 49.460000  86.325000 ;
      RECT 25.945000  86.025000 49.310000  86.175000 ;
      RECT 25.945000  86.025000 49.310000  86.175000 ;
      RECT 26.095000  85.875000 49.160000  86.025000 ;
      RECT 26.095000  85.875000 49.160000  86.025000 ;
      RECT 26.245000  85.725000 49.010000  85.875000 ;
      RECT 26.245000  85.725000 49.010000  85.875000 ;
      RECT 26.395000  85.575000 48.860000  85.725000 ;
      RECT 26.395000  85.575000 48.860000  85.725000 ;
      RECT 26.545000  85.425000 48.710000  85.575000 ;
      RECT 26.545000  85.425000 48.710000  85.575000 ;
      RECT 26.695000  85.275000 48.560000  85.425000 ;
      RECT 26.695000  85.275000 48.560000  85.425000 ;
      RECT 26.845000  85.125000 48.410000  85.275000 ;
      RECT 26.845000  85.125000 48.410000  85.275000 ;
      RECT 26.995000  84.975000 48.260000  85.125000 ;
      RECT 26.995000  84.975000 48.260000  85.125000 ;
      RECT 27.145000  84.825000 48.110000  84.975000 ;
      RECT 27.145000  84.825000 48.110000  84.975000 ;
      RECT 27.295000  84.675000 47.960000  84.825000 ;
      RECT 27.295000  84.675000 47.960000  84.825000 ;
      RECT 27.445000  84.525000 47.810000  84.675000 ;
      RECT 27.445000  84.525000 47.810000  84.675000 ;
      RECT 27.595000  84.375000 47.660000  84.525000 ;
      RECT 27.595000  84.375000 47.660000  84.525000 ;
      RECT 27.745000  84.225000 47.510000  84.375000 ;
      RECT 27.745000  84.225000 47.510000  84.375000 ;
      RECT 27.895000  69.930000 47.360000  84.075000 ;
      RECT 27.895000  84.075000 47.360000  84.225000 ;
      RECT 27.895000  84.075000 47.360000  84.225000 ;
      RECT 27.900000  14.390000 47.355000  25.830000 ;
      RECT 27.900000  58.690000 47.355000  69.930000 ;
      RECT 50.355000   0.000000 75.000000   3.005000 ;
      RECT 50.355000  14.385000 75.000000  17.390000 ;
      RECT 50.355000  22.830000 75.000000  25.835000 ;
      RECT 50.355000  58.685000 75.000000  61.690000 ;
      RECT 50.360000  66.930000 75.000000  67.635000 ;
      RECT 50.360000 194.995000 75.000000 198.000000 ;
      RECT 56.645000  93.360000 75.000000  96.365000 ;
      RECT 71.995000   3.005000 75.000000  14.385000 ;
      RECT 71.995000  25.835000 75.000000  58.685000 ;
      RECT 71.995000  96.365000 75.000000 194.995000 ;
    LAYER met4 ;
      RECT  0.000000   5.885000 75.000000   6.485000 ;
      RECT  0.000000  11.935000  1.365000  12.535000 ;
      RECT  0.000000  16.785000  1.365000  17.385000 ;
      RECT  0.000000  22.835000  1.670000  23.435000 ;
      RECT  0.000000  28.885000  1.670000  29.485000 ;
      RECT  0.000000  33.735000  1.670000  34.335000 ;
      RECT  0.000000  38.585000  1.670000  39.185000 ;
      RECT  0.000000  44.635000  1.670000  45.335000 ;
      RECT  0.000000  55.135000  1.670000  55.835000 ;
      RECT  0.000000  61.085000  1.670000  61.685000 ;
      RECT  0.000000  66.935000 75.000000  67.635000 ;
      RECT  0.000000  93.400000 75.000000 173.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.670000   0.000000 73.330000   5.885000 ;
      RECT  1.670000   6.485000 73.330000  11.935000 ;
      RECT  1.670000  22.835000 73.330000  61.685000 ;
      RECT  1.670000  67.635000 73.330000  67.660000 ;
      RECT  1.670000  93.360000 60.750000  93.365000 ;
      RECT  1.670000  93.360000 60.750000 173.385000 ;
      RECT  1.670000  93.360000 60.750000 173.385000 ;
      RECT  1.670000  93.360000 60.750000 173.385000 ;
      RECT  1.670000  93.360000 60.750000 173.385000 ;
      RECT  1.670000  93.360000 60.750000 173.385000 ;
      RECT  1.670000  93.365000 73.330000  93.400000 ;
      RECT  1.670000  93.365000 73.330000 173.385000 ;
      RECT  1.670000  93.365000 73.330000 173.385000 ;
      RECT  1.670000  93.365000 73.330000 173.385000 ;
      RECT  1.670000  93.365000 73.330000 173.385000 ;
      RECT  1.670000  93.365000 73.330000 173.385000 ;
      RECT  1.670000 173.385000 73.330000 198.000000 ;
      RECT 14.505000  92.110000 60.750000  93.360000 ;
      RECT 14.505000  92.110000 60.750000 173.385000 ;
      RECT 14.505000  92.110000 60.750000 173.385000 ;
      RECT 14.505000  92.110000 60.750000 173.385000 ;
      RECT 14.505000  92.110000 60.750000 173.385000 ;
      RECT 14.505000  92.110000 60.750000 173.385000 ;
      RECT 15.765000  91.220000 59.490000  92.110000 ;
      RECT 16.650000  89.930000 58.605000  91.220000 ;
      RECT 17.925000  88.540000 57.330000  89.930000 ;
      RECT 19.255000  87.415000 56.000000  88.540000 ;
      RECT 20.465000  85.990000 54.790000  87.415000 ;
      RECT 21.850000  84.685000 53.405000  85.990000 ;
      RECT 21.850000  84.685000 53.405000  88.540000 ;
      RECT 23.170000  83.025000 52.085000  84.685000 ;
      RECT 23.170000  83.025000 52.085000  87.415000 ;
      RECT 24.875000  17.385000 50.380000  22.835000 ;
      RECT 24.875000  61.685000 50.380000  66.935000 ;
      RECT 24.900000  67.660000 50.355000  85.990000 ;
      RECT 24.900000  67.660000 50.355000  85.990000 ;
      RECT 24.900000  67.660000 50.355000  85.990000 ;
      RECT 73.330000  22.835000 75.000000  23.435000 ;
      RECT 73.330000  28.885000 75.000000  29.485000 ;
      RECT 73.330000  33.735000 75.000000  34.335000 ;
      RECT 73.330000  38.585000 75.000000  39.185000 ;
      RECT 73.330000  44.635000 75.000000  45.335000 ;
      RECT 73.330000  55.135000 75.000000  55.835000 ;
      RECT 73.330000  61.085000 75.000000  61.685000 ;
      RECT 73.635000  11.935000 75.000000  12.535000 ;
      RECT 73.635000  16.785000 75.000000  17.385000 ;
    LAYER met5 ;
      RECT 0.000000  93.785000 75.000000 172.985000 ;
      RECT 1.765000  12.235000 73.235000  17.085000 ;
      RECT 2.070000   0.000000 72.930000  12.235000 ;
      RECT 2.070000  17.085000 72.930000  93.785000 ;
      RECT 2.070000 172.985000 72.930000 198.000000 ;
  END
END sky130_fd_io__overlay_vddio_lvc


MACRO sky130_fd_io__overlay_vssd_hvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.970000 41.590000 24.395000 46.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 41.590000 74.290000 46.230000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 24.370000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
    PORT
      LAYER via3 ;
        RECT  1.060000 41.660000  1.260000 41.860000 ;
        RECT  1.060000 42.090000  1.260000 42.290000 ;
        RECT  1.060000 42.520000  1.260000 42.720000 ;
        RECT  1.060000 42.950000  1.260000 43.150000 ;
        RECT  1.060000 43.380000  1.260000 43.580000 ;
        RECT  1.060000 43.810000  1.260000 44.010000 ;
        RECT  1.060000 44.240000  1.260000 44.440000 ;
        RECT  1.060000 44.670000  1.260000 44.870000 ;
        RECT  1.060000 45.100000  1.260000 45.300000 ;
        RECT  1.060000 45.530000  1.260000 45.730000 ;
        RECT  1.060000 45.960000  1.260000 46.160000 ;
        RECT  1.465000 41.660000  1.665000 41.860000 ;
        RECT  1.465000 42.090000  1.665000 42.290000 ;
        RECT  1.465000 42.520000  1.665000 42.720000 ;
        RECT  1.465000 42.950000  1.665000 43.150000 ;
        RECT  1.465000 43.380000  1.665000 43.580000 ;
        RECT  1.465000 43.810000  1.665000 44.010000 ;
        RECT  1.465000 44.240000  1.665000 44.440000 ;
        RECT  1.465000 44.670000  1.665000 44.870000 ;
        RECT  1.465000 45.100000  1.665000 45.300000 ;
        RECT  1.465000 45.530000  1.665000 45.730000 ;
        RECT  1.465000 45.960000  1.665000 46.160000 ;
        RECT  1.870000 41.660000  2.070000 41.860000 ;
        RECT  1.870000 42.090000  2.070000 42.290000 ;
        RECT  1.870000 42.520000  2.070000 42.720000 ;
        RECT  1.870000 42.950000  2.070000 43.150000 ;
        RECT  1.870000 43.380000  2.070000 43.580000 ;
        RECT  1.870000 43.810000  2.070000 44.010000 ;
        RECT  1.870000 44.240000  2.070000 44.440000 ;
        RECT  1.870000 44.670000  2.070000 44.870000 ;
        RECT  1.870000 45.100000  2.070000 45.300000 ;
        RECT  1.870000 45.530000  2.070000 45.730000 ;
        RECT  1.870000 45.960000  2.070000 46.160000 ;
        RECT  2.275000 41.660000  2.475000 41.860000 ;
        RECT  2.275000 42.090000  2.475000 42.290000 ;
        RECT  2.275000 42.520000  2.475000 42.720000 ;
        RECT  2.275000 42.950000  2.475000 43.150000 ;
        RECT  2.275000 43.380000  2.475000 43.580000 ;
        RECT  2.275000 43.810000  2.475000 44.010000 ;
        RECT  2.275000 44.240000  2.475000 44.440000 ;
        RECT  2.275000 44.670000  2.475000 44.870000 ;
        RECT  2.275000 45.100000  2.475000 45.300000 ;
        RECT  2.275000 45.530000  2.475000 45.730000 ;
        RECT  2.275000 45.960000  2.475000 46.160000 ;
        RECT  2.680000 41.660000  2.880000 41.860000 ;
        RECT  2.680000 42.090000  2.880000 42.290000 ;
        RECT  2.680000 42.520000  2.880000 42.720000 ;
        RECT  2.680000 42.950000  2.880000 43.150000 ;
        RECT  2.680000 43.380000  2.880000 43.580000 ;
        RECT  2.680000 43.810000  2.880000 44.010000 ;
        RECT  2.680000 44.240000  2.880000 44.440000 ;
        RECT  2.680000 44.670000  2.880000 44.870000 ;
        RECT  2.680000 45.100000  2.880000 45.300000 ;
        RECT  2.680000 45.530000  2.880000 45.730000 ;
        RECT  2.680000 45.960000  2.880000 46.160000 ;
        RECT  3.085000 41.660000  3.285000 41.860000 ;
        RECT  3.085000 42.090000  3.285000 42.290000 ;
        RECT  3.085000 42.520000  3.285000 42.720000 ;
        RECT  3.085000 42.950000  3.285000 43.150000 ;
        RECT  3.085000 43.380000  3.285000 43.580000 ;
        RECT  3.085000 43.810000  3.285000 44.010000 ;
        RECT  3.085000 44.240000  3.285000 44.440000 ;
        RECT  3.085000 44.670000  3.285000 44.870000 ;
        RECT  3.085000 45.100000  3.285000 45.300000 ;
        RECT  3.085000 45.530000  3.285000 45.730000 ;
        RECT  3.085000 45.960000  3.285000 46.160000 ;
        RECT  3.490000 41.660000  3.690000 41.860000 ;
        RECT  3.490000 42.090000  3.690000 42.290000 ;
        RECT  3.490000 42.520000  3.690000 42.720000 ;
        RECT  3.490000 42.950000  3.690000 43.150000 ;
        RECT  3.490000 43.380000  3.690000 43.580000 ;
        RECT  3.490000 43.810000  3.690000 44.010000 ;
        RECT  3.490000 44.240000  3.690000 44.440000 ;
        RECT  3.490000 44.670000  3.690000 44.870000 ;
        RECT  3.490000 45.100000  3.690000 45.300000 ;
        RECT  3.490000 45.530000  3.690000 45.730000 ;
        RECT  3.490000 45.960000  3.690000 46.160000 ;
        RECT  3.895000 41.660000  4.095000 41.860000 ;
        RECT  3.895000 42.090000  4.095000 42.290000 ;
        RECT  3.895000 42.520000  4.095000 42.720000 ;
        RECT  3.895000 42.950000  4.095000 43.150000 ;
        RECT  3.895000 43.380000  4.095000 43.580000 ;
        RECT  3.895000 43.810000  4.095000 44.010000 ;
        RECT  3.895000 44.240000  4.095000 44.440000 ;
        RECT  3.895000 44.670000  4.095000 44.870000 ;
        RECT  3.895000 45.100000  4.095000 45.300000 ;
        RECT  3.895000 45.530000  4.095000 45.730000 ;
        RECT  3.895000 45.960000  4.095000 46.160000 ;
        RECT  4.300000 41.660000  4.500000 41.860000 ;
        RECT  4.300000 42.090000  4.500000 42.290000 ;
        RECT  4.300000 42.520000  4.500000 42.720000 ;
        RECT  4.300000 42.950000  4.500000 43.150000 ;
        RECT  4.300000 43.380000  4.500000 43.580000 ;
        RECT  4.300000 43.810000  4.500000 44.010000 ;
        RECT  4.300000 44.240000  4.500000 44.440000 ;
        RECT  4.300000 44.670000  4.500000 44.870000 ;
        RECT  4.300000 45.100000  4.500000 45.300000 ;
        RECT  4.300000 45.530000  4.500000 45.730000 ;
        RECT  4.300000 45.960000  4.500000 46.160000 ;
        RECT  4.705000 41.660000  4.905000 41.860000 ;
        RECT  4.705000 42.090000  4.905000 42.290000 ;
        RECT  4.705000 42.520000  4.905000 42.720000 ;
        RECT  4.705000 42.950000  4.905000 43.150000 ;
        RECT  4.705000 43.380000  4.905000 43.580000 ;
        RECT  4.705000 43.810000  4.905000 44.010000 ;
        RECT  4.705000 44.240000  4.905000 44.440000 ;
        RECT  4.705000 44.670000  4.905000 44.870000 ;
        RECT  4.705000 45.100000  4.905000 45.300000 ;
        RECT  4.705000 45.530000  4.905000 45.730000 ;
        RECT  4.705000 45.960000  4.905000 46.160000 ;
        RECT  5.110000 41.660000  5.310000 41.860000 ;
        RECT  5.110000 42.090000  5.310000 42.290000 ;
        RECT  5.110000 42.520000  5.310000 42.720000 ;
        RECT  5.110000 42.950000  5.310000 43.150000 ;
        RECT  5.110000 43.380000  5.310000 43.580000 ;
        RECT  5.110000 43.810000  5.310000 44.010000 ;
        RECT  5.110000 44.240000  5.310000 44.440000 ;
        RECT  5.110000 44.670000  5.310000 44.870000 ;
        RECT  5.110000 45.100000  5.310000 45.300000 ;
        RECT  5.110000 45.530000  5.310000 45.730000 ;
        RECT  5.110000 45.960000  5.310000 46.160000 ;
        RECT  5.515000 41.660000  5.715000 41.860000 ;
        RECT  5.515000 42.090000  5.715000 42.290000 ;
        RECT  5.515000 42.520000  5.715000 42.720000 ;
        RECT  5.515000 42.950000  5.715000 43.150000 ;
        RECT  5.515000 43.380000  5.715000 43.580000 ;
        RECT  5.515000 43.810000  5.715000 44.010000 ;
        RECT  5.515000 44.240000  5.715000 44.440000 ;
        RECT  5.515000 44.670000  5.715000 44.870000 ;
        RECT  5.515000 45.100000  5.715000 45.300000 ;
        RECT  5.515000 45.530000  5.715000 45.730000 ;
        RECT  5.515000 45.960000  5.715000 46.160000 ;
        RECT  5.920000 41.660000  6.120000 41.860000 ;
        RECT  5.920000 42.090000  6.120000 42.290000 ;
        RECT  5.920000 42.520000  6.120000 42.720000 ;
        RECT  5.920000 42.950000  6.120000 43.150000 ;
        RECT  5.920000 43.380000  6.120000 43.580000 ;
        RECT  5.920000 43.810000  6.120000 44.010000 ;
        RECT  5.920000 44.240000  6.120000 44.440000 ;
        RECT  5.920000 44.670000  6.120000 44.870000 ;
        RECT  5.920000 45.100000  6.120000 45.300000 ;
        RECT  5.920000 45.530000  6.120000 45.730000 ;
        RECT  5.920000 45.960000  6.120000 46.160000 ;
        RECT  6.325000 41.660000  6.525000 41.860000 ;
        RECT  6.325000 42.090000  6.525000 42.290000 ;
        RECT  6.325000 42.520000  6.525000 42.720000 ;
        RECT  6.325000 42.950000  6.525000 43.150000 ;
        RECT  6.325000 43.380000  6.525000 43.580000 ;
        RECT  6.325000 43.810000  6.525000 44.010000 ;
        RECT  6.325000 44.240000  6.525000 44.440000 ;
        RECT  6.325000 44.670000  6.525000 44.870000 ;
        RECT  6.325000 45.100000  6.525000 45.300000 ;
        RECT  6.325000 45.530000  6.525000 45.730000 ;
        RECT  6.325000 45.960000  6.525000 46.160000 ;
        RECT  6.730000 41.660000  6.930000 41.860000 ;
        RECT  6.730000 42.090000  6.930000 42.290000 ;
        RECT  6.730000 42.520000  6.930000 42.720000 ;
        RECT  6.730000 42.950000  6.930000 43.150000 ;
        RECT  6.730000 43.380000  6.930000 43.580000 ;
        RECT  6.730000 43.810000  6.930000 44.010000 ;
        RECT  6.730000 44.240000  6.930000 44.440000 ;
        RECT  6.730000 44.670000  6.930000 44.870000 ;
        RECT  6.730000 45.100000  6.930000 45.300000 ;
        RECT  6.730000 45.530000  6.930000 45.730000 ;
        RECT  6.730000 45.960000  6.930000 46.160000 ;
        RECT  7.135000 41.660000  7.335000 41.860000 ;
        RECT  7.135000 42.090000  7.335000 42.290000 ;
        RECT  7.135000 42.520000  7.335000 42.720000 ;
        RECT  7.135000 42.950000  7.335000 43.150000 ;
        RECT  7.135000 43.380000  7.335000 43.580000 ;
        RECT  7.135000 43.810000  7.335000 44.010000 ;
        RECT  7.135000 44.240000  7.335000 44.440000 ;
        RECT  7.135000 44.670000  7.335000 44.870000 ;
        RECT  7.135000 45.100000  7.335000 45.300000 ;
        RECT  7.135000 45.530000  7.335000 45.730000 ;
        RECT  7.135000 45.960000  7.335000 46.160000 ;
        RECT  7.540000 41.660000  7.740000 41.860000 ;
        RECT  7.540000 42.090000  7.740000 42.290000 ;
        RECT  7.540000 42.520000  7.740000 42.720000 ;
        RECT  7.540000 42.950000  7.740000 43.150000 ;
        RECT  7.540000 43.380000  7.740000 43.580000 ;
        RECT  7.540000 43.810000  7.740000 44.010000 ;
        RECT  7.540000 44.240000  7.740000 44.440000 ;
        RECT  7.540000 44.670000  7.740000 44.870000 ;
        RECT  7.540000 45.100000  7.740000 45.300000 ;
        RECT  7.540000 45.530000  7.740000 45.730000 ;
        RECT  7.540000 45.960000  7.740000 46.160000 ;
        RECT  7.945000 41.660000  8.145000 41.860000 ;
        RECT  7.945000 42.090000  8.145000 42.290000 ;
        RECT  7.945000 42.520000  8.145000 42.720000 ;
        RECT  7.945000 42.950000  8.145000 43.150000 ;
        RECT  7.945000 43.380000  8.145000 43.580000 ;
        RECT  7.945000 43.810000  8.145000 44.010000 ;
        RECT  7.945000 44.240000  8.145000 44.440000 ;
        RECT  7.945000 44.670000  8.145000 44.870000 ;
        RECT  7.945000 45.100000  8.145000 45.300000 ;
        RECT  7.945000 45.530000  8.145000 45.730000 ;
        RECT  7.945000 45.960000  8.145000 46.160000 ;
        RECT  8.350000 41.660000  8.550000 41.860000 ;
        RECT  8.350000 42.090000  8.550000 42.290000 ;
        RECT  8.350000 42.520000  8.550000 42.720000 ;
        RECT  8.350000 42.950000  8.550000 43.150000 ;
        RECT  8.350000 43.380000  8.550000 43.580000 ;
        RECT  8.350000 43.810000  8.550000 44.010000 ;
        RECT  8.350000 44.240000  8.550000 44.440000 ;
        RECT  8.350000 44.670000  8.550000 44.870000 ;
        RECT  8.350000 45.100000  8.550000 45.300000 ;
        RECT  8.350000 45.530000  8.550000 45.730000 ;
        RECT  8.350000 45.960000  8.550000 46.160000 ;
        RECT  8.755000 41.660000  8.955000 41.860000 ;
        RECT  8.755000 42.090000  8.955000 42.290000 ;
        RECT  8.755000 42.520000  8.955000 42.720000 ;
        RECT  8.755000 42.950000  8.955000 43.150000 ;
        RECT  8.755000 43.380000  8.955000 43.580000 ;
        RECT  8.755000 43.810000  8.955000 44.010000 ;
        RECT  8.755000 44.240000  8.955000 44.440000 ;
        RECT  8.755000 44.670000  8.955000 44.870000 ;
        RECT  8.755000 45.100000  8.955000 45.300000 ;
        RECT  8.755000 45.530000  8.955000 45.730000 ;
        RECT  8.755000 45.960000  8.955000 46.160000 ;
        RECT  9.160000 41.660000  9.360000 41.860000 ;
        RECT  9.160000 42.090000  9.360000 42.290000 ;
        RECT  9.160000 42.520000  9.360000 42.720000 ;
        RECT  9.160000 42.950000  9.360000 43.150000 ;
        RECT  9.160000 43.380000  9.360000 43.580000 ;
        RECT  9.160000 43.810000  9.360000 44.010000 ;
        RECT  9.160000 44.240000  9.360000 44.440000 ;
        RECT  9.160000 44.670000  9.360000 44.870000 ;
        RECT  9.160000 45.100000  9.360000 45.300000 ;
        RECT  9.160000 45.530000  9.360000 45.730000 ;
        RECT  9.160000 45.960000  9.360000 46.160000 ;
        RECT  9.565000 41.660000  9.765000 41.860000 ;
        RECT  9.565000 42.090000  9.765000 42.290000 ;
        RECT  9.565000 42.520000  9.765000 42.720000 ;
        RECT  9.565000 42.950000  9.765000 43.150000 ;
        RECT  9.565000 43.380000  9.765000 43.580000 ;
        RECT  9.565000 43.810000  9.765000 44.010000 ;
        RECT  9.565000 44.240000  9.765000 44.440000 ;
        RECT  9.565000 44.670000  9.765000 44.870000 ;
        RECT  9.565000 45.100000  9.765000 45.300000 ;
        RECT  9.565000 45.530000  9.765000 45.730000 ;
        RECT  9.565000 45.960000  9.765000 46.160000 ;
        RECT  9.970000 41.660000 10.170000 41.860000 ;
        RECT  9.970000 42.090000 10.170000 42.290000 ;
        RECT  9.970000 42.520000 10.170000 42.720000 ;
        RECT  9.970000 42.950000 10.170000 43.150000 ;
        RECT  9.970000 43.380000 10.170000 43.580000 ;
        RECT  9.970000 43.810000 10.170000 44.010000 ;
        RECT  9.970000 44.240000 10.170000 44.440000 ;
        RECT  9.970000 44.670000 10.170000 44.870000 ;
        RECT  9.970000 45.100000 10.170000 45.300000 ;
        RECT  9.970000 45.530000 10.170000 45.730000 ;
        RECT  9.970000 45.960000 10.170000 46.160000 ;
        RECT 10.375000 41.660000 10.575000 41.860000 ;
        RECT 10.375000 42.090000 10.575000 42.290000 ;
        RECT 10.375000 42.520000 10.575000 42.720000 ;
        RECT 10.375000 42.950000 10.575000 43.150000 ;
        RECT 10.375000 43.380000 10.575000 43.580000 ;
        RECT 10.375000 43.810000 10.575000 44.010000 ;
        RECT 10.375000 44.240000 10.575000 44.440000 ;
        RECT 10.375000 44.670000 10.575000 44.870000 ;
        RECT 10.375000 45.100000 10.575000 45.300000 ;
        RECT 10.375000 45.530000 10.575000 45.730000 ;
        RECT 10.375000 45.960000 10.575000 46.160000 ;
        RECT 10.780000 41.660000 10.980000 41.860000 ;
        RECT 10.780000 42.090000 10.980000 42.290000 ;
        RECT 10.780000 42.520000 10.980000 42.720000 ;
        RECT 10.780000 42.950000 10.980000 43.150000 ;
        RECT 10.780000 43.380000 10.980000 43.580000 ;
        RECT 10.780000 43.810000 10.980000 44.010000 ;
        RECT 10.780000 44.240000 10.980000 44.440000 ;
        RECT 10.780000 44.670000 10.980000 44.870000 ;
        RECT 10.780000 45.100000 10.980000 45.300000 ;
        RECT 10.780000 45.530000 10.980000 45.730000 ;
        RECT 10.780000 45.960000 10.980000 46.160000 ;
        RECT 11.185000 41.660000 11.385000 41.860000 ;
        RECT 11.185000 42.090000 11.385000 42.290000 ;
        RECT 11.185000 42.520000 11.385000 42.720000 ;
        RECT 11.185000 42.950000 11.385000 43.150000 ;
        RECT 11.185000 43.380000 11.385000 43.580000 ;
        RECT 11.185000 43.810000 11.385000 44.010000 ;
        RECT 11.185000 44.240000 11.385000 44.440000 ;
        RECT 11.185000 44.670000 11.385000 44.870000 ;
        RECT 11.185000 45.100000 11.385000 45.300000 ;
        RECT 11.185000 45.530000 11.385000 45.730000 ;
        RECT 11.185000 45.960000 11.385000 46.160000 ;
        RECT 11.590000 41.660000 11.790000 41.860000 ;
        RECT 11.590000 42.090000 11.790000 42.290000 ;
        RECT 11.590000 42.520000 11.790000 42.720000 ;
        RECT 11.590000 42.950000 11.790000 43.150000 ;
        RECT 11.590000 43.380000 11.790000 43.580000 ;
        RECT 11.590000 43.810000 11.790000 44.010000 ;
        RECT 11.590000 44.240000 11.790000 44.440000 ;
        RECT 11.590000 44.670000 11.790000 44.870000 ;
        RECT 11.590000 45.100000 11.790000 45.300000 ;
        RECT 11.590000 45.530000 11.790000 45.730000 ;
        RECT 11.590000 45.960000 11.790000 46.160000 ;
        RECT 11.995000 41.660000 12.195000 41.860000 ;
        RECT 11.995000 42.090000 12.195000 42.290000 ;
        RECT 11.995000 42.520000 12.195000 42.720000 ;
        RECT 11.995000 42.950000 12.195000 43.150000 ;
        RECT 11.995000 43.380000 12.195000 43.580000 ;
        RECT 11.995000 43.810000 12.195000 44.010000 ;
        RECT 11.995000 44.240000 12.195000 44.440000 ;
        RECT 11.995000 44.670000 12.195000 44.870000 ;
        RECT 11.995000 45.100000 12.195000 45.300000 ;
        RECT 11.995000 45.530000 12.195000 45.730000 ;
        RECT 11.995000 45.960000 12.195000 46.160000 ;
        RECT 12.400000 41.660000 12.600000 41.860000 ;
        RECT 12.400000 42.090000 12.600000 42.290000 ;
        RECT 12.400000 42.520000 12.600000 42.720000 ;
        RECT 12.400000 42.950000 12.600000 43.150000 ;
        RECT 12.400000 43.380000 12.600000 43.580000 ;
        RECT 12.400000 43.810000 12.600000 44.010000 ;
        RECT 12.400000 44.240000 12.600000 44.440000 ;
        RECT 12.400000 44.670000 12.600000 44.870000 ;
        RECT 12.400000 45.100000 12.600000 45.300000 ;
        RECT 12.400000 45.530000 12.600000 45.730000 ;
        RECT 12.400000 45.960000 12.600000 46.160000 ;
        RECT 12.805000 41.660000 13.005000 41.860000 ;
        RECT 12.805000 42.090000 13.005000 42.290000 ;
        RECT 12.805000 42.520000 13.005000 42.720000 ;
        RECT 12.805000 42.950000 13.005000 43.150000 ;
        RECT 12.805000 43.380000 13.005000 43.580000 ;
        RECT 12.805000 43.810000 13.005000 44.010000 ;
        RECT 12.805000 44.240000 13.005000 44.440000 ;
        RECT 12.805000 44.670000 13.005000 44.870000 ;
        RECT 12.805000 45.100000 13.005000 45.300000 ;
        RECT 12.805000 45.530000 13.005000 45.730000 ;
        RECT 12.805000 45.960000 13.005000 46.160000 ;
        RECT 13.210000 41.660000 13.410000 41.860000 ;
        RECT 13.210000 42.090000 13.410000 42.290000 ;
        RECT 13.210000 42.520000 13.410000 42.720000 ;
        RECT 13.210000 42.950000 13.410000 43.150000 ;
        RECT 13.210000 43.380000 13.410000 43.580000 ;
        RECT 13.210000 43.810000 13.410000 44.010000 ;
        RECT 13.210000 44.240000 13.410000 44.440000 ;
        RECT 13.210000 44.670000 13.410000 44.870000 ;
        RECT 13.210000 45.100000 13.410000 45.300000 ;
        RECT 13.210000 45.530000 13.410000 45.730000 ;
        RECT 13.210000 45.960000 13.410000 46.160000 ;
        RECT 13.615000 41.660000 13.815000 41.860000 ;
        RECT 13.615000 42.090000 13.815000 42.290000 ;
        RECT 13.615000 42.520000 13.815000 42.720000 ;
        RECT 13.615000 42.950000 13.815000 43.150000 ;
        RECT 13.615000 43.380000 13.815000 43.580000 ;
        RECT 13.615000 43.810000 13.815000 44.010000 ;
        RECT 13.615000 44.240000 13.815000 44.440000 ;
        RECT 13.615000 44.670000 13.815000 44.870000 ;
        RECT 13.615000 45.100000 13.815000 45.300000 ;
        RECT 13.615000 45.530000 13.815000 45.730000 ;
        RECT 13.615000 45.960000 13.815000 46.160000 ;
        RECT 14.020000 41.660000 14.220000 41.860000 ;
        RECT 14.020000 42.090000 14.220000 42.290000 ;
        RECT 14.020000 42.520000 14.220000 42.720000 ;
        RECT 14.020000 42.950000 14.220000 43.150000 ;
        RECT 14.020000 43.380000 14.220000 43.580000 ;
        RECT 14.020000 43.810000 14.220000 44.010000 ;
        RECT 14.020000 44.240000 14.220000 44.440000 ;
        RECT 14.020000 44.670000 14.220000 44.870000 ;
        RECT 14.020000 45.100000 14.220000 45.300000 ;
        RECT 14.020000 45.530000 14.220000 45.730000 ;
        RECT 14.020000 45.960000 14.220000 46.160000 ;
        RECT 14.425000 41.660000 14.625000 41.860000 ;
        RECT 14.425000 42.090000 14.625000 42.290000 ;
        RECT 14.425000 42.520000 14.625000 42.720000 ;
        RECT 14.425000 42.950000 14.625000 43.150000 ;
        RECT 14.425000 43.380000 14.625000 43.580000 ;
        RECT 14.425000 43.810000 14.625000 44.010000 ;
        RECT 14.425000 44.240000 14.625000 44.440000 ;
        RECT 14.425000 44.670000 14.625000 44.870000 ;
        RECT 14.425000 45.100000 14.625000 45.300000 ;
        RECT 14.425000 45.530000 14.625000 45.730000 ;
        RECT 14.425000 45.960000 14.625000 46.160000 ;
        RECT 14.830000 41.660000 15.030000 41.860000 ;
        RECT 14.830000 42.090000 15.030000 42.290000 ;
        RECT 14.830000 42.520000 15.030000 42.720000 ;
        RECT 14.830000 42.950000 15.030000 43.150000 ;
        RECT 14.830000 43.380000 15.030000 43.580000 ;
        RECT 14.830000 43.810000 15.030000 44.010000 ;
        RECT 14.830000 44.240000 15.030000 44.440000 ;
        RECT 14.830000 44.670000 15.030000 44.870000 ;
        RECT 14.830000 45.100000 15.030000 45.300000 ;
        RECT 14.830000 45.530000 15.030000 45.730000 ;
        RECT 14.830000 45.960000 15.030000 46.160000 ;
        RECT 15.235000 41.660000 15.435000 41.860000 ;
        RECT 15.235000 42.090000 15.435000 42.290000 ;
        RECT 15.235000 42.520000 15.435000 42.720000 ;
        RECT 15.235000 42.950000 15.435000 43.150000 ;
        RECT 15.235000 43.380000 15.435000 43.580000 ;
        RECT 15.235000 43.810000 15.435000 44.010000 ;
        RECT 15.235000 44.240000 15.435000 44.440000 ;
        RECT 15.235000 44.670000 15.435000 44.870000 ;
        RECT 15.235000 45.100000 15.435000 45.300000 ;
        RECT 15.235000 45.530000 15.435000 45.730000 ;
        RECT 15.235000 45.960000 15.435000 46.160000 ;
        RECT 15.640000 41.660000 15.840000 41.860000 ;
        RECT 15.640000 42.090000 15.840000 42.290000 ;
        RECT 15.640000 42.520000 15.840000 42.720000 ;
        RECT 15.640000 42.950000 15.840000 43.150000 ;
        RECT 15.640000 43.380000 15.840000 43.580000 ;
        RECT 15.640000 43.810000 15.840000 44.010000 ;
        RECT 15.640000 44.240000 15.840000 44.440000 ;
        RECT 15.640000 44.670000 15.840000 44.870000 ;
        RECT 15.640000 45.100000 15.840000 45.300000 ;
        RECT 15.640000 45.530000 15.840000 45.730000 ;
        RECT 15.640000 45.960000 15.840000 46.160000 ;
        RECT 16.045000 41.660000 16.245000 41.860000 ;
        RECT 16.045000 42.090000 16.245000 42.290000 ;
        RECT 16.045000 42.520000 16.245000 42.720000 ;
        RECT 16.045000 42.950000 16.245000 43.150000 ;
        RECT 16.045000 43.380000 16.245000 43.580000 ;
        RECT 16.045000 43.810000 16.245000 44.010000 ;
        RECT 16.045000 44.240000 16.245000 44.440000 ;
        RECT 16.045000 44.670000 16.245000 44.870000 ;
        RECT 16.045000 45.100000 16.245000 45.300000 ;
        RECT 16.045000 45.530000 16.245000 45.730000 ;
        RECT 16.045000 45.960000 16.245000 46.160000 ;
        RECT 16.450000 41.660000 16.650000 41.860000 ;
        RECT 16.450000 42.090000 16.650000 42.290000 ;
        RECT 16.450000 42.520000 16.650000 42.720000 ;
        RECT 16.450000 42.950000 16.650000 43.150000 ;
        RECT 16.450000 43.380000 16.650000 43.580000 ;
        RECT 16.450000 43.810000 16.650000 44.010000 ;
        RECT 16.450000 44.240000 16.650000 44.440000 ;
        RECT 16.450000 44.670000 16.650000 44.870000 ;
        RECT 16.450000 45.100000 16.650000 45.300000 ;
        RECT 16.450000 45.530000 16.650000 45.730000 ;
        RECT 16.450000 45.960000 16.650000 46.160000 ;
        RECT 16.855000 41.660000 17.055000 41.860000 ;
        RECT 16.855000 42.090000 17.055000 42.290000 ;
        RECT 16.855000 42.520000 17.055000 42.720000 ;
        RECT 16.855000 42.950000 17.055000 43.150000 ;
        RECT 16.855000 43.380000 17.055000 43.580000 ;
        RECT 16.855000 43.810000 17.055000 44.010000 ;
        RECT 16.855000 44.240000 17.055000 44.440000 ;
        RECT 16.855000 44.670000 17.055000 44.870000 ;
        RECT 16.855000 45.100000 17.055000 45.300000 ;
        RECT 16.855000 45.530000 17.055000 45.730000 ;
        RECT 16.855000 45.960000 17.055000 46.160000 ;
        RECT 17.260000 41.660000 17.460000 41.860000 ;
        RECT 17.260000 42.090000 17.460000 42.290000 ;
        RECT 17.260000 42.520000 17.460000 42.720000 ;
        RECT 17.260000 42.950000 17.460000 43.150000 ;
        RECT 17.260000 43.380000 17.460000 43.580000 ;
        RECT 17.260000 43.810000 17.460000 44.010000 ;
        RECT 17.260000 44.240000 17.460000 44.440000 ;
        RECT 17.260000 44.670000 17.460000 44.870000 ;
        RECT 17.260000 45.100000 17.460000 45.300000 ;
        RECT 17.260000 45.530000 17.460000 45.730000 ;
        RECT 17.260000 45.960000 17.460000 46.160000 ;
        RECT 17.665000 41.660000 17.865000 41.860000 ;
        RECT 17.665000 42.090000 17.865000 42.290000 ;
        RECT 17.665000 42.520000 17.865000 42.720000 ;
        RECT 17.665000 42.950000 17.865000 43.150000 ;
        RECT 17.665000 43.380000 17.865000 43.580000 ;
        RECT 17.665000 43.810000 17.865000 44.010000 ;
        RECT 17.665000 44.240000 17.865000 44.440000 ;
        RECT 17.665000 44.670000 17.865000 44.870000 ;
        RECT 17.665000 45.100000 17.865000 45.300000 ;
        RECT 17.665000 45.530000 17.865000 45.730000 ;
        RECT 17.665000 45.960000 17.865000 46.160000 ;
        RECT 18.070000 41.660000 18.270000 41.860000 ;
        RECT 18.070000 42.090000 18.270000 42.290000 ;
        RECT 18.070000 42.520000 18.270000 42.720000 ;
        RECT 18.070000 42.950000 18.270000 43.150000 ;
        RECT 18.070000 43.380000 18.270000 43.580000 ;
        RECT 18.070000 43.810000 18.270000 44.010000 ;
        RECT 18.070000 44.240000 18.270000 44.440000 ;
        RECT 18.070000 44.670000 18.270000 44.870000 ;
        RECT 18.070000 45.100000 18.270000 45.300000 ;
        RECT 18.070000 45.530000 18.270000 45.730000 ;
        RECT 18.070000 45.960000 18.270000 46.160000 ;
        RECT 18.475000 41.660000 18.675000 41.860000 ;
        RECT 18.475000 42.090000 18.675000 42.290000 ;
        RECT 18.475000 42.520000 18.675000 42.720000 ;
        RECT 18.475000 42.950000 18.675000 43.150000 ;
        RECT 18.475000 43.380000 18.675000 43.580000 ;
        RECT 18.475000 43.810000 18.675000 44.010000 ;
        RECT 18.475000 44.240000 18.675000 44.440000 ;
        RECT 18.475000 44.670000 18.675000 44.870000 ;
        RECT 18.475000 45.100000 18.675000 45.300000 ;
        RECT 18.475000 45.530000 18.675000 45.730000 ;
        RECT 18.475000 45.960000 18.675000 46.160000 ;
        RECT 18.880000 41.660000 19.080000 41.860000 ;
        RECT 18.880000 42.090000 19.080000 42.290000 ;
        RECT 18.880000 42.520000 19.080000 42.720000 ;
        RECT 18.880000 42.950000 19.080000 43.150000 ;
        RECT 18.880000 43.380000 19.080000 43.580000 ;
        RECT 18.880000 43.810000 19.080000 44.010000 ;
        RECT 18.880000 44.240000 19.080000 44.440000 ;
        RECT 18.880000 44.670000 19.080000 44.870000 ;
        RECT 18.880000 45.100000 19.080000 45.300000 ;
        RECT 18.880000 45.530000 19.080000 45.730000 ;
        RECT 18.880000 45.960000 19.080000 46.160000 ;
        RECT 19.285000 41.660000 19.485000 41.860000 ;
        RECT 19.285000 42.090000 19.485000 42.290000 ;
        RECT 19.285000 42.520000 19.485000 42.720000 ;
        RECT 19.285000 42.950000 19.485000 43.150000 ;
        RECT 19.285000 43.380000 19.485000 43.580000 ;
        RECT 19.285000 43.810000 19.485000 44.010000 ;
        RECT 19.285000 44.240000 19.485000 44.440000 ;
        RECT 19.285000 44.670000 19.485000 44.870000 ;
        RECT 19.285000 45.100000 19.485000 45.300000 ;
        RECT 19.285000 45.530000 19.485000 45.730000 ;
        RECT 19.285000 45.960000 19.485000 46.160000 ;
        RECT 19.690000 41.660000 19.890000 41.860000 ;
        RECT 19.690000 42.090000 19.890000 42.290000 ;
        RECT 19.690000 42.520000 19.890000 42.720000 ;
        RECT 19.690000 42.950000 19.890000 43.150000 ;
        RECT 19.690000 43.380000 19.890000 43.580000 ;
        RECT 19.690000 43.810000 19.890000 44.010000 ;
        RECT 19.690000 44.240000 19.890000 44.440000 ;
        RECT 19.690000 44.670000 19.890000 44.870000 ;
        RECT 19.690000 45.100000 19.890000 45.300000 ;
        RECT 19.690000 45.530000 19.890000 45.730000 ;
        RECT 19.690000 45.960000 19.890000 46.160000 ;
        RECT 20.095000 41.660000 20.295000 41.860000 ;
        RECT 20.095000 42.090000 20.295000 42.290000 ;
        RECT 20.095000 42.520000 20.295000 42.720000 ;
        RECT 20.095000 42.950000 20.295000 43.150000 ;
        RECT 20.095000 43.380000 20.295000 43.580000 ;
        RECT 20.095000 43.810000 20.295000 44.010000 ;
        RECT 20.095000 44.240000 20.295000 44.440000 ;
        RECT 20.095000 44.670000 20.295000 44.870000 ;
        RECT 20.095000 45.100000 20.295000 45.300000 ;
        RECT 20.095000 45.530000 20.295000 45.730000 ;
        RECT 20.095000 45.960000 20.295000 46.160000 ;
        RECT 20.500000 41.660000 20.700000 41.860000 ;
        RECT 20.500000 42.090000 20.700000 42.290000 ;
        RECT 20.500000 42.520000 20.700000 42.720000 ;
        RECT 20.500000 42.950000 20.700000 43.150000 ;
        RECT 20.500000 43.380000 20.700000 43.580000 ;
        RECT 20.500000 43.810000 20.700000 44.010000 ;
        RECT 20.500000 44.240000 20.700000 44.440000 ;
        RECT 20.500000 44.670000 20.700000 44.870000 ;
        RECT 20.500000 45.100000 20.700000 45.300000 ;
        RECT 20.500000 45.530000 20.700000 45.730000 ;
        RECT 20.500000 45.960000 20.700000 46.160000 ;
        RECT 20.905000 41.660000 21.105000 41.860000 ;
        RECT 20.905000 42.090000 21.105000 42.290000 ;
        RECT 20.905000 42.520000 21.105000 42.720000 ;
        RECT 20.905000 42.950000 21.105000 43.150000 ;
        RECT 20.905000 43.380000 21.105000 43.580000 ;
        RECT 20.905000 43.810000 21.105000 44.010000 ;
        RECT 20.905000 44.240000 21.105000 44.440000 ;
        RECT 20.905000 44.670000 21.105000 44.870000 ;
        RECT 20.905000 45.100000 21.105000 45.300000 ;
        RECT 20.905000 45.530000 21.105000 45.730000 ;
        RECT 20.905000 45.960000 21.105000 46.160000 ;
        RECT 21.305000 41.660000 21.505000 41.860000 ;
        RECT 21.305000 42.090000 21.505000 42.290000 ;
        RECT 21.305000 42.520000 21.505000 42.720000 ;
        RECT 21.305000 42.950000 21.505000 43.150000 ;
        RECT 21.305000 43.380000 21.505000 43.580000 ;
        RECT 21.305000 43.810000 21.505000 44.010000 ;
        RECT 21.305000 44.240000 21.505000 44.440000 ;
        RECT 21.305000 44.670000 21.505000 44.870000 ;
        RECT 21.305000 45.100000 21.505000 45.300000 ;
        RECT 21.305000 45.530000 21.505000 45.730000 ;
        RECT 21.305000 45.960000 21.505000 46.160000 ;
        RECT 21.705000 41.660000 21.905000 41.860000 ;
        RECT 21.705000 42.090000 21.905000 42.290000 ;
        RECT 21.705000 42.520000 21.905000 42.720000 ;
        RECT 21.705000 42.950000 21.905000 43.150000 ;
        RECT 21.705000 43.380000 21.905000 43.580000 ;
        RECT 21.705000 43.810000 21.905000 44.010000 ;
        RECT 21.705000 44.240000 21.905000 44.440000 ;
        RECT 21.705000 44.670000 21.905000 44.870000 ;
        RECT 21.705000 45.100000 21.905000 45.300000 ;
        RECT 21.705000 45.530000 21.905000 45.730000 ;
        RECT 21.705000 45.960000 21.905000 46.160000 ;
        RECT 22.105000 41.660000 22.305000 41.860000 ;
        RECT 22.105000 42.090000 22.305000 42.290000 ;
        RECT 22.105000 42.520000 22.305000 42.720000 ;
        RECT 22.105000 42.950000 22.305000 43.150000 ;
        RECT 22.105000 43.380000 22.305000 43.580000 ;
        RECT 22.105000 43.810000 22.305000 44.010000 ;
        RECT 22.105000 44.240000 22.305000 44.440000 ;
        RECT 22.105000 44.670000 22.305000 44.870000 ;
        RECT 22.105000 45.100000 22.305000 45.300000 ;
        RECT 22.105000 45.530000 22.305000 45.730000 ;
        RECT 22.105000 45.960000 22.305000 46.160000 ;
        RECT 22.505000 41.660000 22.705000 41.860000 ;
        RECT 22.505000 42.090000 22.705000 42.290000 ;
        RECT 22.505000 42.520000 22.705000 42.720000 ;
        RECT 22.505000 42.950000 22.705000 43.150000 ;
        RECT 22.505000 43.380000 22.705000 43.580000 ;
        RECT 22.505000 43.810000 22.705000 44.010000 ;
        RECT 22.505000 44.240000 22.705000 44.440000 ;
        RECT 22.505000 44.670000 22.705000 44.870000 ;
        RECT 22.505000 45.100000 22.705000 45.300000 ;
        RECT 22.505000 45.530000 22.705000 45.730000 ;
        RECT 22.505000 45.960000 22.705000 46.160000 ;
        RECT 22.905000 41.660000 23.105000 41.860000 ;
        RECT 22.905000 42.090000 23.105000 42.290000 ;
        RECT 22.905000 42.520000 23.105000 42.720000 ;
        RECT 22.905000 42.950000 23.105000 43.150000 ;
        RECT 22.905000 43.380000 23.105000 43.580000 ;
        RECT 22.905000 43.810000 23.105000 44.010000 ;
        RECT 22.905000 44.240000 23.105000 44.440000 ;
        RECT 22.905000 44.670000 23.105000 44.870000 ;
        RECT 22.905000 45.100000 23.105000 45.300000 ;
        RECT 22.905000 45.530000 23.105000 45.730000 ;
        RECT 22.905000 45.960000 23.105000 46.160000 ;
        RECT 23.305000 41.660000 23.505000 41.860000 ;
        RECT 23.305000 42.090000 23.505000 42.290000 ;
        RECT 23.305000 42.520000 23.505000 42.720000 ;
        RECT 23.305000 42.950000 23.505000 43.150000 ;
        RECT 23.305000 43.380000 23.505000 43.580000 ;
        RECT 23.305000 43.810000 23.505000 44.010000 ;
        RECT 23.305000 44.240000 23.505000 44.440000 ;
        RECT 23.305000 44.670000 23.505000 44.870000 ;
        RECT 23.305000 45.100000 23.505000 45.300000 ;
        RECT 23.305000 45.530000 23.505000 45.730000 ;
        RECT 23.305000 45.960000 23.505000 46.160000 ;
        RECT 23.705000 41.660000 23.905000 41.860000 ;
        RECT 23.705000 42.090000 23.905000 42.290000 ;
        RECT 23.705000 42.520000 23.905000 42.720000 ;
        RECT 23.705000 42.950000 23.905000 43.150000 ;
        RECT 23.705000 43.380000 23.905000 43.580000 ;
        RECT 23.705000 43.810000 23.905000 44.010000 ;
        RECT 23.705000 44.240000 23.905000 44.440000 ;
        RECT 23.705000 44.670000 23.905000 44.870000 ;
        RECT 23.705000 45.100000 23.905000 45.300000 ;
        RECT 23.705000 45.530000 23.905000 45.730000 ;
        RECT 23.705000 45.960000 23.905000 46.160000 ;
        RECT 24.105000 41.660000 24.305000 41.860000 ;
        RECT 24.105000 42.090000 24.305000 42.290000 ;
        RECT 24.105000 42.520000 24.305000 42.720000 ;
        RECT 24.105000 42.950000 24.305000 43.150000 ;
        RECT 24.105000 43.380000 24.305000 43.580000 ;
        RECT 24.105000 43.810000 24.305000 44.010000 ;
        RECT 24.105000 44.240000 24.305000 44.440000 ;
        RECT 24.105000 44.670000 24.305000 44.870000 ;
        RECT 24.105000 45.100000 24.305000 45.300000 ;
        RECT 24.105000 45.530000 24.305000 45.730000 ;
        RECT 24.105000 45.960000 24.305000 46.160000 ;
        RECT 50.480000 41.660000 50.680000 41.860000 ;
        RECT 50.480000 42.090000 50.680000 42.290000 ;
        RECT 50.480000 42.520000 50.680000 42.720000 ;
        RECT 50.480000 42.950000 50.680000 43.150000 ;
        RECT 50.480000 43.380000 50.680000 43.580000 ;
        RECT 50.480000 43.810000 50.680000 44.010000 ;
        RECT 50.480000 44.240000 50.680000 44.440000 ;
        RECT 50.480000 44.670000 50.680000 44.870000 ;
        RECT 50.480000 45.100000 50.680000 45.300000 ;
        RECT 50.480000 45.530000 50.680000 45.730000 ;
        RECT 50.480000 45.960000 50.680000 46.160000 ;
        RECT 50.890000 41.660000 51.090000 41.860000 ;
        RECT 50.890000 42.090000 51.090000 42.290000 ;
        RECT 50.890000 42.520000 51.090000 42.720000 ;
        RECT 50.890000 42.950000 51.090000 43.150000 ;
        RECT 50.890000 43.380000 51.090000 43.580000 ;
        RECT 50.890000 43.810000 51.090000 44.010000 ;
        RECT 50.890000 44.240000 51.090000 44.440000 ;
        RECT 50.890000 44.670000 51.090000 44.870000 ;
        RECT 50.890000 45.100000 51.090000 45.300000 ;
        RECT 50.890000 45.530000 51.090000 45.730000 ;
        RECT 50.890000 45.960000 51.090000 46.160000 ;
        RECT 51.300000 41.660000 51.500000 41.860000 ;
        RECT 51.300000 42.090000 51.500000 42.290000 ;
        RECT 51.300000 42.520000 51.500000 42.720000 ;
        RECT 51.300000 42.950000 51.500000 43.150000 ;
        RECT 51.300000 43.380000 51.500000 43.580000 ;
        RECT 51.300000 43.810000 51.500000 44.010000 ;
        RECT 51.300000 44.240000 51.500000 44.440000 ;
        RECT 51.300000 44.670000 51.500000 44.870000 ;
        RECT 51.300000 45.100000 51.500000 45.300000 ;
        RECT 51.300000 45.530000 51.500000 45.730000 ;
        RECT 51.300000 45.960000 51.500000 46.160000 ;
        RECT 51.710000 41.660000 51.910000 41.860000 ;
        RECT 51.710000 42.090000 51.910000 42.290000 ;
        RECT 51.710000 42.520000 51.910000 42.720000 ;
        RECT 51.710000 42.950000 51.910000 43.150000 ;
        RECT 51.710000 43.380000 51.910000 43.580000 ;
        RECT 51.710000 43.810000 51.910000 44.010000 ;
        RECT 51.710000 44.240000 51.910000 44.440000 ;
        RECT 51.710000 44.670000 51.910000 44.870000 ;
        RECT 51.710000 45.100000 51.910000 45.300000 ;
        RECT 51.710000 45.530000 51.910000 45.730000 ;
        RECT 51.710000 45.960000 51.910000 46.160000 ;
        RECT 52.120000 41.660000 52.320000 41.860000 ;
        RECT 52.120000 42.090000 52.320000 42.290000 ;
        RECT 52.120000 42.520000 52.320000 42.720000 ;
        RECT 52.120000 42.950000 52.320000 43.150000 ;
        RECT 52.120000 43.380000 52.320000 43.580000 ;
        RECT 52.120000 43.810000 52.320000 44.010000 ;
        RECT 52.120000 44.240000 52.320000 44.440000 ;
        RECT 52.120000 44.670000 52.320000 44.870000 ;
        RECT 52.120000 45.100000 52.320000 45.300000 ;
        RECT 52.120000 45.530000 52.320000 45.730000 ;
        RECT 52.120000 45.960000 52.320000 46.160000 ;
        RECT 52.530000 41.660000 52.730000 41.860000 ;
        RECT 52.530000 42.090000 52.730000 42.290000 ;
        RECT 52.530000 42.520000 52.730000 42.720000 ;
        RECT 52.530000 42.950000 52.730000 43.150000 ;
        RECT 52.530000 43.380000 52.730000 43.580000 ;
        RECT 52.530000 43.810000 52.730000 44.010000 ;
        RECT 52.530000 44.240000 52.730000 44.440000 ;
        RECT 52.530000 44.670000 52.730000 44.870000 ;
        RECT 52.530000 45.100000 52.730000 45.300000 ;
        RECT 52.530000 45.530000 52.730000 45.730000 ;
        RECT 52.530000 45.960000 52.730000 46.160000 ;
        RECT 52.940000 41.660000 53.140000 41.860000 ;
        RECT 52.940000 42.090000 53.140000 42.290000 ;
        RECT 52.940000 42.520000 53.140000 42.720000 ;
        RECT 52.940000 42.950000 53.140000 43.150000 ;
        RECT 52.940000 43.380000 53.140000 43.580000 ;
        RECT 52.940000 43.810000 53.140000 44.010000 ;
        RECT 52.940000 44.240000 53.140000 44.440000 ;
        RECT 52.940000 44.670000 53.140000 44.870000 ;
        RECT 52.940000 45.100000 53.140000 45.300000 ;
        RECT 52.940000 45.530000 53.140000 45.730000 ;
        RECT 52.940000 45.960000 53.140000 46.160000 ;
        RECT 53.345000 41.660000 53.545000 41.860000 ;
        RECT 53.345000 42.090000 53.545000 42.290000 ;
        RECT 53.345000 42.520000 53.545000 42.720000 ;
        RECT 53.345000 42.950000 53.545000 43.150000 ;
        RECT 53.345000 43.380000 53.545000 43.580000 ;
        RECT 53.345000 43.810000 53.545000 44.010000 ;
        RECT 53.345000 44.240000 53.545000 44.440000 ;
        RECT 53.345000 44.670000 53.545000 44.870000 ;
        RECT 53.345000 45.100000 53.545000 45.300000 ;
        RECT 53.345000 45.530000 53.545000 45.730000 ;
        RECT 53.345000 45.960000 53.545000 46.160000 ;
        RECT 53.750000 41.660000 53.950000 41.860000 ;
        RECT 53.750000 42.090000 53.950000 42.290000 ;
        RECT 53.750000 42.520000 53.950000 42.720000 ;
        RECT 53.750000 42.950000 53.950000 43.150000 ;
        RECT 53.750000 43.380000 53.950000 43.580000 ;
        RECT 53.750000 43.810000 53.950000 44.010000 ;
        RECT 53.750000 44.240000 53.950000 44.440000 ;
        RECT 53.750000 44.670000 53.950000 44.870000 ;
        RECT 53.750000 45.100000 53.950000 45.300000 ;
        RECT 53.750000 45.530000 53.950000 45.730000 ;
        RECT 53.750000 45.960000 53.950000 46.160000 ;
        RECT 54.155000 41.660000 54.355000 41.860000 ;
        RECT 54.155000 42.090000 54.355000 42.290000 ;
        RECT 54.155000 42.520000 54.355000 42.720000 ;
        RECT 54.155000 42.950000 54.355000 43.150000 ;
        RECT 54.155000 43.380000 54.355000 43.580000 ;
        RECT 54.155000 43.810000 54.355000 44.010000 ;
        RECT 54.155000 44.240000 54.355000 44.440000 ;
        RECT 54.155000 44.670000 54.355000 44.870000 ;
        RECT 54.155000 45.100000 54.355000 45.300000 ;
        RECT 54.155000 45.530000 54.355000 45.730000 ;
        RECT 54.155000 45.960000 54.355000 46.160000 ;
        RECT 54.560000 41.660000 54.760000 41.860000 ;
        RECT 54.560000 42.090000 54.760000 42.290000 ;
        RECT 54.560000 42.520000 54.760000 42.720000 ;
        RECT 54.560000 42.950000 54.760000 43.150000 ;
        RECT 54.560000 43.380000 54.760000 43.580000 ;
        RECT 54.560000 43.810000 54.760000 44.010000 ;
        RECT 54.560000 44.240000 54.760000 44.440000 ;
        RECT 54.560000 44.670000 54.760000 44.870000 ;
        RECT 54.560000 45.100000 54.760000 45.300000 ;
        RECT 54.560000 45.530000 54.760000 45.730000 ;
        RECT 54.560000 45.960000 54.760000 46.160000 ;
        RECT 54.965000 41.660000 55.165000 41.860000 ;
        RECT 54.965000 42.090000 55.165000 42.290000 ;
        RECT 54.965000 42.520000 55.165000 42.720000 ;
        RECT 54.965000 42.950000 55.165000 43.150000 ;
        RECT 54.965000 43.380000 55.165000 43.580000 ;
        RECT 54.965000 43.810000 55.165000 44.010000 ;
        RECT 54.965000 44.240000 55.165000 44.440000 ;
        RECT 54.965000 44.670000 55.165000 44.870000 ;
        RECT 54.965000 45.100000 55.165000 45.300000 ;
        RECT 54.965000 45.530000 55.165000 45.730000 ;
        RECT 54.965000 45.960000 55.165000 46.160000 ;
        RECT 55.370000 41.660000 55.570000 41.860000 ;
        RECT 55.370000 42.090000 55.570000 42.290000 ;
        RECT 55.370000 42.520000 55.570000 42.720000 ;
        RECT 55.370000 42.950000 55.570000 43.150000 ;
        RECT 55.370000 43.380000 55.570000 43.580000 ;
        RECT 55.370000 43.810000 55.570000 44.010000 ;
        RECT 55.370000 44.240000 55.570000 44.440000 ;
        RECT 55.370000 44.670000 55.570000 44.870000 ;
        RECT 55.370000 45.100000 55.570000 45.300000 ;
        RECT 55.370000 45.530000 55.570000 45.730000 ;
        RECT 55.370000 45.960000 55.570000 46.160000 ;
        RECT 55.775000 41.660000 55.975000 41.860000 ;
        RECT 55.775000 42.090000 55.975000 42.290000 ;
        RECT 55.775000 42.520000 55.975000 42.720000 ;
        RECT 55.775000 42.950000 55.975000 43.150000 ;
        RECT 55.775000 43.380000 55.975000 43.580000 ;
        RECT 55.775000 43.810000 55.975000 44.010000 ;
        RECT 55.775000 44.240000 55.975000 44.440000 ;
        RECT 55.775000 44.670000 55.975000 44.870000 ;
        RECT 55.775000 45.100000 55.975000 45.300000 ;
        RECT 55.775000 45.530000 55.975000 45.730000 ;
        RECT 55.775000 45.960000 55.975000 46.160000 ;
        RECT 56.180000 41.660000 56.380000 41.860000 ;
        RECT 56.180000 42.090000 56.380000 42.290000 ;
        RECT 56.180000 42.520000 56.380000 42.720000 ;
        RECT 56.180000 42.950000 56.380000 43.150000 ;
        RECT 56.180000 43.380000 56.380000 43.580000 ;
        RECT 56.180000 43.810000 56.380000 44.010000 ;
        RECT 56.180000 44.240000 56.380000 44.440000 ;
        RECT 56.180000 44.670000 56.380000 44.870000 ;
        RECT 56.180000 45.100000 56.380000 45.300000 ;
        RECT 56.180000 45.530000 56.380000 45.730000 ;
        RECT 56.180000 45.960000 56.380000 46.160000 ;
        RECT 56.585000 41.660000 56.785000 41.860000 ;
        RECT 56.585000 42.090000 56.785000 42.290000 ;
        RECT 56.585000 42.520000 56.785000 42.720000 ;
        RECT 56.585000 42.950000 56.785000 43.150000 ;
        RECT 56.585000 43.380000 56.785000 43.580000 ;
        RECT 56.585000 43.810000 56.785000 44.010000 ;
        RECT 56.585000 44.240000 56.785000 44.440000 ;
        RECT 56.585000 44.670000 56.785000 44.870000 ;
        RECT 56.585000 45.100000 56.785000 45.300000 ;
        RECT 56.585000 45.530000 56.785000 45.730000 ;
        RECT 56.585000 45.960000 56.785000 46.160000 ;
        RECT 56.990000 41.660000 57.190000 41.860000 ;
        RECT 56.990000 42.090000 57.190000 42.290000 ;
        RECT 56.990000 42.520000 57.190000 42.720000 ;
        RECT 56.990000 42.950000 57.190000 43.150000 ;
        RECT 56.990000 43.380000 57.190000 43.580000 ;
        RECT 56.990000 43.810000 57.190000 44.010000 ;
        RECT 56.990000 44.240000 57.190000 44.440000 ;
        RECT 56.990000 44.670000 57.190000 44.870000 ;
        RECT 56.990000 45.100000 57.190000 45.300000 ;
        RECT 56.990000 45.530000 57.190000 45.730000 ;
        RECT 56.990000 45.960000 57.190000 46.160000 ;
        RECT 57.395000 41.660000 57.595000 41.860000 ;
        RECT 57.395000 42.090000 57.595000 42.290000 ;
        RECT 57.395000 42.520000 57.595000 42.720000 ;
        RECT 57.395000 42.950000 57.595000 43.150000 ;
        RECT 57.395000 43.380000 57.595000 43.580000 ;
        RECT 57.395000 43.810000 57.595000 44.010000 ;
        RECT 57.395000 44.240000 57.595000 44.440000 ;
        RECT 57.395000 44.670000 57.595000 44.870000 ;
        RECT 57.395000 45.100000 57.595000 45.300000 ;
        RECT 57.395000 45.530000 57.595000 45.730000 ;
        RECT 57.395000 45.960000 57.595000 46.160000 ;
        RECT 57.800000 41.660000 58.000000 41.860000 ;
        RECT 57.800000 42.090000 58.000000 42.290000 ;
        RECT 57.800000 42.520000 58.000000 42.720000 ;
        RECT 57.800000 42.950000 58.000000 43.150000 ;
        RECT 57.800000 43.380000 58.000000 43.580000 ;
        RECT 57.800000 43.810000 58.000000 44.010000 ;
        RECT 57.800000 44.240000 58.000000 44.440000 ;
        RECT 57.800000 44.670000 58.000000 44.870000 ;
        RECT 57.800000 45.100000 58.000000 45.300000 ;
        RECT 57.800000 45.530000 58.000000 45.730000 ;
        RECT 57.800000 45.960000 58.000000 46.160000 ;
        RECT 58.205000 41.660000 58.405000 41.860000 ;
        RECT 58.205000 42.090000 58.405000 42.290000 ;
        RECT 58.205000 42.520000 58.405000 42.720000 ;
        RECT 58.205000 42.950000 58.405000 43.150000 ;
        RECT 58.205000 43.380000 58.405000 43.580000 ;
        RECT 58.205000 43.810000 58.405000 44.010000 ;
        RECT 58.205000 44.240000 58.405000 44.440000 ;
        RECT 58.205000 44.670000 58.405000 44.870000 ;
        RECT 58.205000 45.100000 58.405000 45.300000 ;
        RECT 58.205000 45.530000 58.405000 45.730000 ;
        RECT 58.205000 45.960000 58.405000 46.160000 ;
        RECT 58.610000 41.660000 58.810000 41.860000 ;
        RECT 58.610000 42.090000 58.810000 42.290000 ;
        RECT 58.610000 42.520000 58.810000 42.720000 ;
        RECT 58.610000 42.950000 58.810000 43.150000 ;
        RECT 58.610000 43.380000 58.810000 43.580000 ;
        RECT 58.610000 43.810000 58.810000 44.010000 ;
        RECT 58.610000 44.240000 58.810000 44.440000 ;
        RECT 58.610000 44.670000 58.810000 44.870000 ;
        RECT 58.610000 45.100000 58.810000 45.300000 ;
        RECT 58.610000 45.530000 58.810000 45.730000 ;
        RECT 58.610000 45.960000 58.810000 46.160000 ;
        RECT 59.015000 41.660000 59.215000 41.860000 ;
        RECT 59.015000 42.090000 59.215000 42.290000 ;
        RECT 59.015000 42.520000 59.215000 42.720000 ;
        RECT 59.015000 42.950000 59.215000 43.150000 ;
        RECT 59.015000 43.380000 59.215000 43.580000 ;
        RECT 59.015000 43.810000 59.215000 44.010000 ;
        RECT 59.015000 44.240000 59.215000 44.440000 ;
        RECT 59.015000 44.670000 59.215000 44.870000 ;
        RECT 59.015000 45.100000 59.215000 45.300000 ;
        RECT 59.015000 45.530000 59.215000 45.730000 ;
        RECT 59.015000 45.960000 59.215000 46.160000 ;
        RECT 59.420000 41.660000 59.620000 41.860000 ;
        RECT 59.420000 42.090000 59.620000 42.290000 ;
        RECT 59.420000 42.520000 59.620000 42.720000 ;
        RECT 59.420000 42.950000 59.620000 43.150000 ;
        RECT 59.420000 43.380000 59.620000 43.580000 ;
        RECT 59.420000 43.810000 59.620000 44.010000 ;
        RECT 59.420000 44.240000 59.620000 44.440000 ;
        RECT 59.420000 44.670000 59.620000 44.870000 ;
        RECT 59.420000 45.100000 59.620000 45.300000 ;
        RECT 59.420000 45.530000 59.620000 45.730000 ;
        RECT 59.420000 45.960000 59.620000 46.160000 ;
        RECT 59.825000 41.660000 60.025000 41.860000 ;
        RECT 59.825000 42.090000 60.025000 42.290000 ;
        RECT 59.825000 42.520000 60.025000 42.720000 ;
        RECT 59.825000 42.950000 60.025000 43.150000 ;
        RECT 59.825000 43.380000 60.025000 43.580000 ;
        RECT 59.825000 43.810000 60.025000 44.010000 ;
        RECT 59.825000 44.240000 60.025000 44.440000 ;
        RECT 59.825000 44.670000 60.025000 44.870000 ;
        RECT 59.825000 45.100000 60.025000 45.300000 ;
        RECT 59.825000 45.530000 60.025000 45.730000 ;
        RECT 59.825000 45.960000 60.025000 46.160000 ;
        RECT 60.230000 41.660000 60.430000 41.860000 ;
        RECT 60.230000 42.090000 60.430000 42.290000 ;
        RECT 60.230000 42.520000 60.430000 42.720000 ;
        RECT 60.230000 42.950000 60.430000 43.150000 ;
        RECT 60.230000 43.380000 60.430000 43.580000 ;
        RECT 60.230000 43.810000 60.430000 44.010000 ;
        RECT 60.230000 44.240000 60.430000 44.440000 ;
        RECT 60.230000 44.670000 60.430000 44.870000 ;
        RECT 60.230000 45.100000 60.430000 45.300000 ;
        RECT 60.230000 45.530000 60.430000 45.730000 ;
        RECT 60.230000 45.960000 60.430000 46.160000 ;
        RECT 60.635000 41.660000 60.835000 41.860000 ;
        RECT 60.635000 42.090000 60.835000 42.290000 ;
        RECT 60.635000 42.520000 60.835000 42.720000 ;
        RECT 60.635000 42.950000 60.835000 43.150000 ;
        RECT 60.635000 43.380000 60.835000 43.580000 ;
        RECT 60.635000 43.810000 60.835000 44.010000 ;
        RECT 60.635000 44.240000 60.835000 44.440000 ;
        RECT 60.635000 44.670000 60.835000 44.870000 ;
        RECT 60.635000 45.100000 60.835000 45.300000 ;
        RECT 60.635000 45.530000 60.835000 45.730000 ;
        RECT 60.635000 45.960000 60.835000 46.160000 ;
        RECT 61.040000 41.660000 61.240000 41.860000 ;
        RECT 61.040000 42.090000 61.240000 42.290000 ;
        RECT 61.040000 42.520000 61.240000 42.720000 ;
        RECT 61.040000 42.950000 61.240000 43.150000 ;
        RECT 61.040000 43.380000 61.240000 43.580000 ;
        RECT 61.040000 43.810000 61.240000 44.010000 ;
        RECT 61.040000 44.240000 61.240000 44.440000 ;
        RECT 61.040000 44.670000 61.240000 44.870000 ;
        RECT 61.040000 45.100000 61.240000 45.300000 ;
        RECT 61.040000 45.530000 61.240000 45.730000 ;
        RECT 61.040000 45.960000 61.240000 46.160000 ;
        RECT 61.445000 41.660000 61.645000 41.860000 ;
        RECT 61.445000 42.090000 61.645000 42.290000 ;
        RECT 61.445000 42.520000 61.645000 42.720000 ;
        RECT 61.445000 42.950000 61.645000 43.150000 ;
        RECT 61.445000 43.380000 61.645000 43.580000 ;
        RECT 61.445000 43.810000 61.645000 44.010000 ;
        RECT 61.445000 44.240000 61.645000 44.440000 ;
        RECT 61.445000 44.670000 61.645000 44.870000 ;
        RECT 61.445000 45.100000 61.645000 45.300000 ;
        RECT 61.445000 45.530000 61.645000 45.730000 ;
        RECT 61.445000 45.960000 61.645000 46.160000 ;
        RECT 61.850000 41.660000 62.050000 41.860000 ;
        RECT 61.850000 42.090000 62.050000 42.290000 ;
        RECT 61.850000 42.520000 62.050000 42.720000 ;
        RECT 61.850000 42.950000 62.050000 43.150000 ;
        RECT 61.850000 43.380000 62.050000 43.580000 ;
        RECT 61.850000 43.810000 62.050000 44.010000 ;
        RECT 61.850000 44.240000 62.050000 44.440000 ;
        RECT 61.850000 44.670000 62.050000 44.870000 ;
        RECT 61.850000 45.100000 62.050000 45.300000 ;
        RECT 61.850000 45.530000 62.050000 45.730000 ;
        RECT 61.850000 45.960000 62.050000 46.160000 ;
        RECT 62.255000 41.660000 62.455000 41.860000 ;
        RECT 62.255000 42.090000 62.455000 42.290000 ;
        RECT 62.255000 42.520000 62.455000 42.720000 ;
        RECT 62.255000 42.950000 62.455000 43.150000 ;
        RECT 62.255000 43.380000 62.455000 43.580000 ;
        RECT 62.255000 43.810000 62.455000 44.010000 ;
        RECT 62.255000 44.240000 62.455000 44.440000 ;
        RECT 62.255000 44.670000 62.455000 44.870000 ;
        RECT 62.255000 45.100000 62.455000 45.300000 ;
        RECT 62.255000 45.530000 62.455000 45.730000 ;
        RECT 62.255000 45.960000 62.455000 46.160000 ;
        RECT 62.660000 41.660000 62.860000 41.860000 ;
        RECT 62.660000 42.090000 62.860000 42.290000 ;
        RECT 62.660000 42.520000 62.860000 42.720000 ;
        RECT 62.660000 42.950000 62.860000 43.150000 ;
        RECT 62.660000 43.380000 62.860000 43.580000 ;
        RECT 62.660000 43.810000 62.860000 44.010000 ;
        RECT 62.660000 44.240000 62.860000 44.440000 ;
        RECT 62.660000 44.670000 62.860000 44.870000 ;
        RECT 62.660000 45.100000 62.860000 45.300000 ;
        RECT 62.660000 45.530000 62.860000 45.730000 ;
        RECT 62.660000 45.960000 62.860000 46.160000 ;
        RECT 63.065000 41.660000 63.265000 41.860000 ;
        RECT 63.065000 42.090000 63.265000 42.290000 ;
        RECT 63.065000 42.520000 63.265000 42.720000 ;
        RECT 63.065000 42.950000 63.265000 43.150000 ;
        RECT 63.065000 43.380000 63.265000 43.580000 ;
        RECT 63.065000 43.810000 63.265000 44.010000 ;
        RECT 63.065000 44.240000 63.265000 44.440000 ;
        RECT 63.065000 44.670000 63.265000 44.870000 ;
        RECT 63.065000 45.100000 63.265000 45.300000 ;
        RECT 63.065000 45.530000 63.265000 45.730000 ;
        RECT 63.065000 45.960000 63.265000 46.160000 ;
        RECT 63.470000 41.660000 63.670000 41.860000 ;
        RECT 63.470000 42.090000 63.670000 42.290000 ;
        RECT 63.470000 42.520000 63.670000 42.720000 ;
        RECT 63.470000 42.950000 63.670000 43.150000 ;
        RECT 63.470000 43.380000 63.670000 43.580000 ;
        RECT 63.470000 43.810000 63.670000 44.010000 ;
        RECT 63.470000 44.240000 63.670000 44.440000 ;
        RECT 63.470000 44.670000 63.670000 44.870000 ;
        RECT 63.470000 45.100000 63.670000 45.300000 ;
        RECT 63.470000 45.530000 63.670000 45.730000 ;
        RECT 63.470000 45.960000 63.670000 46.160000 ;
        RECT 63.875000 41.660000 64.075000 41.860000 ;
        RECT 63.875000 42.090000 64.075000 42.290000 ;
        RECT 63.875000 42.520000 64.075000 42.720000 ;
        RECT 63.875000 42.950000 64.075000 43.150000 ;
        RECT 63.875000 43.380000 64.075000 43.580000 ;
        RECT 63.875000 43.810000 64.075000 44.010000 ;
        RECT 63.875000 44.240000 64.075000 44.440000 ;
        RECT 63.875000 44.670000 64.075000 44.870000 ;
        RECT 63.875000 45.100000 64.075000 45.300000 ;
        RECT 63.875000 45.530000 64.075000 45.730000 ;
        RECT 63.875000 45.960000 64.075000 46.160000 ;
        RECT 64.280000 41.660000 64.480000 41.860000 ;
        RECT 64.280000 42.090000 64.480000 42.290000 ;
        RECT 64.280000 42.520000 64.480000 42.720000 ;
        RECT 64.280000 42.950000 64.480000 43.150000 ;
        RECT 64.280000 43.380000 64.480000 43.580000 ;
        RECT 64.280000 43.810000 64.480000 44.010000 ;
        RECT 64.280000 44.240000 64.480000 44.440000 ;
        RECT 64.280000 44.670000 64.480000 44.870000 ;
        RECT 64.280000 45.100000 64.480000 45.300000 ;
        RECT 64.280000 45.530000 64.480000 45.730000 ;
        RECT 64.280000 45.960000 64.480000 46.160000 ;
        RECT 64.685000 41.660000 64.885000 41.860000 ;
        RECT 64.685000 42.090000 64.885000 42.290000 ;
        RECT 64.685000 42.520000 64.885000 42.720000 ;
        RECT 64.685000 42.950000 64.885000 43.150000 ;
        RECT 64.685000 43.380000 64.885000 43.580000 ;
        RECT 64.685000 43.810000 64.885000 44.010000 ;
        RECT 64.685000 44.240000 64.885000 44.440000 ;
        RECT 64.685000 44.670000 64.885000 44.870000 ;
        RECT 64.685000 45.100000 64.885000 45.300000 ;
        RECT 64.685000 45.530000 64.885000 45.730000 ;
        RECT 64.685000 45.960000 64.885000 46.160000 ;
        RECT 65.090000 41.660000 65.290000 41.860000 ;
        RECT 65.090000 42.090000 65.290000 42.290000 ;
        RECT 65.090000 42.520000 65.290000 42.720000 ;
        RECT 65.090000 42.950000 65.290000 43.150000 ;
        RECT 65.090000 43.380000 65.290000 43.580000 ;
        RECT 65.090000 43.810000 65.290000 44.010000 ;
        RECT 65.090000 44.240000 65.290000 44.440000 ;
        RECT 65.090000 44.670000 65.290000 44.870000 ;
        RECT 65.090000 45.100000 65.290000 45.300000 ;
        RECT 65.090000 45.530000 65.290000 45.730000 ;
        RECT 65.090000 45.960000 65.290000 46.160000 ;
        RECT 65.495000 41.660000 65.695000 41.860000 ;
        RECT 65.495000 42.090000 65.695000 42.290000 ;
        RECT 65.495000 42.520000 65.695000 42.720000 ;
        RECT 65.495000 42.950000 65.695000 43.150000 ;
        RECT 65.495000 43.380000 65.695000 43.580000 ;
        RECT 65.495000 43.810000 65.695000 44.010000 ;
        RECT 65.495000 44.240000 65.695000 44.440000 ;
        RECT 65.495000 44.670000 65.695000 44.870000 ;
        RECT 65.495000 45.100000 65.695000 45.300000 ;
        RECT 65.495000 45.530000 65.695000 45.730000 ;
        RECT 65.495000 45.960000 65.695000 46.160000 ;
        RECT 65.900000 41.660000 66.100000 41.860000 ;
        RECT 65.900000 42.090000 66.100000 42.290000 ;
        RECT 65.900000 42.520000 66.100000 42.720000 ;
        RECT 65.900000 42.950000 66.100000 43.150000 ;
        RECT 65.900000 43.380000 66.100000 43.580000 ;
        RECT 65.900000 43.810000 66.100000 44.010000 ;
        RECT 65.900000 44.240000 66.100000 44.440000 ;
        RECT 65.900000 44.670000 66.100000 44.870000 ;
        RECT 65.900000 45.100000 66.100000 45.300000 ;
        RECT 65.900000 45.530000 66.100000 45.730000 ;
        RECT 65.900000 45.960000 66.100000 46.160000 ;
        RECT 66.305000 41.660000 66.505000 41.860000 ;
        RECT 66.305000 42.090000 66.505000 42.290000 ;
        RECT 66.305000 42.520000 66.505000 42.720000 ;
        RECT 66.305000 42.950000 66.505000 43.150000 ;
        RECT 66.305000 43.380000 66.505000 43.580000 ;
        RECT 66.305000 43.810000 66.505000 44.010000 ;
        RECT 66.305000 44.240000 66.505000 44.440000 ;
        RECT 66.305000 44.670000 66.505000 44.870000 ;
        RECT 66.305000 45.100000 66.505000 45.300000 ;
        RECT 66.305000 45.530000 66.505000 45.730000 ;
        RECT 66.305000 45.960000 66.505000 46.160000 ;
        RECT 66.710000 41.660000 66.910000 41.860000 ;
        RECT 66.710000 42.090000 66.910000 42.290000 ;
        RECT 66.710000 42.520000 66.910000 42.720000 ;
        RECT 66.710000 42.950000 66.910000 43.150000 ;
        RECT 66.710000 43.380000 66.910000 43.580000 ;
        RECT 66.710000 43.810000 66.910000 44.010000 ;
        RECT 66.710000 44.240000 66.910000 44.440000 ;
        RECT 66.710000 44.670000 66.910000 44.870000 ;
        RECT 66.710000 45.100000 66.910000 45.300000 ;
        RECT 66.710000 45.530000 66.910000 45.730000 ;
        RECT 66.710000 45.960000 66.910000 46.160000 ;
        RECT 67.115000 41.660000 67.315000 41.860000 ;
        RECT 67.115000 42.090000 67.315000 42.290000 ;
        RECT 67.115000 42.520000 67.315000 42.720000 ;
        RECT 67.115000 42.950000 67.315000 43.150000 ;
        RECT 67.115000 43.380000 67.315000 43.580000 ;
        RECT 67.115000 43.810000 67.315000 44.010000 ;
        RECT 67.115000 44.240000 67.315000 44.440000 ;
        RECT 67.115000 44.670000 67.315000 44.870000 ;
        RECT 67.115000 45.100000 67.315000 45.300000 ;
        RECT 67.115000 45.530000 67.315000 45.730000 ;
        RECT 67.115000 45.960000 67.315000 46.160000 ;
        RECT 67.520000 41.660000 67.720000 41.860000 ;
        RECT 67.520000 42.090000 67.720000 42.290000 ;
        RECT 67.520000 42.520000 67.720000 42.720000 ;
        RECT 67.520000 42.950000 67.720000 43.150000 ;
        RECT 67.520000 43.380000 67.720000 43.580000 ;
        RECT 67.520000 43.810000 67.720000 44.010000 ;
        RECT 67.520000 44.240000 67.720000 44.440000 ;
        RECT 67.520000 44.670000 67.720000 44.870000 ;
        RECT 67.520000 45.100000 67.720000 45.300000 ;
        RECT 67.520000 45.530000 67.720000 45.730000 ;
        RECT 67.520000 45.960000 67.720000 46.160000 ;
        RECT 67.925000 41.660000 68.125000 41.860000 ;
        RECT 67.925000 42.090000 68.125000 42.290000 ;
        RECT 67.925000 42.520000 68.125000 42.720000 ;
        RECT 67.925000 42.950000 68.125000 43.150000 ;
        RECT 67.925000 43.380000 68.125000 43.580000 ;
        RECT 67.925000 43.810000 68.125000 44.010000 ;
        RECT 67.925000 44.240000 68.125000 44.440000 ;
        RECT 67.925000 44.670000 68.125000 44.870000 ;
        RECT 67.925000 45.100000 68.125000 45.300000 ;
        RECT 67.925000 45.530000 68.125000 45.730000 ;
        RECT 67.925000 45.960000 68.125000 46.160000 ;
        RECT 68.330000 41.660000 68.530000 41.860000 ;
        RECT 68.330000 42.090000 68.530000 42.290000 ;
        RECT 68.330000 42.520000 68.530000 42.720000 ;
        RECT 68.330000 42.950000 68.530000 43.150000 ;
        RECT 68.330000 43.380000 68.530000 43.580000 ;
        RECT 68.330000 43.810000 68.530000 44.010000 ;
        RECT 68.330000 44.240000 68.530000 44.440000 ;
        RECT 68.330000 44.670000 68.530000 44.870000 ;
        RECT 68.330000 45.100000 68.530000 45.300000 ;
        RECT 68.330000 45.530000 68.530000 45.730000 ;
        RECT 68.330000 45.960000 68.530000 46.160000 ;
        RECT 68.735000 41.660000 68.935000 41.860000 ;
        RECT 68.735000 42.090000 68.935000 42.290000 ;
        RECT 68.735000 42.520000 68.935000 42.720000 ;
        RECT 68.735000 42.950000 68.935000 43.150000 ;
        RECT 68.735000 43.380000 68.935000 43.580000 ;
        RECT 68.735000 43.810000 68.935000 44.010000 ;
        RECT 68.735000 44.240000 68.935000 44.440000 ;
        RECT 68.735000 44.670000 68.935000 44.870000 ;
        RECT 68.735000 45.100000 68.935000 45.300000 ;
        RECT 68.735000 45.530000 68.935000 45.730000 ;
        RECT 68.735000 45.960000 68.935000 46.160000 ;
        RECT 69.140000 41.660000 69.340000 41.860000 ;
        RECT 69.140000 42.090000 69.340000 42.290000 ;
        RECT 69.140000 42.520000 69.340000 42.720000 ;
        RECT 69.140000 42.950000 69.340000 43.150000 ;
        RECT 69.140000 43.380000 69.340000 43.580000 ;
        RECT 69.140000 43.810000 69.340000 44.010000 ;
        RECT 69.140000 44.240000 69.340000 44.440000 ;
        RECT 69.140000 44.670000 69.340000 44.870000 ;
        RECT 69.140000 45.100000 69.340000 45.300000 ;
        RECT 69.140000 45.530000 69.340000 45.730000 ;
        RECT 69.140000 45.960000 69.340000 46.160000 ;
        RECT 69.545000 41.660000 69.745000 41.860000 ;
        RECT 69.545000 42.090000 69.745000 42.290000 ;
        RECT 69.545000 42.520000 69.745000 42.720000 ;
        RECT 69.545000 42.950000 69.745000 43.150000 ;
        RECT 69.545000 43.380000 69.745000 43.580000 ;
        RECT 69.545000 43.810000 69.745000 44.010000 ;
        RECT 69.545000 44.240000 69.745000 44.440000 ;
        RECT 69.545000 44.670000 69.745000 44.870000 ;
        RECT 69.545000 45.100000 69.745000 45.300000 ;
        RECT 69.545000 45.530000 69.745000 45.730000 ;
        RECT 69.545000 45.960000 69.745000 46.160000 ;
        RECT 69.950000 41.660000 70.150000 41.860000 ;
        RECT 69.950000 42.090000 70.150000 42.290000 ;
        RECT 69.950000 42.520000 70.150000 42.720000 ;
        RECT 69.950000 42.950000 70.150000 43.150000 ;
        RECT 69.950000 43.380000 70.150000 43.580000 ;
        RECT 69.950000 43.810000 70.150000 44.010000 ;
        RECT 69.950000 44.240000 70.150000 44.440000 ;
        RECT 69.950000 44.670000 70.150000 44.870000 ;
        RECT 69.950000 45.100000 70.150000 45.300000 ;
        RECT 69.950000 45.530000 70.150000 45.730000 ;
        RECT 69.950000 45.960000 70.150000 46.160000 ;
        RECT 70.355000 41.660000 70.555000 41.860000 ;
        RECT 70.355000 42.090000 70.555000 42.290000 ;
        RECT 70.355000 42.520000 70.555000 42.720000 ;
        RECT 70.355000 42.950000 70.555000 43.150000 ;
        RECT 70.355000 43.380000 70.555000 43.580000 ;
        RECT 70.355000 43.810000 70.555000 44.010000 ;
        RECT 70.355000 44.240000 70.555000 44.440000 ;
        RECT 70.355000 44.670000 70.555000 44.870000 ;
        RECT 70.355000 45.100000 70.555000 45.300000 ;
        RECT 70.355000 45.530000 70.555000 45.730000 ;
        RECT 70.355000 45.960000 70.555000 46.160000 ;
        RECT 70.760000 41.660000 70.960000 41.860000 ;
        RECT 70.760000 42.090000 70.960000 42.290000 ;
        RECT 70.760000 42.520000 70.960000 42.720000 ;
        RECT 70.760000 42.950000 70.960000 43.150000 ;
        RECT 70.760000 43.380000 70.960000 43.580000 ;
        RECT 70.760000 43.810000 70.960000 44.010000 ;
        RECT 70.760000 44.240000 70.960000 44.440000 ;
        RECT 70.760000 44.670000 70.960000 44.870000 ;
        RECT 70.760000 45.100000 70.960000 45.300000 ;
        RECT 70.760000 45.530000 70.960000 45.730000 ;
        RECT 70.760000 45.960000 70.960000 46.160000 ;
        RECT 71.165000 41.660000 71.365000 41.860000 ;
        RECT 71.165000 42.090000 71.365000 42.290000 ;
        RECT 71.165000 42.520000 71.365000 42.720000 ;
        RECT 71.165000 42.950000 71.365000 43.150000 ;
        RECT 71.165000 43.380000 71.365000 43.580000 ;
        RECT 71.165000 43.810000 71.365000 44.010000 ;
        RECT 71.165000 44.240000 71.365000 44.440000 ;
        RECT 71.165000 44.670000 71.365000 44.870000 ;
        RECT 71.165000 45.100000 71.365000 45.300000 ;
        RECT 71.165000 45.530000 71.365000 45.730000 ;
        RECT 71.165000 45.960000 71.365000 46.160000 ;
        RECT 71.570000 41.660000 71.770000 41.860000 ;
        RECT 71.570000 42.090000 71.770000 42.290000 ;
        RECT 71.570000 42.520000 71.770000 42.720000 ;
        RECT 71.570000 42.950000 71.770000 43.150000 ;
        RECT 71.570000 43.380000 71.770000 43.580000 ;
        RECT 71.570000 43.810000 71.770000 44.010000 ;
        RECT 71.570000 44.240000 71.770000 44.440000 ;
        RECT 71.570000 44.670000 71.770000 44.870000 ;
        RECT 71.570000 45.100000 71.770000 45.300000 ;
        RECT 71.570000 45.530000 71.770000 45.730000 ;
        RECT 71.570000 45.960000 71.770000 46.160000 ;
        RECT 71.975000 41.660000 72.175000 41.860000 ;
        RECT 71.975000 42.090000 72.175000 42.290000 ;
        RECT 71.975000 42.520000 72.175000 42.720000 ;
        RECT 71.975000 42.950000 72.175000 43.150000 ;
        RECT 71.975000 43.380000 72.175000 43.580000 ;
        RECT 71.975000 43.810000 72.175000 44.010000 ;
        RECT 71.975000 44.240000 72.175000 44.440000 ;
        RECT 71.975000 44.670000 72.175000 44.870000 ;
        RECT 71.975000 45.100000 72.175000 45.300000 ;
        RECT 71.975000 45.530000 72.175000 45.730000 ;
        RECT 71.975000 45.960000 72.175000 46.160000 ;
        RECT 72.380000 41.660000 72.580000 41.860000 ;
        RECT 72.380000 42.090000 72.580000 42.290000 ;
        RECT 72.380000 42.520000 72.580000 42.720000 ;
        RECT 72.380000 42.950000 72.580000 43.150000 ;
        RECT 72.380000 43.380000 72.580000 43.580000 ;
        RECT 72.380000 43.810000 72.580000 44.010000 ;
        RECT 72.380000 44.240000 72.580000 44.440000 ;
        RECT 72.380000 44.670000 72.580000 44.870000 ;
        RECT 72.380000 45.100000 72.580000 45.300000 ;
        RECT 72.380000 45.530000 72.580000 45.730000 ;
        RECT 72.380000 45.960000 72.580000 46.160000 ;
        RECT 72.785000 41.660000 72.985000 41.860000 ;
        RECT 72.785000 42.090000 72.985000 42.290000 ;
        RECT 72.785000 42.520000 72.985000 42.720000 ;
        RECT 72.785000 42.950000 72.985000 43.150000 ;
        RECT 72.785000 43.380000 72.985000 43.580000 ;
        RECT 72.785000 43.810000 72.985000 44.010000 ;
        RECT 72.785000 44.240000 72.985000 44.440000 ;
        RECT 72.785000 44.670000 72.985000 44.870000 ;
        RECT 72.785000 45.100000 72.985000 45.300000 ;
        RECT 72.785000 45.530000 72.985000 45.730000 ;
        RECT 72.785000 45.960000 72.985000 46.160000 ;
        RECT 73.190000 41.660000 73.390000 41.860000 ;
        RECT 73.190000 42.090000 73.390000 42.290000 ;
        RECT 73.190000 42.520000 73.390000 42.720000 ;
        RECT 73.190000 42.950000 73.390000 43.150000 ;
        RECT 73.190000 43.380000 73.390000 43.580000 ;
        RECT 73.190000 43.810000 73.390000 44.010000 ;
        RECT 73.190000 44.240000 73.390000 44.440000 ;
        RECT 73.190000 44.670000 73.390000 44.870000 ;
        RECT 73.190000 45.100000 73.390000 45.300000 ;
        RECT 73.190000 45.530000 73.390000 45.730000 ;
        RECT 73.190000 45.960000 73.390000 46.160000 ;
        RECT 73.595000 41.660000 73.795000 41.860000 ;
        RECT 73.595000 42.090000 73.795000 42.290000 ;
        RECT 73.595000 42.520000 73.795000 42.720000 ;
        RECT 73.595000 42.950000 73.795000 43.150000 ;
        RECT 73.595000 43.380000 73.795000 43.580000 ;
        RECT 73.595000 43.810000 73.795000 44.010000 ;
        RECT 73.595000 44.240000 73.795000 44.440000 ;
        RECT 73.595000 44.670000 73.795000 44.870000 ;
        RECT 73.595000 45.100000 73.795000 45.300000 ;
        RECT 73.595000 45.530000 73.795000 45.730000 ;
        RECT 73.595000 45.960000 73.795000 46.160000 ;
        RECT 74.000000 41.660000 74.200000 41.860000 ;
        RECT 74.000000 42.090000 74.200000 42.290000 ;
        RECT 74.000000 42.520000 74.200000 42.720000 ;
        RECT 74.000000 42.950000 74.200000 43.150000 ;
        RECT 74.000000 43.380000 74.200000 43.580000 ;
        RECT 74.000000 43.810000 74.200000 44.010000 ;
        RECT 74.000000 44.240000 74.200000 44.440000 ;
        RECT 74.000000 44.670000 74.200000 44.870000 ;
        RECT 74.000000 45.100000 74.200000 45.300000 ;
        RECT 74.000000 45.530000 74.200000 45.730000 ;
        RECT 74.000000 45.960000 74.200000 46.160000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 75.000000  41.190000 ;
      RECT  0.000000 41.190000  0.570000  46.630000 ;
      RECT  0.000000 46.630000 75.000000 200.000000 ;
      RECT 24.795000 41.190000 49.990000  46.630000 ;
      RECT 74.690000 41.190000 75.000000  46.630000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000  19.385000 73.330000  41.185000 ;
      RECT  1.670000  46.635000 73.330000  95.400000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT 24.770000  41.185000 50.015000  46.635000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT 0.000000   0.000000 75.000000   1.335000 ;
      RECT 0.000000  95.785000 75.000000 174.985000 ;
      RECT 1.765000  14.235000 73.235000  19.085000 ;
      RECT 2.070000   1.335000 72.930000  14.235000 ;
      RECT 2.070000  19.085000 72.930000  95.785000 ;
      RECT 2.070000 174.985000 72.930000 200.000000 ;
  END
END sky130_fd_io__overlay_vssd_hvc


MACRO sky130_fd_io__overlay_vssa_hvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.495000 51.650000 24.395000 52.820000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 47.740000 24.395000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 56.410000 24.395000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.970000 36.740000 24.395000 40.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 36.740000 74.290000 40.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 47.740000 74.290000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 51.650000 74.290000 52.820000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 56.410000 74.290000 56.730000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 24.370000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 24.370000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 24.370000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 24.370000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.585000 51.715000  0.785000 51.915000 ;
        RECT  0.585000 52.135000  0.785000 52.335000 ;
        RECT  0.585000 52.555000  0.785000 52.755000 ;
        RECT  0.620000 47.800000  0.820000 48.000000 ;
        RECT  0.620000 56.470000  0.820000 56.670000 ;
        RECT  0.995000 51.715000  1.195000 51.915000 ;
        RECT  0.995000 52.135000  1.195000 52.335000 ;
        RECT  0.995000 52.555000  1.195000 52.755000 ;
        RECT  1.025000 47.800000  1.225000 48.000000 ;
        RECT  1.025000 56.470000  1.225000 56.670000 ;
        RECT  1.060000 36.820000  1.260000 37.020000 ;
        RECT  1.060000 37.260000  1.260000 37.460000 ;
        RECT  1.060000 37.700000  1.260000 37.900000 ;
        RECT  1.060000 38.140000  1.260000 38.340000 ;
        RECT  1.060000 38.580000  1.260000 38.780000 ;
        RECT  1.060000 39.020000  1.260000 39.220000 ;
        RECT  1.060000 39.460000  1.260000 39.660000 ;
        RECT  1.060000 39.900000  1.260000 40.100000 ;
        RECT  1.405000 51.715000  1.605000 51.915000 ;
        RECT  1.405000 52.135000  1.605000 52.335000 ;
        RECT  1.405000 52.555000  1.605000 52.755000 ;
        RECT  1.430000 47.800000  1.630000 48.000000 ;
        RECT  1.430000 56.470000  1.630000 56.670000 ;
        RECT  1.465000 36.820000  1.665000 37.020000 ;
        RECT  1.465000 37.260000  1.665000 37.460000 ;
        RECT  1.465000 37.700000  1.665000 37.900000 ;
        RECT  1.465000 38.140000  1.665000 38.340000 ;
        RECT  1.465000 38.580000  1.665000 38.780000 ;
        RECT  1.465000 39.020000  1.665000 39.220000 ;
        RECT  1.465000 39.460000  1.665000 39.660000 ;
        RECT  1.465000 39.900000  1.665000 40.100000 ;
        RECT  1.815000 51.715000  2.015000 51.915000 ;
        RECT  1.815000 52.135000  2.015000 52.335000 ;
        RECT  1.815000 52.555000  2.015000 52.755000 ;
        RECT  1.835000 47.800000  2.035000 48.000000 ;
        RECT  1.835000 56.470000  2.035000 56.670000 ;
        RECT  1.870000 36.820000  2.070000 37.020000 ;
        RECT  1.870000 37.260000  2.070000 37.460000 ;
        RECT  1.870000 37.700000  2.070000 37.900000 ;
        RECT  1.870000 38.140000  2.070000 38.340000 ;
        RECT  1.870000 38.580000  2.070000 38.780000 ;
        RECT  1.870000 39.020000  2.070000 39.220000 ;
        RECT  1.870000 39.460000  2.070000 39.660000 ;
        RECT  1.870000 39.900000  2.070000 40.100000 ;
        RECT  2.225000 51.715000  2.425000 51.915000 ;
        RECT  2.225000 52.135000  2.425000 52.335000 ;
        RECT  2.225000 52.555000  2.425000 52.755000 ;
        RECT  2.240000 47.800000  2.440000 48.000000 ;
        RECT  2.240000 56.470000  2.440000 56.670000 ;
        RECT  2.275000 36.820000  2.475000 37.020000 ;
        RECT  2.275000 37.260000  2.475000 37.460000 ;
        RECT  2.275000 37.700000  2.475000 37.900000 ;
        RECT  2.275000 38.140000  2.475000 38.340000 ;
        RECT  2.275000 38.580000  2.475000 38.780000 ;
        RECT  2.275000 39.020000  2.475000 39.220000 ;
        RECT  2.275000 39.460000  2.475000 39.660000 ;
        RECT  2.275000 39.900000  2.475000 40.100000 ;
        RECT  2.635000 51.715000  2.835000 51.915000 ;
        RECT  2.635000 52.135000  2.835000 52.335000 ;
        RECT  2.635000 52.555000  2.835000 52.755000 ;
        RECT  2.645000 47.800000  2.845000 48.000000 ;
        RECT  2.645000 56.470000  2.845000 56.670000 ;
        RECT  2.680000 36.820000  2.880000 37.020000 ;
        RECT  2.680000 37.260000  2.880000 37.460000 ;
        RECT  2.680000 37.700000  2.880000 37.900000 ;
        RECT  2.680000 38.140000  2.880000 38.340000 ;
        RECT  2.680000 38.580000  2.880000 38.780000 ;
        RECT  2.680000 39.020000  2.880000 39.220000 ;
        RECT  2.680000 39.460000  2.880000 39.660000 ;
        RECT  2.680000 39.900000  2.880000 40.100000 ;
        RECT  3.045000 51.715000  3.245000 51.915000 ;
        RECT  3.045000 52.135000  3.245000 52.335000 ;
        RECT  3.045000 52.555000  3.245000 52.755000 ;
        RECT  3.050000 47.800000  3.250000 48.000000 ;
        RECT  3.050000 56.470000  3.250000 56.670000 ;
        RECT  3.085000 36.820000  3.285000 37.020000 ;
        RECT  3.085000 37.260000  3.285000 37.460000 ;
        RECT  3.085000 37.700000  3.285000 37.900000 ;
        RECT  3.085000 38.140000  3.285000 38.340000 ;
        RECT  3.085000 38.580000  3.285000 38.780000 ;
        RECT  3.085000 39.020000  3.285000 39.220000 ;
        RECT  3.085000 39.460000  3.285000 39.660000 ;
        RECT  3.085000 39.900000  3.285000 40.100000 ;
        RECT  3.450000 51.715000  3.650000 51.915000 ;
        RECT  3.450000 52.135000  3.650000 52.335000 ;
        RECT  3.450000 52.555000  3.650000 52.755000 ;
        RECT  3.455000 47.800000  3.655000 48.000000 ;
        RECT  3.455000 56.470000  3.655000 56.670000 ;
        RECT  3.490000 36.820000  3.690000 37.020000 ;
        RECT  3.490000 37.260000  3.690000 37.460000 ;
        RECT  3.490000 37.700000  3.690000 37.900000 ;
        RECT  3.490000 38.140000  3.690000 38.340000 ;
        RECT  3.490000 38.580000  3.690000 38.780000 ;
        RECT  3.490000 39.020000  3.690000 39.220000 ;
        RECT  3.490000 39.460000  3.690000 39.660000 ;
        RECT  3.490000 39.900000  3.690000 40.100000 ;
        RECT  3.855000 51.715000  4.055000 51.915000 ;
        RECT  3.855000 52.135000  4.055000 52.335000 ;
        RECT  3.855000 52.555000  4.055000 52.755000 ;
        RECT  3.860000 47.800000  4.060000 48.000000 ;
        RECT  3.860000 56.470000  4.060000 56.670000 ;
        RECT  3.895000 36.820000  4.095000 37.020000 ;
        RECT  3.895000 37.260000  4.095000 37.460000 ;
        RECT  3.895000 37.700000  4.095000 37.900000 ;
        RECT  3.895000 38.140000  4.095000 38.340000 ;
        RECT  3.895000 38.580000  4.095000 38.780000 ;
        RECT  3.895000 39.020000  4.095000 39.220000 ;
        RECT  3.895000 39.460000  4.095000 39.660000 ;
        RECT  3.895000 39.900000  4.095000 40.100000 ;
        RECT  4.260000 51.715000  4.460000 51.915000 ;
        RECT  4.260000 52.135000  4.460000 52.335000 ;
        RECT  4.260000 52.555000  4.460000 52.755000 ;
        RECT  4.265000 47.800000  4.465000 48.000000 ;
        RECT  4.265000 56.470000  4.465000 56.670000 ;
        RECT  4.300000 36.820000  4.500000 37.020000 ;
        RECT  4.300000 37.260000  4.500000 37.460000 ;
        RECT  4.300000 37.700000  4.500000 37.900000 ;
        RECT  4.300000 38.140000  4.500000 38.340000 ;
        RECT  4.300000 38.580000  4.500000 38.780000 ;
        RECT  4.300000 39.020000  4.500000 39.220000 ;
        RECT  4.300000 39.460000  4.500000 39.660000 ;
        RECT  4.300000 39.900000  4.500000 40.100000 ;
        RECT  4.665000 51.715000  4.865000 51.915000 ;
        RECT  4.665000 52.135000  4.865000 52.335000 ;
        RECT  4.665000 52.555000  4.865000 52.755000 ;
        RECT  4.670000 47.800000  4.870000 48.000000 ;
        RECT  4.670000 56.470000  4.870000 56.670000 ;
        RECT  4.705000 36.820000  4.905000 37.020000 ;
        RECT  4.705000 37.260000  4.905000 37.460000 ;
        RECT  4.705000 37.700000  4.905000 37.900000 ;
        RECT  4.705000 38.140000  4.905000 38.340000 ;
        RECT  4.705000 38.580000  4.905000 38.780000 ;
        RECT  4.705000 39.020000  4.905000 39.220000 ;
        RECT  4.705000 39.460000  4.905000 39.660000 ;
        RECT  4.705000 39.900000  4.905000 40.100000 ;
        RECT  5.070000 51.715000  5.270000 51.915000 ;
        RECT  5.070000 52.135000  5.270000 52.335000 ;
        RECT  5.070000 52.555000  5.270000 52.755000 ;
        RECT  5.075000 47.800000  5.275000 48.000000 ;
        RECT  5.075000 56.470000  5.275000 56.670000 ;
        RECT  5.110000 36.820000  5.310000 37.020000 ;
        RECT  5.110000 37.260000  5.310000 37.460000 ;
        RECT  5.110000 37.700000  5.310000 37.900000 ;
        RECT  5.110000 38.140000  5.310000 38.340000 ;
        RECT  5.110000 38.580000  5.310000 38.780000 ;
        RECT  5.110000 39.020000  5.310000 39.220000 ;
        RECT  5.110000 39.460000  5.310000 39.660000 ;
        RECT  5.110000 39.900000  5.310000 40.100000 ;
        RECT  5.475000 51.715000  5.675000 51.915000 ;
        RECT  5.475000 52.135000  5.675000 52.335000 ;
        RECT  5.475000 52.555000  5.675000 52.755000 ;
        RECT  5.480000 47.800000  5.680000 48.000000 ;
        RECT  5.480000 56.470000  5.680000 56.670000 ;
        RECT  5.515000 36.820000  5.715000 37.020000 ;
        RECT  5.515000 37.260000  5.715000 37.460000 ;
        RECT  5.515000 37.700000  5.715000 37.900000 ;
        RECT  5.515000 38.140000  5.715000 38.340000 ;
        RECT  5.515000 38.580000  5.715000 38.780000 ;
        RECT  5.515000 39.020000  5.715000 39.220000 ;
        RECT  5.515000 39.460000  5.715000 39.660000 ;
        RECT  5.515000 39.900000  5.715000 40.100000 ;
        RECT  5.880000 51.715000  6.080000 51.915000 ;
        RECT  5.880000 52.135000  6.080000 52.335000 ;
        RECT  5.880000 52.555000  6.080000 52.755000 ;
        RECT  5.885000 47.800000  6.085000 48.000000 ;
        RECT  5.885000 56.470000  6.085000 56.670000 ;
        RECT  5.920000 36.820000  6.120000 37.020000 ;
        RECT  5.920000 37.260000  6.120000 37.460000 ;
        RECT  5.920000 37.700000  6.120000 37.900000 ;
        RECT  5.920000 38.140000  6.120000 38.340000 ;
        RECT  5.920000 38.580000  6.120000 38.780000 ;
        RECT  5.920000 39.020000  6.120000 39.220000 ;
        RECT  5.920000 39.460000  6.120000 39.660000 ;
        RECT  5.920000 39.900000  6.120000 40.100000 ;
        RECT  6.285000 51.715000  6.485000 51.915000 ;
        RECT  6.285000 52.135000  6.485000 52.335000 ;
        RECT  6.285000 52.555000  6.485000 52.755000 ;
        RECT  6.290000 47.800000  6.490000 48.000000 ;
        RECT  6.290000 56.470000  6.490000 56.670000 ;
        RECT  6.325000 36.820000  6.525000 37.020000 ;
        RECT  6.325000 37.260000  6.525000 37.460000 ;
        RECT  6.325000 37.700000  6.525000 37.900000 ;
        RECT  6.325000 38.140000  6.525000 38.340000 ;
        RECT  6.325000 38.580000  6.525000 38.780000 ;
        RECT  6.325000 39.020000  6.525000 39.220000 ;
        RECT  6.325000 39.460000  6.525000 39.660000 ;
        RECT  6.325000 39.900000  6.525000 40.100000 ;
        RECT  6.690000 51.715000  6.890000 51.915000 ;
        RECT  6.690000 52.135000  6.890000 52.335000 ;
        RECT  6.690000 52.555000  6.890000 52.755000 ;
        RECT  6.695000 47.800000  6.895000 48.000000 ;
        RECT  6.695000 56.470000  6.895000 56.670000 ;
        RECT  6.730000 36.820000  6.930000 37.020000 ;
        RECT  6.730000 37.260000  6.930000 37.460000 ;
        RECT  6.730000 37.700000  6.930000 37.900000 ;
        RECT  6.730000 38.140000  6.930000 38.340000 ;
        RECT  6.730000 38.580000  6.930000 38.780000 ;
        RECT  6.730000 39.020000  6.930000 39.220000 ;
        RECT  6.730000 39.460000  6.930000 39.660000 ;
        RECT  6.730000 39.900000  6.930000 40.100000 ;
        RECT  7.095000 51.715000  7.295000 51.915000 ;
        RECT  7.095000 52.135000  7.295000 52.335000 ;
        RECT  7.095000 52.555000  7.295000 52.755000 ;
        RECT  7.100000 47.800000  7.300000 48.000000 ;
        RECT  7.100000 56.470000  7.300000 56.670000 ;
        RECT  7.135000 36.820000  7.335000 37.020000 ;
        RECT  7.135000 37.260000  7.335000 37.460000 ;
        RECT  7.135000 37.700000  7.335000 37.900000 ;
        RECT  7.135000 38.140000  7.335000 38.340000 ;
        RECT  7.135000 38.580000  7.335000 38.780000 ;
        RECT  7.135000 39.020000  7.335000 39.220000 ;
        RECT  7.135000 39.460000  7.335000 39.660000 ;
        RECT  7.135000 39.900000  7.335000 40.100000 ;
        RECT  7.500000 51.715000  7.700000 51.915000 ;
        RECT  7.500000 52.135000  7.700000 52.335000 ;
        RECT  7.500000 52.555000  7.700000 52.755000 ;
        RECT  7.505000 47.800000  7.705000 48.000000 ;
        RECT  7.505000 56.470000  7.705000 56.670000 ;
        RECT  7.540000 36.820000  7.740000 37.020000 ;
        RECT  7.540000 37.260000  7.740000 37.460000 ;
        RECT  7.540000 37.700000  7.740000 37.900000 ;
        RECT  7.540000 38.140000  7.740000 38.340000 ;
        RECT  7.540000 38.580000  7.740000 38.780000 ;
        RECT  7.540000 39.020000  7.740000 39.220000 ;
        RECT  7.540000 39.460000  7.740000 39.660000 ;
        RECT  7.540000 39.900000  7.740000 40.100000 ;
        RECT  7.905000 51.715000  8.105000 51.915000 ;
        RECT  7.905000 52.135000  8.105000 52.335000 ;
        RECT  7.905000 52.555000  8.105000 52.755000 ;
        RECT  7.910000 47.800000  8.110000 48.000000 ;
        RECT  7.910000 56.470000  8.110000 56.670000 ;
        RECT  7.945000 36.820000  8.145000 37.020000 ;
        RECT  7.945000 37.260000  8.145000 37.460000 ;
        RECT  7.945000 37.700000  8.145000 37.900000 ;
        RECT  7.945000 38.140000  8.145000 38.340000 ;
        RECT  7.945000 38.580000  8.145000 38.780000 ;
        RECT  7.945000 39.020000  8.145000 39.220000 ;
        RECT  7.945000 39.460000  8.145000 39.660000 ;
        RECT  7.945000 39.900000  8.145000 40.100000 ;
        RECT  8.310000 51.715000  8.510000 51.915000 ;
        RECT  8.310000 52.135000  8.510000 52.335000 ;
        RECT  8.310000 52.555000  8.510000 52.755000 ;
        RECT  8.315000 47.800000  8.515000 48.000000 ;
        RECT  8.315000 56.470000  8.515000 56.670000 ;
        RECT  8.350000 36.820000  8.550000 37.020000 ;
        RECT  8.350000 37.260000  8.550000 37.460000 ;
        RECT  8.350000 37.700000  8.550000 37.900000 ;
        RECT  8.350000 38.140000  8.550000 38.340000 ;
        RECT  8.350000 38.580000  8.550000 38.780000 ;
        RECT  8.350000 39.020000  8.550000 39.220000 ;
        RECT  8.350000 39.460000  8.550000 39.660000 ;
        RECT  8.350000 39.900000  8.550000 40.100000 ;
        RECT  8.715000 51.715000  8.915000 51.915000 ;
        RECT  8.715000 52.135000  8.915000 52.335000 ;
        RECT  8.715000 52.555000  8.915000 52.755000 ;
        RECT  8.720000 47.800000  8.920000 48.000000 ;
        RECT  8.720000 56.470000  8.920000 56.670000 ;
        RECT  8.755000 36.820000  8.955000 37.020000 ;
        RECT  8.755000 37.260000  8.955000 37.460000 ;
        RECT  8.755000 37.700000  8.955000 37.900000 ;
        RECT  8.755000 38.140000  8.955000 38.340000 ;
        RECT  8.755000 38.580000  8.955000 38.780000 ;
        RECT  8.755000 39.020000  8.955000 39.220000 ;
        RECT  8.755000 39.460000  8.955000 39.660000 ;
        RECT  8.755000 39.900000  8.955000 40.100000 ;
        RECT  9.120000 51.715000  9.320000 51.915000 ;
        RECT  9.120000 52.135000  9.320000 52.335000 ;
        RECT  9.120000 52.555000  9.320000 52.755000 ;
        RECT  9.125000 47.800000  9.325000 48.000000 ;
        RECT  9.125000 56.470000  9.325000 56.670000 ;
        RECT  9.160000 36.820000  9.360000 37.020000 ;
        RECT  9.160000 37.260000  9.360000 37.460000 ;
        RECT  9.160000 37.700000  9.360000 37.900000 ;
        RECT  9.160000 38.140000  9.360000 38.340000 ;
        RECT  9.160000 38.580000  9.360000 38.780000 ;
        RECT  9.160000 39.020000  9.360000 39.220000 ;
        RECT  9.160000 39.460000  9.360000 39.660000 ;
        RECT  9.160000 39.900000  9.360000 40.100000 ;
        RECT  9.525000 51.715000  9.725000 51.915000 ;
        RECT  9.525000 52.135000  9.725000 52.335000 ;
        RECT  9.525000 52.555000  9.725000 52.755000 ;
        RECT  9.530000 47.800000  9.730000 48.000000 ;
        RECT  9.530000 56.470000  9.730000 56.670000 ;
        RECT  9.565000 36.820000  9.765000 37.020000 ;
        RECT  9.565000 37.260000  9.765000 37.460000 ;
        RECT  9.565000 37.700000  9.765000 37.900000 ;
        RECT  9.565000 38.140000  9.765000 38.340000 ;
        RECT  9.565000 38.580000  9.765000 38.780000 ;
        RECT  9.565000 39.020000  9.765000 39.220000 ;
        RECT  9.565000 39.460000  9.765000 39.660000 ;
        RECT  9.565000 39.900000  9.765000 40.100000 ;
        RECT  9.930000 51.715000 10.130000 51.915000 ;
        RECT  9.930000 52.135000 10.130000 52.335000 ;
        RECT  9.930000 52.555000 10.130000 52.755000 ;
        RECT  9.935000 47.800000 10.135000 48.000000 ;
        RECT  9.935000 56.470000 10.135000 56.670000 ;
        RECT  9.970000 36.820000 10.170000 37.020000 ;
        RECT  9.970000 37.260000 10.170000 37.460000 ;
        RECT  9.970000 37.700000 10.170000 37.900000 ;
        RECT  9.970000 38.140000 10.170000 38.340000 ;
        RECT  9.970000 38.580000 10.170000 38.780000 ;
        RECT  9.970000 39.020000 10.170000 39.220000 ;
        RECT  9.970000 39.460000 10.170000 39.660000 ;
        RECT  9.970000 39.900000 10.170000 40.100000 ;
        RECT 10.335000 51.715000 10.535000 51.915000 ;
        RECT 10.335000 52.135000 10.535000 52.335000 ;
        RECT 10.335000 52.555000 10.535000 52.755000 ;
        RECT 10.340000 47.800000 10.540000 48.000000 ;
        RECT 10.340000 56.470000 10.540000 56.670000 ;
        RECT 10.375000 36.820000 10.575000 37.020000 ;
        RECT 10.375000 37.260000 10.575000 37.460000 ;
        RECT 10.375000 37.700000 10.575000 37.900000 ;
        RECT 10.375000 38.140000 10.575000 38.340000 ;
        RECT 10.375000 38.580000 10.575000 38.780000 ;
        RECT 10.375000 39.020000 10.575000 39.220000 ;
        RECT 10.375000 39.460000 10.575000 39.660000 ;
        RECT 10.375000 39.900000 10.575000 40.100000 ;
        RECT 10.740000 51.715000 10.940000 51.915000 ;
        RECT 10.740000 52.135000 10.940000 52.335000 ;
        RECT 10.740000 52.555000 10.940000 52.755000 ;
        RECT 10.745000 47.800000 10.945000 48.000000 ;
        RECT 10.745000 56.470000 10.945000 56.670000 ;
        RECT 10.780000 36.820000 10.980000 37.020000 ;
        RECT 10.780000 37.260000 10.980000 37.460000 ;
        RECT 10.780000 37.700000 10.980000 37.900000 ;
        RECT 10.780000 38.140000 10.980000 38.340000 ;
        RECT 10.780000 38.580000 10.980000 38.780000 ;
        RECT 10.780000 39.020000 10.980000 39.220000 ;
        RECT 10.780000 39.460000 10.980000 39.660000 ;
        RECT 10.780000 39.900000 10.980000 40.100000 ;
        RECT 11.145000 51.715000 11.345000 51.915000 ;
        RECT 11.145000 52.135000 11.345000 52.335000 ;
        RECT 11.145000 52.555000 11.345000 52.755000 ;
        RECT 11.150000 47.800000 11.350000 48.000000 ;
        RECT 11.150000 56.470000 11.350000 56.670000 ;
        RECT 11.185000 36.820000 11.385000 37.020000 ;
        RECT 11.185000 37.260000 11.385000 37.460000 ;
        RECT 11.185000 37.700000 11.385000 37.900000 ;
        RECT 11.185000 38.140000 11.385000 38.340000 ;
        RECT 11.185000 38.580000 11.385000 38.780000 ;
        RECT 11.185000 39.020000 11.385000 39.220000 ;
        RECT 11.185000 39.460000 11.385000 39.660000 ;
        RECT 11.185000 39.900000 11.385000 40.100000 ;
        RECT 11.550000 51.715000 11.750000 51.915000 ;
        RECT 11.550000 52.135000 11.750000 52.335000 ;
        RECT 11.550000 52.555000 11.750000 52.755000 ;
        RECT 11.555000 47.800000 11.755000 48.000000 ;
        RECT 11.555000 56.470000 11.755000 56.670000 ;
        RECT 11.590000 36.820000 11.790000 37.020000 ;
        RECT 11.590000 37.260000 11.790000 37.460000 ;
        RECT 11.590000 37.700000 11.790000 37.900000 ;
        RECT 11.590000 38.140000 11.790000 38.340000 ;
        RECT 11.590000 38.580000 11.790000 38.780000 ;
        RECT 11.590000 39.020000 11.790000 39.220000 ;
        RECT 11.590000 39.460000 11.790000 39.660000 ;
        RECT 11.590000 39.900000 11.790000 40.100000 ;
        RECT 11.955000 51.715000 12.155000 51.915000 ;
        RECT 11.955000 52.135000 12.155000 52.335000 ;
        RECT 11.955000 52.555000 12.155000 52.755000 ;
        RECT 11.960000 47.800000 12.160000 48.000000 ;
        RECT 11.960000 56.470000 12.160000 56.670000 ;
        RECT 11.995000 36.820000 12.195000 37.020000 ;
        RECT 11.995000 37.260000 12.195000 37.460000 ;
        RECT 11.995000 37.700000 12.195000 37.900000 ;
        RECT 11.995000 38.140000 12.195000 38.340000 ;
        RECT 11.995000 38.580000 12.195000 38.780000 ;
        RECT 11.995000 39.020000 12.195000 39.220000 ;
        RECT 11.995000 39.460000 12.195000 39.660000 ;
        RECT 11.995000 39.900000 12.195000 40.100000 ;
        RECT 12.360000 51.715000 12.560000 51.915000 ;
        RECT 12.360000 52.135000 12.560000 52.335000 ;
        RECT 12.360000 52.555000 12.560000 52.755000 ;
        RECT 12.365000 47.800000 12.565000 48.000000 ;
        RECT 12.365000 56.470000 12.565000 56.670000 ;
        RECT 12.400000 36.820000 12.600000 37.020000 ;
        RECT 12.400000 37.260000 12.600000 37.460000 ;
        RECT 12.400000 37.700000 12.600000 37.900000 ;
        RECT 12.400000 38.140000 12.600000 38.340000 ;
        RECT 12.400000 38.580000 12.600000 38.780000 ;
        RECT 12.400000 39.020000 12.600000 39.220000 ;
        RECT 12.400000 39.460000 12.600000 39.660000 ;
        RECT 12.400000 39.900000 12.600000 40.100000 ;
        RECT 12.765000 51.715000 12.965000 51.915000 ;
        RECT 12.765000 52.135000 12.965000 52.335000 ;
        RECT 12.765000 52.555000 12.965000 52.755000 ;
        RECT 12.770000 47.800000 12.970000 48.000000 ;
        RECT 12.770000 56.470000 12.970000 56.670000 ;
        RECT 12.805000 36.820000 13.005000 37.020000 ;
        RECT 12.805000 37.260000 13.005000 37.460000 ;
        RECT 12.805000 37.700000 13.005000 37.900000 ;
        RECT 12.805000 38.140000 13.005000 38.340000 ;
        RECT 12.805000 38.580000 13.005000 38.780000 ;
        RECT 12.805000 39.020000 13.005000 39.220000 ;
        RECT 12.805000 39.460000 13.005000 39.660000 ;
        RECT 12.805000 39.900000 13.005000 40.100000 ;
        RECT 13.170000 51.715000 13.370000 51.915000 ;
        RECT 13.170000 52.135000 13.370000 52.335000 ;
        RECT 13.170000 52.555000 13.370000 52.755000 ;
        RECT 13.175000 47.800000 13.375000 48.000000 ;
        RECT 13.175000 56.470000 13.375000 56.670000 ;
        RECT 13.210000 36.820000 13.410000 37.020000 ;
        RECT 13.210000 37.260000 13.410000 37.460000 ;
        RECT 13.210000 37.700000 13.410000 37.900000 ;
        RECT 13.210000 38.140000 13.410000 38.340000 ;
        RECT 13.210000 38.580000 13.410000 38.780000 ;
        RECT 13.210000 39.020000 13.410000 39.220000 ;
        RECT 13.210000 39.460000 13.410000 39.660000 ;
        RECT 13.210000 39.900000 13.410000 40.100000 ;
        RECT 13.575000 51.715000 13.775000 51.915000 ;
        RECT 13.575000 52.135000 13.775000 52.335000 ;
        RECT 13.575000 52.555000 13.775000 52.755000 ;
        RECT 13.580000 47.800000 13.780000 48.000000 ;
        RECT 13.580000 56.470000 13.780000 56.670000 ;
        RECT 13.615000 36.820000 13.815000 37.020000 ;
        RECT 13.615000 37.260000 13.815000 37.460000 ;
        RECT 13.615000 37.700000 13.815000 37.900000 ;
        RECT 13.615000 38.140000 13.815000 38.340000 ;
        RECT 13.615000 38.580000 13.815000 38.780000 ;
        RECT 13.615000 39.020000 13.815000 39.220000 ;
        RECT 13.615000 39.460000 13.815000 39.660000 ;
        RECT 13.615000 39.900000 13.815000 40.100000 ;
        RECT 13.980000 51.715000 14.180000 51.915000 ;
        RECT 13.980000 52.135000 14.180000 52.335000 ;
        RECT 13.980000 52.555000 14.180000 52.755000 ;
        RECT 13.985000 47.800000 14.185000 48.000000 ;
        RECT 13.985000 56.470000 14.185000 56.670000 ;
        RECT 14.020000 36.820000 14.220000 37.020000 ;
        RECT 14.020000 37.260000 14.220000 37.460000 ;
        RECT 14.020000 37.700000 14.220000 37.900000 ;
        RECT 14.020000 38.140000 14.220000 38.340000 ;
        RECT 14.020000 38.580000 14.220000 38.780000 ;
        RECT 14.020000 39.020000 14.220000 39.220000 ;
        RECT 14.020000 39.460000 14.220000 39.660000 ;
        RECT 14.020000 39.900000 14.220000 40.100000 ;
        RECT 14.385000 51.715000 14.585000 51.915000 ;
        RECT 14.385000 52.135000 14.585000 52.335000 ;
        RECT 14.385000 52.555000 14.585000 52.755000 ;
        RECT 14.390000 47.800000 14.590000 48.000000 ;
        RECT 14.390000 56.470000 14.590000 56.670000 ;
        RECT 14.425000 36.820000 14.625000 37.020000 ;
        RECT 14.425000 37.260000 14.625000 37.460000 ;
        RECT 14.425000 37.700000 14.625000 37.900000 ;
        RECT 14.425000 38.140000 14.625000 38.340000 ;
        RECT 14.425000 38.580000 14.625000 38.780000 ;
        RECT 14.425000 39.020000 14.625000 39.220000 ;
        RECT 14.425000 39.460000 14.625000 39.660000 ;
        RECT 14.425000 39.900000 14.625000 40.100000 ;
        RECT 14.790000 51.715000 14.990000 51.915000 ;
        RECT 14.790000 52.135000 14.990000 52.335000 ;
        RECT 14.790000 52.555000 14.990000 52.755000 ;
        RECT 14.795000 47.800000 14.995000 48.000000 ;
        RECT 14.795000 56.470000 14.995000 56.670000 ;
        RECT 14.830000 36.820000 15.030000 37.020000 ;
        RECT 14.830000 37.260000 15.030000 37.460000 ;
        RECT 14.830000 37.700000 15.030000 37.900000 ;
        RECT 14.830000 38.140000 15.030000 38.340000 ;
        RECT 14.830000 38.580000 15.030000 38.780000 ;
        RECT 14.830000 39.020000 15.030000 39.220000 ;
        RECT 14.830000 39.460000 15.030000 39.660000 ;
        RECT 14.830000 39.900000 15.030000 40.100000 ;
        RECT 15.195000 51.715000 15.395000 51.915000 ;
        RECT 15.195000 52.135000 15.395000 52.335000 ;
        RECT 15.195000 52.555000 15.395000 52.755000 ;
        RECT 15.200000 47.800000 15.400000 48.000000 ;
        RECT 15.200000 56.470000 15.400000 56.670000 ;
        RECT 15.235000 36.820000 15.435000 37.020000 ;
        RECT 15.235000 37.260000 15.435000 37.460000 ;
        RECT 15.235000 37.700000 15.435000 37.900000 ;
        RECT 15.235000 38.140000 15.435000 38.340000 ;
        RECT 15.235000 38.580000 15.435000 38.780000 ;
        RECT 15.235000 39.020000 15.435000 39.220000 ;
        RECT 15.235000 39.460000 15.435000 39.660000 ;
        RECT 15.235000 39.900000 15.435000 40.100000 ;
        RECT 15.600000 51.715000 15.800000 51.915000 ;
        RECT 15.600000 52.135000 15.800000 52.335000 ;
        RECT 15.600000 52.555000 15.800000 52.755000 ;
        RECT 15.605000 47.800000 15.805000 48.000000 ;
        RECT 15.605000 56.470000 15.805000 56.670000 ;
        RECT 15.640000 36.820000 15.840000 37.020000 ;
        RECT 15.640000 37.260000 15.840000 37.460000 ;
        RECT 15.640000 37.700000 15.840000 37.900000 ;
        RECT 15.640000 38.140000 15.840000 38.340000 ;
        RECT 15.640000 38.580000 15.840000 38.780000 ;
        RECT 15.640000 39.020000 15.840000 39.220000 ;
        RECT 15.640000 39.460000 15.840000 39.660000 ;
        RECT 15.640000 39.900000 15.840000 40.100000 ;
        RECT 16.005000 51.715000 16.205000 51.915000 ;
        RECT 16.005000 52.135000 16.205000 52.335000 ;
        RECT 16.005000 52.555000 16.205000 52.755000 ;
        RECT 16.010000 47.800000 16.210000 48.000000 ;
        RECT 16.010000 56.470000 16.210000 56.670000 ;
        RECT 16.045000 36.820000 16.245000 37.020000 ;
        RECT 16.045000 37.260000 16.245000 37.460000 ;
        RECT 16.045000 37.700000 16.245000 37.900000 ;
        RECT 16.045000 38.140000 16.245000 38.340000 ;
        RECT 16.045000 38.580000 16.245000 38.780000 ;
        RECT 16.045000 39.020000 16.245000 39.220000 ;
        RECT 16.045000 39.460000 16.245000 39.660000 ;
        RECT 16.045000 39.900000 16.245000 40.100000 ;
        RECT 16.410000 51.715000 16.610000 51.915000 ;
        RECT 16.410000 52.135000 16.610000 52.335000 ;
        RECT 16.410000 52.555000 16.610000 52.755000 ;
        RECT 16.415000 47.800000 16.615000 48.000000 ;
        RECT 16.415000 56.470000 16.615000 56.670000 ;
        RECT 16.450000 36.820000 16.650000 37.020000 ;
        RECT 16.450000 37.260000 16.650000 37.460000 ;
        RECT 16.450000 37.700000 16.650000 37.900000 ;
        RECT 16.450000 38.140000 16.650000 38.340000 ;
        RECT 16.450000 38.580000 16.650000 38.780000 ;
        RECT 16.450000 39.020000 16.650000 39.220000 ;
        RECT 16.450000 39.460000 16.650000 39.660000 ;
        RECT 16.450000 39.900000 16.650000 40.100000 ;
        RECT 16.815000 51.715000 17.015000 51.915000 ;
        RECT 16.815000 52.135000 17.015000 52.335000 ;
        RECT 16.815000 52.555000 17.015000 52.755000 ;
        RECT 16.820000 47.800000 17.020000 48.000000 ;
        RECT 16.820000 56.470000 17.020000 56.670000 ;
        RECT 16.855000 36.820000 17.055000 37.020000 ;
        RECT 16.855000 37.260000 17.055000 37.460000 ;
        RECT 16.855000 37.700000 17.055000 37.900000 ;
        RECT 16.855000 38.140000 17.055000 38.340000 ;
        RECT 16.855000 38.580000 17.055000 38.780000 ;
        RECT 16.855000 39.020000 17.055000 39.220000 ;
        RECT 16.855000 39.460000 17.055000 39.660000 ;
        RECT 16.855000 39.900000 17.055000 40.100000 ;
        RECT 17.220000 51.715000 17.420000 51.915000 ;
        RECT 17.220000 52.135000 17.420000 52.335000 ;
        RECT 17.220000 52.555000 17.420000 52.755000 ;
        RECT 17.225000 47.800000 17.425000 48.000000 ;
        RECT 17.225000 56.470000 17.425000 56.670000 ;
        RECT 17.260000 36.820000 17.460000 37.020000 ;
        RECT 17.260000 37.260000 17.460000 37.460000 ;
        RECT 17.260000 37.700000 17.460000 37.900000 ;
        RECT 17.260000 38.140000 17.460000 38.340000 ;
        RECT 17.260000 38.580000 17.460000 38.780000 ;
        RECT 17.260000 39.020000 17.460000 39.220000 ;
        RECT 17.260000 39.460000 17.460000 39.660000 ;
        RECT 17.260000 39.900000 17.460000 40.100000 ;
        RECT 17.625000 51.715000 17.825000 51.915000 ;
        RECT 17.625000 52.135000 17.825000 52.335000 ;
        RECT 17.625000 52.555000 17.825000 52.755000 ;
        RECT 17.630000 47.800000 17.830000 48.000000 ;
        RECT 17.630000 56.470000 17.830000 56.670000 ;
        RECT 17.665000 36.820000 17.865000 37.020000 ;
        RECT 17.665000 37.260000 17.865000 37.460000 ;
        RECT 17.665000 37.700000 17.865000 37.900000 ;
        RECT 17.665000 38.140000 17.865000 38.340000 ;
        RECT 17.665000 38.580000 17.865000 38.780000 ;
        RECT 17.665000 39.020000 17.865000 39.220000 ;
        RECT 17.665000 39.460000 17.865000 39.660000 ;
        RECT 17.665000 39.900000 17.865000 40.100000 ;
        RECT 18.030000 51.715000 18.230000 51.915000 ;
        RECT 18.030000 52.135000 18.230000 52.335000 ;
        RECT 18.030000 52.555000 18.230000 52.755000 ;
        RECT 18.035000 47.800000 18.235000 48.000000 ;
        RECT 18.035000 56.470000 18.235000 56.670000 ;
        RECT 18.070000 36.820000 18.270000 37.020000 ;
        RECT 18.070000 37.260000 18.270000 37.460000 ;
        RECT 18.070000 37.700000 18.270000 37.900000 ;
        RECT 18.070000 38.140000 18.270000 38.340000 ;
        RECT 18.070000 38.580000 18.270000 38.780000 ;
        RECT 18.070000 39.020000 18.270000 39.220000 ;
        RECT 18.070000 39.460000 18.270000 39.660000 ;
        RECT 18.070000 39.900000 18.270000 40.100000 ;
        RECT 18.435000 51.715000 18.635000 51.915000 ;
        RECT 18.435000 52.135000 18.635000 52.335000 ;
        RECT 18.435000 52.555000 18.635000 52.755000 ;
        RECT 18.440000 47.800000 18.640000 48.000000 ;
        RECT 18.440000 56.470000 18.640000 56.670000 ;
        RECT 18.475000 36.820000 18.675000 37.020000 ;
        RECT 18.475000 37.260000 18.675000 37.460000 ;
        RECT 18.475000 37.700000 18.675000 37.900000 ;
        RECT 18.475000 38.140000 18.675000 38.340000 ;
        RECT 18.475000 38.580000 18.675000 38.780000 ;
        RECT 18.475000 39.020000 18.675000 39.220000 ;
        RECT 18.475000 39.460000 18.675000 39.660000 ;
        RECT 18.475000 39.900000 18.675000 40.100000 ;
        RECT 18.840000 51.715000 19.040000 51.915000 ;
        RECT 18.840000 52.135000 19.040000 52.335000 ;
        RECT 18.840000 52.555000 19.040000 52.755000 ;
        RECT 18.845000 47.800000 19.045000 48.000000 ;
        RECT 18.845000 56.470000 19.045000 56.670000 ;
        RECT 18.880000 36.820000 19.080000 37.020000 ;
        RECT 18.880000 37.260000 19.080000 37.460000 ;
        RECT 18.880000 37.700000 19.080000 37.900000 ;
        RECT 18.880000 38.140000 19.080000 38.340000 ;
        RECT 18.880000 38.580000 19.080000 38.780000 ;
        RECT 18.880000 39.020000 19.080000 39.220000 ;
        RECT 18.880000 39.460000 19.080000 39.660000 ;
        RECT 18.880000 39.900000 19.080000 40.100000 ;
        RECT 19.245000 51.715000 19.445000 51.915000 ;
        RECT 19.245000 52.135000 19.445000 52.335000 ;
        RECT 19.245000 52.555000 19.445000 52.755000 ;
        RECT 19.250000 47.800000 19.450000 48.000000 ;
        RECT 19.250000 56.470000 19.450000 56.670000 ;
        RECT 19.285000 36.820000 19.485000 37.020000 ;
        RECT 19.285000 37.260000 19.485000 37.460000 ;
        RECT 19.285000 37.700000 19.485000 37.900000 ;
        RECT 19.285000 38.140000 19.485000 38.340000 ;
        RECT 19.285000 38.580000 19.485000 38.780000 ;
        RECT 19.285000 39.020000 19.485000 39.220000 ;
        RECT 19.285000 39.460000 19.485000 39.660000 ;
        RECT 19.285000 39.900000 19.485000 40.100000 ;
        RECT 19.650000 51.715000 19.850000 51.915000 ;
        RECT 19.650000 52.135000 19.850000 52.335000 ;
        RECT 19.650000 52.555000 19.850000 52.755000 ;
        RECT 19.655000 47.800000 19.855000 48.000000 ;
        RECT 19.655000 56.470000 19.855000 56.670000 ;
        RECT 19.690000 36.820000 19.890000 37.020000 ;
        RECT 19.690000 37.260000 19.890000 37.460000 ;
        RECT 19.690000 37.700000 19.890000 37.900000 ;
        RECT 19.690000 38.140000 19.890000 38.340000 ;
        RECT 19.690000 38.580000 19.890000 38.780000 ;
        RECT 19.690000 39.020000 19.890000 39.220000 ;
        RECT 19.690000 39.460000 19.890000 39.660000 ;
        RECT 19.690000 39.900000 19.890000 40.100000 ;
        RECT 20.055000 51.715000 20.255000 51.915000 ;
        RECT 20.055000 52.135000 20.255000 52.335000 ;
        RECT 20.055000 52.555000 20.255000 52.755000 ;
        RECT 20.060000 47.800000 20.260000 48.000000 ;
        RECT 20.060000 56.470000 20.260000 56.670000 ;
        RECT 20.095000 36.820000 20.295000 37.020000 ;
        RECT 20.095000 37.260000 20.295000 37.460000 ;
        RECT 20.095000 37.700000 20.295000 37.900000 ;
        RECT 20.095000 38.140000 20.295000 38.340000 ;
        RECT 20.095000 38.580000 20.295000 38.780000 ;
        RECT 20.095000 39.020000 20.295000 39.220000 ;
        RECT 20.095000 39.460000 20.295000 39.660000 ;
        RECT 20.095000 39.900000 20.295000 40.100000 ;
        RECT 20.460000 51.715000 20.660000 51.915000 ;
        RECT 20.460000 52.135000 20.660000 52.335000 ;
        RECT 20.460000 52.555000 20.660000 52.755000 ;
        RECT 20.465000 47.800000 20.665000 48.000000 ;
        RECT 20.465000 56.470000 20.665000 56.670000 ;
        RECT 20.500000 36.820000 20.700000 37.020000 ;
        RECT 20.500000 37.260000 20.700000 37.460000 ;
        RECT 20.500000 37.700000 20.700000 37.900000 ;
        RECT 20.500000 38.140000 20.700000 38.340000 ;
        RECT 20.500000 38.580000 20.700000 38.780000 ;
        RECT 20.500000 39.020000 20.700000 39.220000 ;
        RECT 20.500000 39.460000 20.700000 39.660000 ;
        RECT 20.500000 39.900000 20.700000 40.100000 ;
        RECT 20.865000 51.715000 21.065000 51.915000 ;
        RECT 20.865000 52.135000 21.065000 52.335000 ;
        RECT 20.865000 52.555000 21.065000 52.755000 ;
        RECT 20.870000 47.800000 21.070000 48.000000 ;
        RECT 20.870000 56.470000 21.070000 56.670000 ;
        RECT 20.905000 36.820000 21.105000 37.020000 ;
        RECT 20.905000 37.260000 21.105000 37.460000 ;
        RECT 20.905000 37.700000 21.105000 37.900000 ;
        RECT 20.905000 38.140000 21.105000 38.340000 ;
        RECT 20.905000 38.580000 21.105000 38.780000 ;
        RECT 20.905000 39.020000 21.105000 39.220000 ;
        RECT 20.905000 39.460000 21.105000 39.660000 ;
        RECT 20.905000 39.900000 21.105000 40.100000 ;
        RECT 21.270000 51.715000 21.470000 51.915000 ;
        RECT 21.270000 52.135000 21.470000 52.335000 ;
        RECT 21.270000 52.555000 21.470000 52.755000 ;
        RECT 21.275000 47.800000 21.475000 48.000000 ;
        RECT 21.275000 56.470000 21.475000 56.670000 ;
        RECT 21.305000 36.820000 21.505000 37.020000 ;
        RECT 21.305000 37.260000 21.505000 37.460000 ;
        RECT 21.305000 37.700000 21.505000 37.900000 ;
        RECT 21.305000 38.140000 21.505000 38.340000 ;
        RECT 21.305000 38.580000 21.505000 38.780000 ;
        RECT 21.305000 39.020000 21.505000 39.220000 ;
        RECT 21.305000 39.460000 21.505000 39.660000 ;
        RECT 21.305000 39.900000 21.505000 40.100000 ;
        RECT 21.675000 51.715000 21.875000 51.915000 ;
        RECT 21.675000 52.135000 21.875000 52.335000 ;
        RECT 21.675000 52.555000 21.875000 52.755000 ;
        RECT 21.680000 47.800000 21.880000 48.000000 ;
        RECT 21.680000 56.470000 21.880000 56.670000 ;
        RECT 21.705000 36.820000 21.905000 37.020000 ;
        RECT 21.705000 37.260000 21.905000 37.460000 ;
        RECT 21.705000 37.700000 21.905000 37.900000 ;
        RECT 21.705000 38.140000 21.905000 38.340000 ;
        RECT 21.705000 38.580000 21.905000 38.780000 ;
        RECT 21.705000 39.020000 21.905000 39.220000 ;
        RECT 21.705000 39.460000 21.905000 39.660000 ;
        RECT 21.705000 39.900000 21.905000 40.100000 ;
        RECT 22.080000 51.715000 22.280000 51.915000 ;
        RECT 22.080000 52.135000 22.280000 52.335000 ;
        RECT 22.080000 52.555000 22.280000 52.755000 ;
        RECT 22.085000 47.800000 22.285000 48.000000 ;
        RECT 22.085000 56.470000 22.285000 56.670000 ;
        RECT 22.105000 36.820000 22.305000 37.020000 ;
        RECT 22.105000 37.260000 22.305000 37.460000 ;
        RECT 22.105000 37.700000 22.305000 37.900000 ;
        RECT 22.105000 38.140000 22.305000 38.340000 ;
        RECT 22.105000 38.580000 22.305000 38.780000 ;
        RECT 22.105000 39.020000 22.305000 39.220000 ;
        RECT 22.105000 39.460000 22.305000 39.660000 ;
        RECT 22.105000 39.900000 22.305000 40.100000 ;
        RECT 22.485000 51.715000 22.685000 51.915000 ;
        RECT 22.485000 52.135000 22.685000 52.335000 ;
        RECT 22.485000 52.555000 22.685000 52.755000 ;
        RECT 22.490000 47.800000 22.690000 48.000000 ;
        RECT 22.490000 56.470000 22.690000 56.670000 ;
        RECT 22.505000 36.820000 22.705000 37.020000 ;
        RECT 22.505000 37.260000 22.705000 37.460000 ;
        RECT 22.505000 37.700000 22.705000 37.900000 ;
        RECT 22.505000 38.140000 22.705000 38.340000 ;
        RECT 22.505000 38.580000 22.705000 38.780000 ;
        RECT 22.505000 39.020000 22.705000 39.220000 ;
        RECT 22.505000 39.460000 22.705000 39.660000 ;
        RECT 22.505000 39.900000 22.705000 40.100000 ;
        RECT 22.890000 51.715000 23.090000 51.915000 ;
        RECT 22.890000 52.135000 23.090000 52.335000 ;
        RECT 22.890000 52.555000 23.090000 52.755000 ;
        RECT 22.895000 47.800000 23.095000 48.000000 ;
        RECT 22.895000 56.470000 23.095000 56.670000 ;
        RECT 22.905000 36.820000 23.105000 37.020000 ;
        RECT 22.905000 37.260000 23.105000 37.460000 ;
        RECT 22.905000 37.700000 23.105000 37.900000 ;
        RECT 22.905000 38.140000 23.105000 38.340000 ;
        RECT 22.905000 38.580000 23.105000 38.780000 ;
        RECT 22.905000 39.020000 23.105000 39.220000 ;
        RECT 22.905000 39.460000 23.105000 39.660000 ;
        RECT 22.905000 39.900000 23.105000 40.100000 ;
        RECT 23.295000 51.715000 23.495000 51.915000 ;
        RECT 23.295000 52.135000 23.495000 52.335000 ;
        RECT 23.295000 52.555000 23.495000 52.755000 ;
        RECT 23.300000 47.800000 23.500000 48.000000 ;
        RECT 23.300000 56.470000 23.500000 56.670000 ;
        RECT 23.305000 36.820000 23.505000 37.020000 ;
        RECT 23.305000 37.260000 23.505000 37.460000 ;
        RECT 23.305000 37.700000 23.505000 37.900000 ;
        RECT 23.305000 38.140000 23.505000 38.340000 ;
        RECT 23.305000 38.580000 23.505000 38.780000 ;
        RECT 23.305000 39.020000 23.505000 39.220000 ;
        RECT 23.305000 39.460000 23.505000 39.660000 ;
        RECT 23.305000 39.900000 23.505000 40.100000 ;
        RECT 23.700000 51.715000 23.900000 51.915000 ;
        RECT 23.700000 52.135000 23.900000 52.335000 ;
        RECT 23.700000 52.555000 23.900000 52.755000 ;
        RECT 23.705000 36.820000 23.905000 37.020000 ;
        RECT 23.705000 37.260000 23.905000 37.460000 ;
        RECT 23.705000 37.700000 23.905000 37.900000 ;
        RECT 23.705000 38.140000 23.905000 38.340000 ;
        RECT 23.705000 38.580000 23.905000 38.780000 ;
        RECT 23.705000 39.020000 23.905000 39.220000 ;
        RECT 23.705000 39.460000 23.905000 39.660000 ;
        RECT 23.705000 39.900000 23.905000 40.100000 ;
        RECT 23.705000 47.800000 23.905000 48.000000 ;
        RECT 23.705000 56.470000 23.905000 56.670000 ;
        RECT 24.105000 36.820000 24.305000 37.020000 ;
        RECT 24.105000 37.260000 24.305000 37.460000 ;
        RECT 24.105000 37.700000 24.305000 37.900000 ;
        RECT 24.105000 38.140000 24.305000 38.340000 ;
        RECT 24.105000 38.580000 24.305000 38.780000 ;
        RECT 24.105000 39.020000 24.305000 39.220000 ;
        RECT 24.105000 39.460000 24.305000 39.660000 ;
        RECT 24.105000 39.900000 24.305000 40.100000 ;
        RECT 24.105000 47.800000 24.305000 48.000000 ;
        RECT 24.105000 51.715000 24.305000 51.915000 ;
        RECT 24.105000 52.135000 24.305000 52.335000 ;
        RECT 24.105000 52.555000 24.305000 52.755000 ;
        RECT 24.105000 56.470000 24.305000 56.670000 ;
        RECT 50.480000 36.820000 50.680000 37.020000 ;
        RECT 50.480000 37.260000 50.680000 37.460000 ;
        RECT 50.480000 37.700000 50.680000 37.900000 ;
        RECT 50.480000 38.140000 50.680000 38.340000 ;
        RECT 50.480000 38.580000 50.680000 38.780000 ;
        RECT 50.480000 39.020000 50.680000 39.220000 ;
        RECT 50.480000 39.460000 50.680000 39.660000 ;
        RECT 50.480000 39.900000 50.680000 40.100000 ;
        RECT 50.480000 47.800000 50.680000 48.000000 ;
        RECT 50.480000 51.715000 50.680000 51.915000 ;
        RECT 50.480000 52.135000 50.680000 52.335000 ;
        RECT 50.480000 52.555000 50.680000 52.755000 ;
        RECT 50.480000 56.470000 50.680000 56.670000 ;
        RECT 50.885000 47.800000 51.085000 48.000000 ;
        RECT 50.885000 56.470000 51.085000 56.670000 ;
        RECT 50.890000 36.820000 51.090000 37.020000 ;
        RECT 50.890000 37.260000 51.090000 37.460000 ;
        RECT 50.890000 37.700000 51.090000 37.900000 ;
        RECT 50.890000 38.140000 51.090000 38.340000 ;
        RECT 50.890000 38.580000 51.090000 38.780000 ;
        RECT 50.890000 39.020000 51.090000 39.220000 ;
        RECT 50.890000 39.460000 51.090000 39.660000 ;
        RECT 50.890000 39.900000 51.090000 40.100000 ;
        RECT 50.890000 51.715000 51.090000 51.915000 ;
        RECT 50.890000 52.135000 51.090000 52.335000 ;
        RECT 50.890000 52.555000 51.090000 52.755000 ;
        RECT 51.290000 47.800000 51.490000 48.000000 ;
        RECT 51.290000 56.470000 51.490000 56.670000 ;
        RECT 51.300000 36.820000 51.500000 37.020000 ;
        RECT 51.300000 37.260000 51.500000 37.460000 ;
        RECT 51.300000 37.700000 51.500000 37.900000 ;
        RECT 51.300000 38.140000 51.500000 38.340000 ;
        RECT 51.300000 38.580000 51.500000 38.780000 ;
        RECT 51.300000 39.020000 51.500000 39.220000 ;
        RECT 51.300000 39.460000 51.500000 39.660000 ;
        RECT 51.300000 39.900000 51.500000 40.100000 ;
        RECT 51.300000 51.715000 51.500000 51.915000 ;
        RECT 51.300000 52.135000 51.500000 52.335000 ;
        RECT 51.300000 52.555000 51.500000 52.755000 ;
        RECT 51.695000 47.800000 51.895000 48.000000 ;
        RECT 51.695000 56.470000 51.895000 56.670000 ;
        RECT 51.710000 36.820000 51.910000 37.020000 ;
        RECT 51.710000 37.260000 51.910000 37.460000 ;
        RECT 51.710000 37.700000 51.910000 37.900000 ;
        RECT 51.710000 38.140000 51.910000 38.340000 ;
        RECT 51.710000 38.580000 51.910000 38.780000 ;
        RECT 51.710000 39.020000 51.910000 39.220000 ;
        RECT 51.710000 39.460000 51.910000 39.660000 ;
        RECT 51.710000 39.900000 51.910000 40.100000 ;
        RECT 51.710000 51.715000 51.910000 51.915000 ;
        RECT 51.710000 52.135000 51.910000 52.335000 ;
        RECT 51.710000 52.555000 51.910000 52.755000 ;
        RECT 52.100000 47.800000 52.300000 48.000000 ;
        RECT 52.100000 56.470000 52.300000 56.670000 ;
        RECT 52.120000 36.820000 52.320000 37.020000 ;
        RECT 52.120000 37.260000 52.320000 37.460000 ;
        RECT 52.120000 37.700000 52.320000 37.900000 ;
        RECT 52.120000 38.140000 52.320000 38.340000 ;
        RECT 52.120000 38.580000 52.320000 38.780000 ;
        RECT 52.120000 39.020000 52.320000 39.220000 ;
        RECT 52.120000 39.460000 52.320000 39.660000 ;
        RECT 52.120000 39.900000 52.320000 40.100000 ;
        RECT 52.120000 51.715000 52.320000 51.915000 ;
        RECT 52.120000 52.135000 52.320000 52.335000 ;
        RECT 52.120000 52.555000 52.320000 52.755000 ;
        RECT 52.505000 47.800000 52.705000 48.000000 ;
        RECT 52.505000 56.470000 52.705000 56.670000 ;
        RECT 52.530000 36.820000 52.730000 37.020000 ;
        RECT 52.530000 37.260000 52.730000 37.460000 ;
        RECT 52.530000 37.700000 52.730000 37.900000 ;
        RECT 52.530000 38.140000 52.730000 38.340000 ;
        RECT 52.530000 38.580000 52.730000 38.780000 ;
        RECT 52.530000 39.020000 52.730000 39.220000 ;
        RECT 52.530000 39.460000 52.730000 39.660000 ;
        RECT 52.530000 39.900000 52.730000 40.100000 ;
        RECT 52.530000 51.715000 52.730000 51.915000 ;
        RECT 52.530000 52.135000 52.730000 52.335000 ;
        RECT 52.530000 52.555000 52.730000 52.755000 ;
        RECT 52.910000 47.800000 53.110000 48.000000 ;
        RECT 52.910000 56.470000 53.110000 56.670000 ;
        RECT 52.940000 36.820000 53.140000 37.020000 ;
        RECT 52.940000 37.260000 53.140000 37.460000 ;
        RECT 52.940000 37.700000 53.140000 37.900000 ;
        RECT 52.940000 38.140000 53.140000 38.340000 ;
        RECT 52.940000 38.580000 53.140000 38.780000 ;
        RECT 52.940000 39.020000 53.140000 39.220000 ;
        RECT 52.940000 39.460000 53.140000 39.660000 ;
        RECT 52.940000 39.900000 53.140000 40.100000 ;
        RECT 52.940000 51.715000 53.140000 51.915000 ;
        RECT 52.940000 52.135000 53.140000 52.335000 ;
        RECT 52.940000 52.555000 53.140000 52.755000 ;
        RECT 53.315000 47.800000 53.515000 48.000000 ;
        RECT 53.315000 56.470000 53.515000 56.670000 ;
        RECT 53.345000 36.820000 53.545000 37.020000 ;
        RECT 53.345000 37.260000 53.545000 37.460000 ;
        RECT 53.345000 37.700000 53.545000 37.900000 ;
        RECT 53.345000 38.140000 53.545000 38.340000 ;
        RECT 53.345000 38.580000 53.545000 38.780000 ;
        RECT 53.345000 39.020000 53.545000 39.220000 ;
        RECT 53.345000 39.460000 53.545000 39.660000 ;
        RECT 53.345000 39.900000 53.545000 40.100000 ;
        RECT 53.345000 51.715000 53.545000 51.915000 ;
        RECT 53.345000 52.135000 53.545000 52.335000 ;
        RECT 53.345000 52.555000 53.545000 52.755000 ;
        RECT 53.720000 47.800000 53.920000 48.000000 ;
        RECT 53.720000 56.470000 53.920000 56.670000 ;
        RECT 53.750000 36.820000 53.950000 37.020000 ;
        RECT 53.750000 37.260000 53.950000 37.460000 ;
        RECT 53.750000 37.700000 53.950000 37.900000 ;
        RECT 53.750000 38.140000 53.950000 38.340000 ;
        RECT 53.750000 38.580000 53.950000 38.780000 ;
        RECT 53.750000 39.020000 53.950000 39.220000 ;
        RECT 53.750000 39.460000 53.950000 39.660000 ;
        RECT 53.750000 39.900000 53.950000 40.100000 ;
        RECT 53.750000 51.715000 53.950000 51.915000 ;
        RECT 53.750000 52.135000 53.950000 52.335000 ;
        RECT 53.750000 52.555000 53.950000 52.755000 ;
        RECT 54.125000 47.800000 54.325000 48.000000 ;
        RECT 54.125000 56.470000 54.325000 56.670000 ;
        RECT 54.155000 36.820000 54.355000 37.020000 ;
        RECT 54.155000 37.260000 54.355000 37.460000 ;
        RECT 54.155000 37.700000 54.355000 37.900000 ;
        RECT 54.155000 38.140000 54.355000 38.340000 ;
        RECT 54.155000 38.580000 54.355000 38.780000 ;
        RECT 54.155000 39.020000 54.355000 39.220000 ;
        RECT 54.155000 39.460000 54.355000 39.660000 ;
        RECT 54.155000 39.900000 54.355000 40.100000 ;
        RECT 54.155000 51.715000 54.355000 51.915000 ;
        RECT 54.155000 52.135000 54.355000 52.335000 ;
        RECT 54.155000 52.555000 54.355000 52.755000 ;
        RECT 54.530000 47.800000 54.730000 48.000000 ;
        RECT 54.530000 56.470000 54.730000 56.670000 ;
        RECT 54.560000 36.820000 54.760000 37.020000 ;
        RECT 54.560000 37.260000 54.760000 37.460000 ;
        RECT 54.560000 37.700000 54.760000 37.900000 ;
        RECT 54.560000 38.140000 54.760000 38.340000 ;
        RECT 54.560000 38.580000 54.760000 38.780000 ;
        RECT 54.560000 39.020000 54.760000 39.220000 ;
        RECT 54.560000 39.460000 54.760000 39.660000 ;
        RECT 54.560000 39.900000 54.760000 40.100000 ;
        RECT 54.560000 51.715000 54.760000 51.915000 ;
        RECT 54.560000 52.135000 54.760000 52.335000 ;
        RECT 54.560000 52.555000 54.760000 52.755000 ;
        RECT 54.935000 47.800000 55.135000 48.000000 ;
        RECT 54.935000 56.470000 55.135000 56.670000 ;
        RECT 54.965000 36.820000 55.165000 37.020000 ;
        RECT 54.965000 37.260000 55.165000 37.460000 ;
        RECT 54.965000 37.700000 55.165000 37.900000 ;
        RECT 54.965000 38.140000 55.165000 38.340000 ;
        RECT 54.965000 38.580000 55.165000 38.780000 ;
        RECT 54.965000 39.020000 55.165000 39.220000 ;
        RECT 54.965000 39.460000 55.165000 39.660000 ;
        RECT 54.965000 39.900000 55.165000 40.100000 ;
        RECT 54.965000 51.715000 55.165000 51.915000 ;
        RECT 54.965000 52.135000 55.165000 52.335000 ;
        RECT 54.965000 52.555000 55.165000 52.755000 ;
        RECT 55.340000 47.800000 55.540000 48.000000 ;
        RECT 55.340000 56.470000 55.540000 56.670000 ;
        RECT 55.370000 36.820000 55.570000 37.020000 ;
        RECT 55.370000 37.260000 55.570000 37.460000 ;
        RECT 55.370000 37.700000 55.570000 37.900000 ;
        RECT 55.370000 38.140000 55.570000 38.340000 ;
        RECT 55.370000 38.580000 55.570000 38.780000 ;
        RECT 55.370000 39.020000 55.570000 39.220000 ;
        RECT 55.370000 39.460000 55.570000 39.660000 ;
        RECT 55.370000 39.900000 55.570000 40.100000 ;
        RECT 55.370000 51.715000 55.570000 51.915000 ;
        RECT 55.370000 52.135000 55.570000 52.335000 ;
        RECT 55.370000 52.555000 55.570000 52.755000 ;
        RECT 55.745000 47.800000 55.945000 48.000000 ;
        RECT 55.745000 56.470000 55.945000 56.670000 ;
        RECT 55.775000 36.820000 55.975000 37.020000 ;
        RECT 55.775000 37.260000 55.975000 37.460000 ;
        RECT 55.775000 37.700000 55.975000 37.900000 ;
        RECT 55.775000 38.140000 55.975000 38.340000 ;
        RECT 55.775000 38.580000 55.975000 38.780000 ;
        RECT 55.775000 39.020000 55.975000 39.220000 ;
        RECT 55.775000 39.460000 55.975000 39.660000 ;
        RECT 55.775000 39.900000 55.975000 40.100000 ;
        RECT 55.775000 51.715000 55.975000 51.915000 ;
        RECT 55.775000 52.135000 55.975000 52.335000 ;
        RECT 55.775000 52.555000 55.975000 52.755000 ;
        RECT 56.150000 47.800000 56.350000 48.000000 ;
        RECT 56.150000 56.470000 56.350000 56.670000 ;
        RECT 56.180000 36.820000 56.380000 37.020000 ;
        RECT 56.180000 37.260000 56.380000 37.460000 ;
        RECT 56.180000 37.700000 56.380000 37.900000 ;
        RECT 56.180000 38.140000 56.380000 38.340000 ;
        RECT 56.180000 38.580000 56.380000 38.780000 ;
        RECT 56.180000 39.020000 56.380000 39.220000 ;
        RECT 56.180000 39.460000 56.380000 39.660000 ;
        RECT 56.180000 39.900000 56.380000 40.100000 ;
        RECT 56.180000 51.715000 56.380000 51.915000 ;
        RECT 56.180000 52.135000 56.380000 52.335000 ;
        RECT 56.180000 52.555000 56.380000 52.755000 ;
        RECT 56.555000 47.800000 56.755000 48.000000 ;
        RECT 56.555000 56.470000 56.755000 56.670000 ;
        RECT 56.585000 36.820000 56.785000 37.020000 ;
        RECT 56.585000 37.260000 56.785000 37.460000 ;
        RECT 56.585000 37.700000 56.785000 37.900000 ;
        RECT 56.585000 38.140000 56.785000 38.340000 ;
        RECT 56.585000 38.580000 56.785000 38.780000 ;
        RECT 56.585000 39.020000 56.785000 39.220000 ;
        RECT 56.585000 39.460000 56.785000 39.660000 ;
        RECT 56.585000 39.900000 56.785000 40.100000 ;
        RECT 56.585000 51.715000 56.785000 51.915000 ;
        RECT 56.585000 52.135000 56.785000 52.335000 ;
        RECT 56.585000 52.555000 56.785000 52.755000 ;
        RECT 56.960000 47.800000 57.160000 48.000000 ;
        RECT 56.960000 56.470000 57.160000 56.670000 ;
        RECT 56.990000 36.820000 57.190000 37.020000 ;
        RECT 56.990000 37.260000 57.190000 37.460000 ;
        RECT 56.990000 37.700000 57.190000 37.900000 ;
        RECT 56.990000 38.140000 57.190000 38.340000 ;
        RECT 56.990000 38.580000 57.190000 38.780000 ;
        RECT 56.990000 39.020000 57.190000 39.220000 ;
        RECT 56.990000 39.460000 57.190000 39.660000 ;
        RECT 56.990000 39.900000 57.190000 40.100000 ;
        RECT 56.990000 51.715000 57.190000 51.915000 ;
        RECT 56.990000 52.135000 57.190000 52.335000 ;
        RECT 56.990000 52.555000 57.190000 52.755000 ;
        RECT 57.365000 47.800000 57.565000 48.000000 ;
        RECT 57.365000 56.470000 57.565000 56.670000 ;
        RECT 57.395000 36.820000 57.595000 37.020000 ;
        RECT 57.395000 37.260000 57.595000 37.460000 ;
        RECT 57.395000 37.700000 57.595000 37.900000 ;
        RECT 57.395000 38.140000 57.595000 38.340000 ;
        RECT 57.395000 38.580000 57.595000 38.780000 ;
        RECT 57.395000 39.020000 57.595000 39.220000 ;
        RECT 57.395000 39.460000 57.595000 39.660000 ;
        RECT 57.395000 39.900000 57.595000 40.100000 ;
        RECT 57.395000 51.715000 57.595000 51.915000 ;
        RECT 57.395000 52.135000 57.595000 52.335000 ;
        RECT 57.395000 52.555000 57.595000 52.755000 ;
        RECT 57.770000 47.800000 57.970000 48.000000 ;
        RECT 57.770000 56.470000 57.970000 56.670000 ;
        RECT 57.800000 36.820000 58.000000 37.020000 ;
        RECT 57.800000 37.260000 58.000000 37.460000 ;
        RECT 57.800000 37.700000 58.000000 37.900000 ;
        RECT 57.800000 38.140000 58.000000 38.340000 ;
        RECT 57.800000 38.580000 58.000000 38.780000 ;
        RECT 57.800000 39.020000 58.000000 39.220000 ;
        RECT 57.800000 39.460000 58.000000 39.660000 ;
        RECT 57.800000 39.900000 58.000000 40.100000 ;
        RECT 57.800000 51.715000 58.000000 51.915000 ;
        RECT 57.800000 52.135000 58.000000 52.335000 ;
        RECT 57.800000 52.555000 58.000000 52.755000 ;
        RECT 58.175000 47.800000 58.375000 48.000000 ;
        RECT 58.175000 56.470000 58.375000 56.670000 ;
        RECT 58.205000 36.820000 58.405000 37.020000 ;
        RECT 58.205000 37.260000 58.405000 37.460000 ;
        RECT 58.205000 37.700000 58.405000 37.900000 ;
        RECT 58.205000 38.140000 58.405000 38.340000 ;
        RECT 58.205000 38.580000 58.405000 38.780000 ;
        RECT 58.205000 39.020000 58.405000 39.220000 ;
        RECT 58.205000 39.460000 58.405000 39.660000 ;
        RECT 58.205000 39.900000 58.405000 40.100000 ;
        RECT 58.205000 51.715000 58.405000 51.915000 ;
        RECT 58.205000 52.135000 58.405000 52.335000 ;
        RECT 58.205000 52.555000 58.405000 52.755000 ;
        RECT 58.580000 47.800000 58.780000 48.000000 ;
        RECT 58.580000 56.470000 58.780000 56.670000 ;
        RECT 58.610000 36.820000 58.810000 37.020000 ;
        RECT 58.610000 37.260000 58.810000 37.460000 ;
        RECT 58.610000 37.700000 58.810000 37.900000 ;
        RECT 58.610000 38.140000 58.810000 38.340000 ;
        RECT 58.610000 38.580000 58.810000 38.780000 ;
        RECT 58.610000 39.020000 58.810000 39.220000 ;
        RECT 58.610000 39.460000 58.810000 39.660000 ;
        RECT 58.610000 39.900000 58.810000 40.100000 ;
        RECT 58.610000 51.715000 58.810000 51.915000 ;
        RECT 58.610000 52.135000 58.810000 52.335000 ;
        RECT 58.610000 52.555000 58.810000 52.755000 ;
        RECT 58.985000 47.800000 59.185000 48.000000 ;
        RECT 58.985000 56.470000 59.185000 56.670000 ;
        RECT 59.015000 36.820000 59.215000 37.020000 ;
        RECT 59.015000 37.260000 59.215000 37.460000 ;
        RECT 59.015000 37.700000 59.215000 37.900000 ;
        RECT 59.015000 38.140000 59.215000 38.340000 ;
        RECT 59.015000 38.580000 59.215000 38.780000 ;
        RECT 59.015000 39.020000 59.215000 39.220000 ;
        RECT 59.015000 39.460000 59.215000 39.660000 ;
        RECT 59.015000 39.900000 59.215000 40.100000 ;
        RECT 59.015000 51.715000 59.215000 51.915000 ;
        RECT 59.015000 52.135000 59.215000 52.335000 ;
        RECT 59.015000 52.555000 59.215000 52.755000 ;
        RECT 59.390000 47.800000 59.590000 48.000000 ;
        RECT 59.390000 56.470000 59.590000 56.670000 ;
        RECT 59.420000 36.820000 59.620000 37.020000 ;
        RECT 59.420000 37.260000 59.620000 37.460000 ;
        RECT 59.420000 37.700000 59.620000 37.900000 ;
        RECT 59.420000 38.140000 59.620000 38.340000 ;
        RECT 59.420000 38.580000 59.620000 38.780000 ;
        RECT 59.420000 39.020000 59.620000 39.220000 ;
        RECT 59.420000 39.460000 59.620000 39.660000 ;
        RECT 59.420000 39.900000 59.620000 40.100000 ;
        RECT 59.420000 51.715000 59.620000 51.915000 ;
        RECT 59.420000 52.135000 59.620000 52.335000 ;
        RECT 59.420000 52.555000 59.620000 52.755000 ;
        RECT 59.795000 47.800000 59.995000 48.000000 ;
        RECT 59.795000 56.470000 59.995000 56.670000 ;
        RECT 59.825000 36.820000 60.025000 37.020000 ;
        RECT 59.825000 37.260000 60.025000 37.460000 ;
        RECT 59.825000 37.700000 60.025000 37.900000 ;
        RECT 59.825000 38.140000 60.025000 38.340000 ;
        RECT 59.825000 38.580000 60.025000 38.780000 ;
        RECT 59.825000 39.020000 60.025000 39.220000 ;
        RECT 59.825000 39.460000 60.025000 39.660000 ;
        RECT 59.825000 39.900000 60.025000 40.100000 ;
        RECT 59.825000 51.715000 60.025000 51.915000 ;
        RECT 59.825000 52.135000 60.025000 52.335000 ;
        RECT 59.825000 52.555000 60.025000 52.755000 ;
        RECT 60.200000 47.800000 60.400000 48.000000 ;
        RECT 60.200000 56.470000 60.400000 56.670000 ;
        RECT 60.230000 36.820000 60.430000 37.020000 ;
        RECT 60.230000 37.260000 60.430000 37.460000 ;
        RECT 60.230000 37.700000 60.430000 37.900000 ;
        RECT 60.230000 38.140000 60.430000 38.340000 ;
        RECT 60.230000 38.580000 60.430000 38.780000 ;
        RECT 60.230000 39.020000 60.430000 39.220000 ;
        RECT 60.230000 39.460000 60.430000 39.660000 ;
        RECT 60.230000 39.900000 60.430000 40.100000 ;
        RECT 60.230000 51.715000 60.430000 51.915000 ;
        RECT 60.230000 52.135000 60.430000 52.335000 ;
        RECT 60.230000 52.555000 60.430000 52.755000 ;
        RECT 60.605000 47.800000 60.805000 48.000000 ;
        RECT 60.605000 56.470000 60.805000 56.670000 ;
        RECT 60.635000 36.820000 60.835000 37.020000 ;
        RECT 60.635000 37.260000 60.835000 37.460000 ;
        RECT 60.635000 37.700000 60.835000 37.900000 ;
        RECT 60.635000 38.140000 60.835000 38.340000 ;
        RECT 60.635000 38.580000 60.835000 38.780000 ;
        RECT 60.635000 39.020000 60.835000 39.220000 ;
        RECT 60.635000 39.460000 60.835000 39.660000 ;
        RECT 60.635000 39.900000 60.835000 40.100000 ;
        RECT 60.635000 51.715000 60.835000 51.915000 ;
        RECT 60.635000 52.135000 60.835000 52.335000 ;
        RECT 60.635000 52.555000 60.835000 52.755000 ;
        RECT 61.010000 47.800000 61.210000 48.000000 ;
        RECT 61.010000 56.470000 61.210000 56.670000 ;
        RECT 61.040000 36.820000 61.240000 37.020000 ;
        RECT 61.040000 37.260000 61.240000 37.460000 ;
        RECT 61.040000 37.700000 61.240000 37.900000 ;
        RECT 61.040000 38.140000 61.240000 38.340000 ;
        RECT 61.040000 38.580000 61.240000 38.780000 ;
        RECT 61.040000 39.020000 61.240000 39.220000 ;
        RECT 61.040000 39.460000 61.240000 39.660000 ;
        RECT 61.040000 39.900000 61.240000 40.100000 ;
        RECT 61.040000 51.715000 61.240000 51.915000 ;
        RECT 61.040000 52.135000 61.240000 52.335000 ;
        RECT 61.040000 52.555000 61.240000 52.755000 ;
        RECT 61.415000 47.800000 61.615000 48.000000 ;
        RECT 61.415000 56.470000 61.615000 56.670000 ;
        RECT 61.445000 36.820000 61.645000 37.020000 ;
        RECT 61.445000 37.260000 61.645000 37.460000 ;
        RECT 61.445000 37.700000 61.645000 37.900000 ;
        RECT 61.445000 38.140000 61.645000 38.340000 ;
        RECT 61.445000 38.580000 61.645000 38.780000 ;
        RECT 61.445000 39.020000 61.645000 39.220000 ;
        RECT 61.445000 39.460000 61.645000 39.660000 ;
        RECT 61.445000 39.900000 61.645000 40.100000 ;
        RECT 61.445000 51.715000 61.645000 51.915000 ;
        RECT 61.445000 52.135000 61.645000 52.335000 ;
        RECT 61.445000 52.555000 61.645000 52.755000 ;
        RECT 61.820000 47.800000 62.020000 48.000000 ;
        RECT 61.820000 56.470000 62.020000 56.670000 ;
        RECT 61.850000 36.820000 62.050000 37.020000 ;
        RECT 61.850000 37.260000 62.050000 37.460000 ;
        RECT 61.850000 37.700000 62.050000 37.900000 ;
        RECT 61.850000 38.140000 62.050000 38.340000 ;
        RECT 61.850000 38.580000 62.050000 38.780000 ;
        RECT 61.850000 39.020000 62.050000 39.220000 ;
        RECT 61.850000 39.460000 62.050000 39.660000 ;
        RECT 61.850000 39.900000 62.050000 40.100000 ;
        RECT 61.850000 51.715000 62.050000 51.915000 ;
        RECT 61.850000 52.135000 62.050000 52.335000 ;
        RECT 61.850000 52.555000 62.050000 52.755000 ;
        RECT 62.225000 47.800000 62.425000 48.000000 ;
        RECT 62.225000 56.470000 62.425000 56.670000 ;
        RECT 62.255000 36.820000 62.455000 37.020000 ;
        RECT 62.255000 37.260000 62.455000 37.460000 ;
        RECT 62.255000 37.700000 62.455000 37.900000 ;
        RECT 62.255000 38.140000 62.455000 38.340000 ;
        RECT 62.255000 38.580000 62.455000 38.780000 ;
        RECT 62.255000 39.020000 62.455000 39.220000 ;
        RECT 62.255000 39.460000 62.455000 39.660000 ;
        RECT 62.255000 39.900000 62.455000 40.100000 ;
        RECT 62.255000 51.715000 62.455000 51.915000 ;
        RECT 62.255000 52.135000 62.455000 52.335000 ;
        RECT 62.255000 52.555000 62.455000 52.755000 ;
        RECT 62.630000 47.800000 62.830000 48.000000 ;
        RECT 62.630000 56.470000 62.830000 56.670000 ;
        RECT 62.660000 36.820000 62.860000 37.020000 ;
        RECT 62.660000 37.260000 62.860000 37.460000 ;
        RECT 62.660000 37.700000 62.860000 37.900000 ;
        RECT 62.660000 38.140000 62.860000 38.340000 ;
        RECT 62.660000 38.580000 62.860000 38.780000 ;
        RECT 62.660000 39.020000 62.860000 39.220000 ;
        RECT 62.660000 39.460000 62.860000 39.660000 ;
        RECT 62.660000 39.900000 62.860000 40.100000 ;
        RECT 62.660000 51.715000 62.860000 51.915000 ;
        RECT 62.660000 52.135000 62.860000 52.335000 ;
        RECT 62.660000 52.555000 62.860000 52.755000 ;
        RECT 63.035000 47.800000 63.235000 48.000000 ;
        RECT 63.035000 56.470000 63.235000 56.670000 ;
        RECT 63.065000 36.820000 63.265000 37.020000 ;
        RECT 63.065000 37.260000 63.265000 37.460000 ;
        RECT 63.065000 37.700000 63.265000 37.900000 ;
        RECT 63.065000 38.140000 63.265000 38.340000 ;
        RECT 63.065000 38.580000 63.265000 38.780000 ;
        RECT 63.065000 39.020000 63.265000 39.220000 ;
        RECT 63.065000 39.460000 63.265000 39.660000 ;
        RECT 63.065000 39.900000 63.265000 40.100000 ;
        RECT 63.065000 51.715000 63.265000 51.915000 ;
        RECT 63.065000 52.135000 63.265000 52.335000 ;
        RECT 63.065000 52.555000 63.265000 52.755000 ;
        RECT 63.440000 47.800000 63.640000 48.000000 ;
        RECT 63.440000 56.470000 63.640000 56.670000 ;
        RECT 63.470000 36.820000 63.670000 37.020000 ;
        RECT 63.470000 37.260000 63.670000 37.460000 ;
        RECT 63.470000 37.700000 63.670000 37.900000 ;
        RECT 63.470000 38.140000 63.670000 38.340000 ;
        RECT 63.470000 38.580000 63.670000 38.780000 ;
        RECT 63.470000 39.020000 63.670000 39.220000 ;
        RECT 63.470000 39.460000 63.670000 39.660000 ;
        RECT 63.470000 39.900000 63.670000 40.100000 ;
        RECT 63.470000 51.715000 63.670000 51.915000 ;
        RECT 63.470000 52.135000 63.670000 52.335000 ;
        RECT 63.470000 52.555000 63.670000 52.755000 ;
        RECT 63.845000 47.800000 64.045000 48.000000 ;
        RECT 63.845000 56.470000 64.045000 56.670000 ;
        RECT 63.875000 36.820000 64.075000 37.020000 ;
        RECT 63.875000 37.260000 64.075000 37.460000 ;
        RECT 63.875000 37.700000 64.075000 37.900000 ;
        RECT 63.875000 38.140000 64.075000 38.340000 ;
        RECT 63.875000 38.580000 64.075000 38.780000 ;
        RECT 63.875000 39.020000 64.075000 39.220000 ;
        RECT 63.875000 39.460000 64.075000 39.660000 ;
        RECT 63.875000 39.900000 64.075000 40.100000 ;
        RECT 63.875000 51.715000 64.075000 51.915000 ;
        RECT 63.875000 52.135000 64.075000 52.335000 ;
        RECT 63.875000 52.555000 64.075000 52.755000 ;
        RECT 64.250000 47.800000 64.450000 48.000000 ;
        RECT 64.250000 56.470000 64.450000 56.670000 ;
        RECT 64.280000 36.820000 64.480000 37.020000 ;
        RECT 64.280000 37.260000 64.480000 37.460000 ;
        RECT 64.280000 37.700000 64.480000 37.900000 ;
        RECT 64.280000 38.140000 64.480000 38.340000 ;
        RECT 64.280000 38.580000 64.480000 38.780000 ;
        RECT 64.280000 39.020000 64.480000 39.220000 ;
        RECT 64.280000 39.460000 64.480000 39.660000 ;
        RECT 64.280000 39.900000 64.480000 40.100000 ;
        RECT 64.280000 51.715000 64.480000 51.915000 ;
        RECT 64.280000 52.135000 64.480000 52.335000 ;
        RECT 64.280000 52.555000 64.480000 52.755000 ;
        RECT 64.655000 47.800000 64.855000 48.000000 ;
        RECT 64.655000 56.470000 64.855000 56.670000 ;
        RECT 64.685000 36.820000 64.885000 37.020000 ;
        RECT 64.685000 37.260000 64.885000 37.460000 ;
        RECT 64.685000 37.700000 64.885000 37.900000 ;
        RECT 64.685000 38.140000 64.885000 38.340000 ;
        RECT 64.685000 38.580000 64.885000 38.780000 ;
        RECT 64.685000 39.020000 64.885000 39.220000 ;
        RECT 64.685000 39.460000 64.885000 39.660000 ;
        RECT 64.685000 39.900000 64.885000 40.100000 ;
        RECT 64.685000 51.715000 64.885000 51.915000 ;
        RECT 64.685000 52.135000 64.885000 52.335000 ;
        RECT 64.685000 52.555000 64.885000 52.755000 ;
        RECT 65.060000 47.800000 65.260000 48.000000 ;
        RECT 65.060000 56.470000 65.260000 56.670000 ;
        RECT 65.090000 36.820000 65.290000 37.020000 ;
        RECT 65.090000 37.260000 65.290000 37.460000 ;
        RECT 65.090000 37.700000 65.290000 37.900000 ;
        RECT 65.090000 38.140000 65.290000 38.340000 ;
        RECT 65.090000 38.580000 65.290000 38.780000 ;
        RECT 65.090000 39.020000 65.290000 39.220000 ;
        RECT 65.090000 39.460000 65.290000 39.660000 ;
        RECT 65.090000 39.900000 65.290000 40.100000 ;
        RECT 65.090000 51.715000 65.290000 51.915000 ;
        RECT 65.090000 52.135000 65.290000 52.335000 ;
        RECT 65.090000 52.555000 65.290000 52.755000 ;
        RECT 65.465000 47.800000 65.665000 48.000000 ;
        RECT 65.465000 56.470000 65.665000 56.670000 ;
        RECT 65.495000 36.820000 65.695000 37.020000 ;
        RECT 65.495000 37.260000 65.695000 37.460000 ;
        RECT 65.495000 37.700000 65.695000 37.900000 ;
        RECT 65.495000 38.140000 65.695000 38.340000 ;
        RECT 65.495000 38.580000 65.695000 38.780000 ;
        RECT 65.495000 39.020000 65.695000 39.220000 ;
        RECT 65.495000 39.460000 65.695000 39.660000 ;
        RECT 65.495000 39.900000 65.695000 40.100000 ;
        RECT 65.495000 51.715000 65.695000 51.915000 ;
        RECT 65.495000 52.135000 65.695000 52.335000 ;
        RECT 65.495000 52.555000 65.695000 52.755000 ;
        RECT 65.870000 47.800000 66.070000 48.000000 ;
        RECT 65.870000 56.470000 66.070000 56.670000 ;
        RECT 65.900000 36.820000 66.100000 37.020000 ;
        RECT 65.900000 37.260000 66.100000 37.460000 ;
        RECT 65.900000 37.700000 66.100000 37.900000 ;
        RECT 65.900000 38.140000 66.100000 38.340000 ;
        RECT 65.900000 38.580000 66.100000 38.780000 ;
        RECT 65.900000 39.020000 66.100000 39.220000 ;
        RECT 65.900000 39.460000 66.100000 39.660000 ;
        RECT 65.900000 39.900000 66.100000 40.100000 ;
        RECT 65.900000 51.715000 66.100000 51.915000 ;
        RECT 65.900000 52.135000 66.100000 52.335000 ;
        RECT 65.900000 52.555000 66.100000 52.755000 ;
        RECT 66.275000 47.800000 66.475000 48.000000 ;
        RECT 66.275000 56.470000 66.475000 56.670000 ;
        RECT 66.305000 36.820000 66.505000 37.020000 ;
        RECT 66.305000 37.260000 66.505000 37.460000 ;
        RECT 66.305000 37.700000 66.505000 37.900000 ;
        RECT 66.305000 38.140000 66.505000 38.340000 ;
        RECT 66.305000 38.580000 66.505000 38.780000 ;
        RECT 66.305000 39.020000 66.505000 39.220000 ;
        RECT 66.305000 39.460000 66.505000 39.660000 ;
        RECT 66.305000 39.900000 66.505000 40.100000 ;
        RECT 66.305000 51.715000 66.505000 51.915000 ;
        RECT 66.305000 52.135000 66.505000 52.335000 ;
        RECT 66.305000 52.555000 66.505000 52.755000 ;
        RECT 66.680000 47.800000 66.880000 48.000000 ;
        RECT 66.680000 56.470000 66.880000 56.670000 ;
        RECT 66.710000 36.820000 66.910000 37.020000 ;
        RECT 66.710000 37.260000 66.910000 37.460000 ;
        RECT 66.710000 37.700000 66.910000 37.900000 ;
        RECT 66.710000 38.140000 66.910000 38.340000 ;
        RECT 66.710000 38.580000 66.910000 38.780000 ;
        RECT 66.710000 39.020000 66.910000 39.220000 ;
        RECT 66.710000 39.460000 66.910000 39.660000 ;
        RECT 66.710000 39.900000 66.910000 40.100000 ;
        RECT 66.710000 51.715000 66.910000 51.915000 ;
        RECT 66.710000 52.135000 66.910000 52.335000 ;
        RECT 66.710000 52.555000 66.910000 52.755000 ;
        RECT 67.085000 47.800000 67.285000 48.000000 ;
        RECT 67.085000 56.470000 67.285000 56.670000 ;
        RECT 67.115000 36.820000 67.315000 37.020000 ;
        RECT 67.115000 37.260000 67.315000 37.460000 ;
        RECT 67.115000 37.700000 67.315000 37.900000 ;
        RECT 67.115000 38.140000 67.315000 38.340000 ;
        RECT 67.115000 38.580000 67.315000 38.780000 ;
        RECT 67.115000 39.020000 67.315000 39.220000 ;
        RECT 67.115000 39.460000 67.315000 39.660000 ;
        RECT 67.115000 39.900000 67.315000 40.100000 ;
        RECT 67.115000 51.715000 67.315000 51.915000 ;
        RECT 67.115000 52.135000 67.315000 52.335000 ;
        RECT 67.115000 52.555000 67.315000 52.755000 ;
        RECT 67.490000 47.800000 67.690000 48.000000 ;
        RECT 67.490000 56.470000 67.690000 56.670000 ;
        RECT 67.520000 36.820000 67.720000 37.020000 ;
        RECT 67.520000 37.260000 67.720000 37.460000 ;
        RECT 67.520000 37.700000 67.720000 37.900000 ;
        RECT 67.520000 38.140000 67.720000 38.340000 ;
        RECT 67.520000 38.580000 67.720000 38.780000 ;
        RECT 67.520000 39.020000 67.720000 39.220000 ;
        RECT 67.520000 39.460000 67.720000 39.660000 ;
        RECT 67.520000 39.900000 67.720000 40.100000 ;
        RECT 67.520000 51.715000 67.720000 51.915000 ;
        RECT 67.520000 52.135000 67.720000 52.335000 ;
        RECT 67.520000 52.555000 67.720000 52.755000 ;
        RECT 67.895000 47.800000 68.095000 48.000000 ;
        RECT 67.895000 56.470000 68.095000 56.670000 ;
        RECT 67.925000 36.820000 68.125000 37.020000 ;
        RECT 67.925000 37.260000 68.125000 37.460000 ;
        RECT 67.925000 37.700000 68.125000 37.900000 ;
        RECT 67.925000 38.140000 68.125000 38.340000 ;
        RECT 67.925000 38.580000 68.125000 38.780000 ;
        RECT 67.925000 39.020000 68.125000 39.220000 ;
        RECT 67.925000 39.460000 68.125000 39.660000 ;
        RECT 67.925000 39.900000 68.125000 40.100000 ;
        RECT 67.925000 51.715000 68.125000 51.915000 ;
        RECT 67.925000 52.135000 68.125000 52.335000 ;
        RECT 67.925000 52.555000 68.125000 52.755000 ;
        RECT 68.300000 47.800000 68.500000 48.000000 ;
        RECT 68.300000 56.470000 68.500000 56.670000 ;
        RECT 68.330000 36.820000 68.530000 37.020000 ;
        RECT 68.330000 37.260000 68.530000 37.460000 ;
        RECT 68.330000 37.700000 68.530000 37.900000 ;
        RECT 68.330000 38.140000 68.530000 38.340000 ;
        RECT 68.330000 38.580000 68.530000 38.780000 ;
        RECT 68.330000 39.020000 68.530000 39.220000 ;
        RECT 68.330000 39.460000 68.530000 39.660000 ;
        RECT 68.330000 39.900000 68.530000 40.100000 ;
        RECT 68.330000 51.715000 68.530000 51.915000 ;
        RECT 68.330000 52.135000 68.530000 52.335000 ;
        RECT 68.330000 52.555000 68.530000 52.755000 ;
        RECT 68.705000 47.800000 68.905000 48.000000 ;
        RECT 68.705000 56.470000 68.905000 56.670000 ;
        RECT 68.735000 36.820000 68.935000 37.020000 ;
        RECT 68.735000 37.260000 68.935000 37.460000 ;
        RECT 68.735000 37.700000 68.935000 37.900000 ;
        RECT 68.735000 38.140000 68.935000 38.340000 ;
        RECT 68.735000 38.580000 68.935000 38.780000 ;
        RECT 68.735000 39.020000 68.935000 39.220000 ;
        RECT 68.735000 39.460000 68.935000 39.660000 ;
        RECT 68.735000 39.900000 68.935000 40.100000 ;
        RECT 68.735000 51.715000 68.935000 51.915000 ;
        RECT 68.735000 52.135000 68.935000 52.335000 ;
        RECT 68.735000 52.555000 68.935000 52.755000 ;
        RECT 69.110000 47.800000 69.310000 48.000000 ;
        RECT 69.110000 56.470000 69.310000 56.670000 ;
        RECT 69.140000 36.820000 69.340000 37.020000 ;
        RECT 69.140000 37.260000 69.340000 37.460000 ;
        RECT 69.140000 37.700000 69.340000 37.900000 ;
        RECT 69.140000 38.140000 69.340000 38.340000 ;
        RECT 69.140000 38.580000 69.340000 38.780000 ;
        RECT 69.140000 39.020000 69.340000 39.220000 ;
        RECT 69.140000 39.460000 69.340000 39.660000 ;
        RECT 69.140000 39.900000 69.340000 40.100000 ;
        RECT 69.140000 51.715000 69.340000 51.915000 ;
        RECT 69.140000 52.135000 69.340000 52.335000 ;
        RECT 69.140000 52.555000 69.340000 52.755000 ;
        RECT 69.515000 47.800000 69.715000 48.000000 ;
        RECT 69.515000 56.470000 69.715000 56.670000 ;
        RECT 69.545000 36.820000 69.745000 37.020000 ;
        RECT 69.545000 37.260000 69.745000 37.460000 ;
        RECT 69.545000 37.700000 69.745000 37.900000 ;
        RECT 69.545000 38.140000 69.745000 38.340000 ;
        RECT 69.545000 38.580000 69.745000 38.780000 ;
        RECT 69.545000 39.020000 69.745000 39.220000 ;
        RECT 69.545000 39.460000 69.745000 39.660000 ;
        RECT 69.545000 39.900000 69.745000 40.100000 ;
        RECT 69.545000 51.715000 69.745000 51.915000 ;
        RECT 69.545000 52.135000 69.745000 52.335000 ;
        RECT 69.545000 52.555000 69.745000 52.755000 ;
        RECT 69.920000 47.800000 70.120000 48.000000 ;
        RECT 69.920000 56.470000 70.120000 56.670000 ;
        RECT 69.950000 36.820000 70.150000 37.020000 ;
        RECT 69.950000 37.260000 70.150000 37.460000 ;
        RECT 69.950000 37.700000 70.150000 37.900000 ;
        RECT 69.950000 38.140000 70.150000 38.340000 ;
        RECT 69.950000 38.580000 70.150000 38.780000 ;
        RECT 69.950000 39.020000 70.150000 39.220000 ;
        RECT 69.950000 39.460000 70.150000 39.660000 ;
        RECT 69.950000 39.900000 70.150000 40.100000 ;
        RECT 69.950000 51.715000 70.150000 51.915000 ;
        RECT 69.950000 52.135000 70.150000 52.335000 ;
        RECT 69.950000 52.555000 70.150000 52.755000 ;
        RECT 70.325000 47.800000 70.525000 48.000000 ;
        RECT 70.325000 56.470000 70.525000 56.670000 ;
        RECT 70.355000 36.820000 70.555000 37.020000 ;
        RECT 70.355000 37.260000 70.555000 37.460000 ;
        RECT 70.355000 37.700000 70.555000 37.900000 ;
        RECT 70.355000 38.140000 70.555000 38.340000 ;
        RECT 70.355000 38.580000 70.555000 38.780000 ;
        RECT 70.355000 39.020000 70.555000 39.220000 ;
        RECT 70.355000 39.460000 70.555000 39.660000 ;
        RECT 70.355000 39.900000 70.555000 40.100000 ;
        RECT 70.355000 51.715000 70.555000 51.915000 ;
        RECT 70.355000 52.135000 70.555000 52.335000 ;
        RECT 70.355000 52.555000 70.555000 52.755000 ;
        RECT 70.730000 47.800000 70.930000 48.000000 ;
        RECT 70.730000 56.470000 70.930000 56.670000 ;
        RECT 70.760000 36.820000 70.960000 37.020000 ;
        RECT 70.760000 37.260000 70.960000 37.460000 ;
        RECT 70.760000 37.700000 70.960000 37.900000 ;
        RECT 70.760000 38.140000 70.960000 38.340000 ;
        RECT 70.760000 38.580000 70.960000 38.780000 ;
        RECT 70.760000 39.020000 70.960000 39.220000 ;
        RECT 70.760000 39.460000 70.960000 39.660000 ;
        RECT 70.760000 39.900000 70.960000 40.100000 ;
        RECT 70.760000 51.715000 70.960000 51.915000 ;
        RECT 70.760000 52.135000 70.960000 52.335000 ;
        RECT 70.760000 52.555000 70.960000 52.755000 ;
        RECT 71.135000 47.800000 71.335000 48.000000 ;
        RECT 71.135000 56.470000 71.335000 56.670000 ;
        RECT 71.165000 36.820000 71.365000 37.020000 ;
        RECT 71.165000 37.260000 71.365000 37.460000 ;
        RECT 71.165000 37.700000 71.365000 37.900000 ;
        RECT 71.165000 38.140000 71.365000 38.340000 ;
        RECT 71.165000 38.580000 71.365000 38.780000 ;
        RECT 71.165000 39.020000 71.365000 39.220000 ;
        RECT 71.165000 39.460000 71.365000 39.660000 ;
        RECT 71.165000 39.900000 71.365000 40.100000 ;
        RECT 71.165000 51.715000 71.365000 51.915000 ;
        RECT 71.165000 52.135000 71.365000 52.335000 ;
        RECT 71.165000 52.555000 71.365000 52.755000 ;
        RECT 71.540000 47.800000 71.740000 48.000000 ;
        RECT 71.540000 56.470000 71.740000 56.670000 ;
        RECT 71.570000 36.820000 71.770000 37.020000 ;
        RECT 71.570000 37.260000 71.770000 37.460000 ;
        RECT 71.570000 37.700000 71.770000 37.900000 ;
        RECT 71.570000 38.140000 71.770000 38.340000 ;
        RECT 71.570000 38.580000 71.770000 38.780000 ;
        RECT 71.570000 39.020000 71.770000 39.220000 ;
        RECT 71.570000 39.460000 71.770000 39.660000 ;
        RECT 71.570000 39.900000 71.770000 40.100000 ;
        RECT 71.570000 51.715000 71.770000 51.915000 ;
        RECT 71.570000 52.135000 71.770000 52.335000 ;
        RECT 71.570000 52.555000 71.770000 52.755000 ;
        RECT 71.950000 47.800000 72.150000 48.000000 ;
        RECT 71.950000 56.470000 72.150000 56.670000 ;
        RECT 71.975000 36.820000 72.175000 37.020000 ;
        RECT 71.975000 37.260000 72.175000 37.460000 ;
        RECT 71.975000 37.700000 72.175000 37.900000 ;
        RECT 71.975000 38.140000 72.175000 38.340000 ;
        RECT 71.975000 38.580000 72.175000 38.780000 ;
        RECT 71.975000 39.020000 72.175000 39.220000 ;
        RECT 71.975000 39.460000 72.175000 39.660000 ;
        RECT 71.975000 39.900000 72.175000 40.100000 ;
        RECT 71.975000 51.715000 72.175000 51.915000 ;
        RECT 71.975000 52.135000 72.175000 52.335000 ;
        RECT 71.975000 52.555000 72.175000 52.755000 ;
        RECT 72.360000 47.800000 72.560000 48.000000 ;
        RECT 72.360000 56.470000 72.560000 56.670000 ;
        RECT 72.380000 36.820000 72.580000 37.020000 ;
        RECT 72.380000 37.260000 72.580000 37.460000 ;
        RECT 72.380000 37.700000 72.580000 37.900000 ;
        RECT 72.380000 38.140000 72.580000 38.340000 ;
        RECT 72.380000 38.580000 72.580000 38.780000 ;
        RECT 72.380000 39.020000 72.580000 39.220000 ;
        RECT 72.380000 39.460000 72.580000 39.660000 ;
        RECT 72.380000 39.900000 72.580000 40.100000 ;
        RECT 72.380000 51.715000 72.580000 51.915000 ;
        RECT 72.380000 52.135000 72.580000 52.335000 ;
        RECT 72.380000 52.555000 72.580000 52.755000 ;
        RECT 72.770000 47.800000 72.970000 48.000000 ;
        RECT 72.770000 56.470000 72.970000 56.670000 ;
        RECT 72.785000 36.820000 72.985000 37.020000 ;
        RECT 72.785000 37.260000 72.985000 37.460000 ;
        RECT 72.785000 37.700000 72.985000 37.900000 ;
        RECT 72.785000 38.140000 72.985000 38.340000 ;
        RECT 72.785000 38.580000 72.985000 38.780000 ;
        RECT 72.785000 39.020000 72.985000 39.220000 ;
        RECT 72.785000 39.460000 72.985000 39.660000 ;
        RECT 72.785000 39.900000 72.985000 40.100000 ;
        RECT 72.785000 51.715000 72.985000 51.915000 ;
        RECT 72.785000 52.135000 72.985000 52.335000 ;
        RECT 72.785000 52.555000 72.985000 52.755000 ;
        RECT 73.180000 47.800000 73.380000 48.000000 ;
        RECT 73.180000 56.470000 73.380000 56.670000 ;
        RECT 73.190000 36.820000 73.390000 37.020000 ;
        RECT 73.190000 37.260000 73.390000 37.460000 ;
        RECT 73.190000 37.700000 73.390000 37.900000 ;
        RECT 73.190000 38.140000 73.390000 38.340000 ;
        RECT 73.190000 38.580000 73.390000 38.780000 ;
        RECT 73.190000 39.020000 73.390000 39.220000 ;
        RECT 73.190000 39.460000 73.390000 39.660000 ;
        RECT 73.190000 39.900000 73.390000 40.100000 ;
        RECT 73.190000 51.715000 73.390000 51.915000 ;
        RECT 73.190000 52.135000 73.390000 52.335000 ;
        RECT 73.190000 52.555000 73.390000 52.755000 ;
        RECT 73.590000 47.800000 73.790000 48.000000 ;
        RECT 73.590000 56.470000 73.790000 56.670000 ;
        RECT 73.595000 36.820000 73.795000 37.020000 ;
        RECT 73.595000 37.260000 73.795000 37.460000 ;
        RECT 73.595000 37.700000 73.795000 37.900000 ;
        RECT 73.595000 38.140000 73.795000 38.340000 ;
        RECT 73.595000 38.580000 73.795000 38.780000 ;
        RECT 73.595000 39.020000 73.795000 39.220000 ;
        RECT 73.595000 39.460000 73.795000 39.660000 ;
        RECT 73.595000 39.900000 73.795000 40.100000 ;
        RECT 73.595000 51.715000 73.795000 51.915000 ;
        RECT 73.595000 52.135000 73.795000 52.335000 ;
        RECT 73.595000 52.555000 73.795000 52.755000 ;
        RECT 74.000000 36.820000 74.200000 37.020000 ;
        RECT 74.000000 37.260000 74.200000 37.460000 ;
        RECT 74.000000 37.700000 74.200000 37.900000 ;
        RECT 74.000000 38.140000 74.200000 38.340000 ;
        RECT 74.000000 38.580000 74.200000 38.780000 ;
        RECT 74.000000 39.020000 74.200000 39.220000 ;
        RECT 74.000000 39.460000 74.200000 39.660000 ;
        RECT 74.000000 39.900000 74.200000 40.100000 ;
        RECT 74.000000 47.800000 74.200000 48.000000 ;
        RECT 74.000000 51.715000 74.200000 51.915000 ;
        RECT 74.000000 52.135000 74.200000 52.335000 ;
        RECT 74.000000 52.555000 74.200000 52.755000 ;
        RECT 74.000000 56.470000 74.200000 56.670000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 75.000000  36.340000 ;
      RECT  0.000000 36.340000  0.570000  40.580000 ;
      RECT  0.000000 40.580000 75.000000  47.340000 ;
      RECT  0.000000 48.460000 24.795000  51.250000 ;
      RECT  0.000000 53.220000 24.795000  56.010000 ;
      RECT  0.000000 57.130000 75.000000 200.000000 ;
      RECT 24.795000 36.340000 49.990000  40.580000 ;
      RECT 24.795000 47.340000 49.990000  57.130000 ;
      RECT 49.990000 48.460000 75.000000  51.250000 ;
      RECT 49.990000 53.220000 75.000000  56.010000 ;
      RECT 74.690000 36.340000 75.000000  40.580000 ;
      RECT 74.690000 47.340000 75.000000  48.460000 ;
      RECT 74.690000 51.250000 75.000000  53.220000 ;
      RECT 74.690000 56.010000 75.000000  57.130000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000  19.385000 73.330000  36.335000 ;
      RECT  1.670000  40.585000 73.330000  47.335000 ;
      RECT  1.670000  48.465000 24.770000  51.245000 ;
      RECT  1.670000  53.225000 24.770000  56.005000 ;
      RECT  1.670000  57.135000 73.330000  95.400000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT 24.770000  36.335000 50.015000  40.585000 ;
      RECT 24.770000  47.335000 50.015000  57.135000 ;
      RECT 50.015000  48.465000 73.330000  51.245000 ;
      RECT 50.015000  53.225000 73.330000  56.005000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT 0.000000   0.000000 75.000000   1.335000 ;
      RECT 0.000000  95.785000 75.000000 174.985000 ;
      RECT 1.765000  14.235000 73.235000  19.085000 ;
      RECT 2.070000   1.335000 72.930000  14.235000 ;
      RECT 2.070000  19.085000 72.930000  95.785000 ;
      RECT 2.070000 174.985000 72.930000 200.000000 ;
  END
END sky130_fd_io__overlay_vssa_hvc


END LIBRARY
