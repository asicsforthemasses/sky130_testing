
# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0
#
# Autogenerated by https://www.asicsforthemasses.com
#

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;


MACRO sky130_fd_sc_hdll__clkmux2_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.232200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.290000 0.255000 2.615000 1.415000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.232200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.810000 1.950000 1.615000 ;
        RECT 1.780000 1.615000 3.075000 1.785000 ;
        RECT 2.785000 0.255000 3.075000 1.615000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.479400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 0.995000 1.270000 1.325000 ;
        RECT 1.070000 1.325000 1.270000 2.295000 ;
        RECT 1.070000 2.295000 3.415000 2.465000 ;
        RECT 3.245000 1.440000 3.995000 1.630000 ;
        RECT 3.245000 1.630000 3.415000 2.295000 ;
        RECT 3.805000 1.055000 3.995000 1.440000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.405200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.255000 0.345000 1.495000 ;
        RECT 0.090000 1.495000 0.425000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.515000  0.085000 0.895000 0.485000 ;
      RECT 0.515000  0.655000 1.610000 0.825000 ;
      RECT 0.515000  0.825000 0.685000 1.325000 ;
      RECT 0.645000  1.495000 0.815000 2.635000 ;
      RECT 1.435000  0.255000 1.955000 0.620000 ;
      RECT 1.435000  0.620000 1.610000 0.655000 ;
      RECT 1.440000  0.825000 1.610000 1.955000 ;
      RECT 1.440000  1.955000 2.885000 2.125000 ;
      RECT 3.250000  0.085000 3.765000 0.525000 ;
      RECT 3.325000  0.695000 4.385000 0.865000 ;
      RECT 3.325000  0.865000 3.495000 1.185000 ;
      RECT 3.585000  1.835000 3.815000 2.635000 ;
      RECT 3.985000  1.835000 4.385000 2.465000 ;
      RECT 4.035000  0.255000 4.280000 0.695000 ;
      RECT 4.215000  0.865000 4.385000 1.835000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkmux2_1


MACRO sky130_fd_sc_hdll__clkmux2_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.232200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.670000 0.255000 3.995000 1.415000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.232200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.160000 0.810000 3.330000 1.615000 ;
        RECT 3.160000 1.615000 4.455000 1.785000 ;
        RECT 4.165000 0.255000 4.455000 1.615000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.479400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 0.995000 2.650000 1.325000 ;
        RECT 2.450000 1.325000 2.650000 2.295000 ;
        RECT 2.450000 2.295000 4.795000 2.465000 ;
        RECT 4.625000 1.440000 5.375000 1.630000 ;
        RECT 4.625000 1.630000 4.795000 2.295000 ;
        RECT 5.185000 1.055000 5.375000 1.440000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.860800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.495000 0.895000 2.465000 ;
        RECT 0.590000 0.255000 0.850000 1.065000 ;
        RECT 0.590000 1.065000 1.745000 1.325000 ;
        RECT 0.590000 1.325000 0.850000 1.495000 ;
        RECT 1.475000 0.255000 1.745000 1.065000 ;
        RECT 1.475000 1.325000 1.745000 1.495000 ;
        RECT 1.475000 1.495000 1.835000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.135000  1.495000 0.395000 2.635000 ;
      RECT 0.175000  0.085000 0.420000 0.655000 ;
      RECT 1.055000  0.085000 1.305000 0.655000 ;
      RECT 1.065000  1.495000 1.305000 2.635000 ;
      RECT 1.915000  0.085000 2.275000 0.485000 ;
      RECT 1.915000  0.655000 2.990000 0.825000 ;
      RECT 1.915000  0.825000 2.085000 1.325000 ;
      RECT 2.005000  1.495000 2.280000 2.635000 ;
      RECT 2.815000  0.255000 3.500000 0.620000 ;
      RECT 2.815000  0.620000 2.990000 0.655000 ;
      RECT 2.820000  0.825000 2.990000 1.955000 ;
      RECT 2.820000  1.955000 4.265000 2.125000 ;
      RECT 4.630000  0.085000 5.145000 0.525000 ;
      RECT 4.705000  0.695000 5.765000 0.865000 ;
      RECT 4.705000  0.865000 4.875000 1.185000 ;
      RECT 4.965000  1.835000 5.195000 2.635000 ;
      RECT 5.365000  1.835000 5.765000 2.465000 ;
      RECT 5.415000  0.255000 5.660000 0.695000 ;
      RECT 5.595000  0.865000 5.765000 1.835000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkmux2_4


MACRO sky130_fd_sc_hdll__clkmux2_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.232200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.750000 0.255000 3.075000 1.415000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.232200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.240000 0.810000 2.410000 1.615000 ;
        RECT 2.240000 1.615000 3.535000 1.785000 ;
        RECT 3.245000 0.255000 3.535000 1.615000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.479400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.995000 1.730000 1.325000 ;
        RECT 1.530000 1.325000 1.730000 2.295000 ;
        RECT 1.530000 2.295000 3.875000 2.465000 ;
        RECT 3.705000 1.440000 4.455000 1.630000 ;
        RECT 3.705000 1.630000 3.875000 2.295000 ;
        RECT 4.265000 1.055000 4.455000 1.440000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.430400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.255000 0.805000 1.495000 ;
        RECT 0.555000 1.495000 0.895000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.135000  0.085000 0.385000 0.655000 ;
      RECT 0.135000  1.495000 0.380000 2.635000 ;
      RECT 0.975000  0.085000 1.355000 0.485000 ;
      RECT 0.975000  0.655000 2.070000 0.825000 ;
      RECT 0.975000  0.825000 1.145000 1.325000 ;
      RECT 1.075000  1.495000 1.325000 2.635000 ;
      RECT 1.895000  0.255000 2.580000 0.620000 ;
      RECT 1.895000  0.620000 2.070000 0.655000 ;
      RECT 1.900000  0.825000 2.070000 1.955000 ;
      RECT 1.900000  1.955000 3.345000 2.125000 ;
      RECT 3.710000  0.085000 4.225000 0.525000 ;
      RECT 3.785000  0.695000 4.845000 0.865000 ;
      RECT 3.785000  0.865000 3.955000 1.185000 ;
      RECT 4.045000  1.835000 4.275000 2.635000 ;
      RECT 4.445000  1.835000 4.845000 2.465000 ;
      RECT 4.495000  0.255000 4.740000 0.695000 ;
      RECT 4.675000  0.865000 4.845000 1.835000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkmux2_2


MACRO sky130_fd_sc_hdll__nor4b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 1.340000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.075000 2.650000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.860000 1.075000 3.660000 1.285000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.205000 1.075000 5.885000 1.285000 ;
        RECT 5.615000 1.285000 5.885000 1.955000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.219500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.895000 0.725000 ;
        RECT 0.515000 0.725000 4.270000 0.905000 ;
        RECT 1.455000 0.255000 1.835000 0.725000 ;
        RECT 2.950000 0.255000 3.330000 0.725000 ;
        RECT 3.890000 0.255000 4.270000 0.725000 ;
        RECT 3.980000 1.455000 4.490000 1.625000 ;
        RECT 3.980000 1.625000 4.230000 2.125000 ;
        RECT 4.065000 0.905000 4.270000 1.075000 ;
        RECT 4.065000 1.075000 4.490000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.905000 ;
      RECT 0.085000  1.455000 2.305000 1.625000 ;
      RECT 0.085000  1.625000 0.425000 2.465000 ;
      RECT 0.645000  1.795000 0.855000 2.635000 ;
      RECT 1.075000  1.625000 1.325000 2.465000 ;
      RECT 1.115000  0.085000 1.285000 0.555000 ;
      RECT 1.545000  1.795000 1.755000 2.295000 ;
      RECT 1.545000  2.295000 3.290000 2.465000 ;
      RECT 1.925000  1.625000 2.305000 2.125000 ;
      RECT 2.055000  0.085000 2.780000 0.555000 ;
      RECT 2.475000  1.455000 3.760000 1.625000 ;
      RECT 2.475000  1.625000 2.860000 2.125000 ;
      RECT 3.080000  1.795000 3.290000 2.295000 ;
      RECT 3.510000  1.625000 3.760000 2.295000 ;
      RECT 3.510000  2.295000 4.695000 2.465000 ;
      RECT 3.550000  0.085000 3.720000 0.555000 ;
      RECT 4.450000  1.795000 4.695000 2.295000 ;
      RECT 4.490000  0.085000 4.695000 0.895000 ;
      RECT 4.720000  1.075000 5.035000 1.245000 ;
      RECT 4.865000  0.380000 5.220000 0.905000 ;
      RECT 4.865000  0.905000 5.035000 1.075000 ;
      RECT 4.865000  1.245000 5.035000 2.035000 ;
      RECT 4.865000  2.035000 5.220000 2.450000 ;
      RECT 5.440000  0.085000 5.690000 0.825000 ;
      RECT 5.440000  2.135000 5.690000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4b_2


MACRO sky130_fd_sc_hdll__nor4b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.660000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 1.075000 2.005000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275000 1.075000 4.150000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.385000 1.075000 6.285000 1.285000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855000 1.075000 9.550000 1.285000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  2.341500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.895000 0.725000 ;
        RECT 0.515000 0.725000 7.995000 0.905000 ;
        RECT 1.455000 0.255000 1.835000 0.725000 ;
        RECT 2.395000 0.255000 2.775000 0.725000 ;
        RECT 3.335000 0.255000 3.715000 0.725000 ;
        RECT 4.795000 0.255000 5.175000 0.725000 ;
        RECT 5.735000 0.255000 6.115000 0.725000 ;
        RECT 6.675000 0.255000 7.055000 0.725000 ;
        RECT 6.765000 0.905000 7.250000 1.455000 ;
        RECT 6.765000 1.455000 7.955000 1.625000 ;
        RECT 6.765000 1.625000 7.015000 2.125000 ;
        RECT 7.615000 0.255000 7.995000 0.725000 ;
        RECT 7.705000 1.625000 7.955000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.095000  1.455000 2.265000 1.625000 ;
      RECT 0.095000  1.625000 0.425000 2.465000 ;
      RECT 0.175000  0.085000 0.345000 0.895000 ;
      RECT 0.645000  1.795000 0.855000 2.635000 ;
      RECT 1.075000  1.625000 1.325000 2.465000 ;
      RECT 1.115000  0.085000 1.285000 0.555000 ;
      RECT 1.545000  1.795000 1.795000 2.635000 ;
      RECT 2.015000  1.625000 2.265000 2.295000 ;
      RECT 2.015000  2.295000 4.145000 2.465000 ;
      RECT 2.055000  0.085000 2.225000 0.555000 ;
      RECT 2.485000  1.455000 6.075000 1.625000 ;
      RECT 2.485000  1.625000 2.735000 2.125000 ;
      RECT 2.955000  1.795000 3.205000 2.295000 ;
      RECT 2.995000  0.085000 3.165000 0.555000 ;
      RECT 3.425000  1.625000 3.675000 2.125000 ;
      RECT 3.895000  1.795000 4.145000 2.295000 ;
      RECT 3.935000  0.085000 4.625000 0.555000 ;
      RECT 4.415000  1.795000 4.665000 2.295000 ;
      RECT 4.415000  2.295000 8.425000 2.465000 ;
      RECT 4.885000  1.625000 5.135000 2.125000 ;
      RECT 5.355000  1.795000 5.605000 2.295000 ;
      RECT 5.395000  0.085000 5.565000 0.555000 ;
      RECT 5.825000  1.625000 6.075000 2.125000 ;
      RECT 6.295000  1.455000 6.545000 2.295000 ;
      RECT 6.335000  0.085000 6.505000 0.555000 ;
      RECT 7.235000  1.795000 7.485000 2.295000 ;
      RECT 7.275000  0.085000 7.445000 0.555000 ;
      RECT 7.420000  1.075000 8.440000 1.285000 ;
      RECT 8.175000  1.795000 8.425000 2.295000 ;
      RECT 8.215000  0.085000 8.385000 0.555000 ;
      RECT 8.270000  0.735000 8.985000 0.905000 ;
      RECT 8.270000  0.905000 8.440000 1.075000 ;
      RECT 8.270000  1.285000 8.440000 1.455000 ;
      RECT 8.270000  1.455000 8.985000 1.625000 ;
      RECT 8.610000  0.255000 8.985000 0.735000 ;
      RECT 8.650000  1.625000 8.985000 2.465000 ;
      RECT 9.205000  0.085000 9.435000 0.905000 ;
      RECT 9.205000  1.455000 9.435000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4b_4


MACRO sky130_fd_sc_hdll__nor4b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.175000 0.995000 2.655000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 0.995000 1.935000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 0.995000 1.285000 1.615000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.825000 0.995000 3.225000 1.615000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.913500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.655000 2.075000 0.825000 ;
        RECT 0.085000 0.825000 0.345000 2.450000 ;
        RECT 0.905000 0.300000 1.105000 0.655000 ;
        RECT 1.875000 0.310000 2.075000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.355000  0.085000 0.685000 0.480000 ;
      RECT 0.525000  0.995000 0.745000 1.795000 ;
      RECT 0.525000  1.795000 3.565000 2.005000 ;
      RECT 1.325000  0.085000 1.655000 0.485000 ;
      RECT 2.245000  0.085000 2.735000 0.825000 ;
      RECT 2.325000  2.185000 2.705000 2.635000 ;
      RECT 3.090000  0.405000 3.260000 0.655000 ;
      RECT 3.090000  0.655000 3.565000 0.825000 ;
      RECT 3.395000  0.825000 3.565000 1.795000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4b_1


MACRO sky130_fd_sc_hdll__conb_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  1.380000 BY  2.720000 ;
  SITE unithd ;
  PIN HI
    ANTENNADIFFAREA  0.000000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.605000 1.740000 ;
    END
  END HI
  PIN LO
    ANTENNADIFFAREA  0.000000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.775000 0.915000 1.295000 2.465000 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.275000  1.910000 0.605000 2.635000 ;
      RECT 0.775000  0.085000 1.115000 0.745000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__conb_1


MACRO sky130_fd_sc_hdll__buf_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  1.840000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.220200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.985000 0.545000 1.355000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.348500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.255000 1.395000 0.760000 ;
        RECT 1.065000 1.560000 1.395000 2.465000 ;
        RECT 1.215000 0.760000 1.395000 1.560000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 1.840000 0.085000 ;
        RECT 0.525000  0.085000 0.895000 0.465000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 1.840000 2.805000 ;
        RECT 0.525000 1.875000 0.895000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.165000 1.535000 0.890000 1.705000 ;
      RECT 0.165000 1.705000 0.345000 2.465000 ;
      RECT 0.175000 0.255000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 0.890000 0.805000 ;
      RECT 0.720000 0.805000 0.890000 1.060000 ;
      RECT 0.720000 1.060000 1.035000 1.390000 ;
      RECT 0.720000 1.390000 0.890000 1.535000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_1


MACRO sky130_fd_sc_hdll__buf_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.832500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.340000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055000 0.255000 2.225000 0.735000 ;
        RECT 2.055000 0.735000 5.045000 0.905000 ;
        RECT 2.055000 1.445000 5.045000 1.615000 ;
        RECT 2.055000 1.615000 2.225000 2.465000 ;
        RECT 2.995000 0.255000 3.165000 0.735000 ;
        RECT 2.995000 1.615000 3.165000 2.465000 ;
        RECT 3.935000 0.255000 4.105000 0.735000 ;
        RECT 3.935000 1.615000 4.105000 2.465000 ;
        RECT 4.690000 0.905000 5.045000 1.445000 ;
        RECT 4.875000 0.255000 5.045000 0.735000 ;
        RECT 4.875000 1.615000 5.045000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.515000  0.085000 0.895000 0.565000 ;
        RECT 1.455000  0.085000 1.835000 0.565000 ;
        RECT 2.395000  0.085000 2.775000 0.565000 ;
        RECT 3.335000  0.085000 3.715000 0.565000 ;
        RECT 4.275000  0.085000 4.655000 0.565000 ;
        RECT 5.215000  0.085000 5.595000 0.885000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.645000 1.835000 0.815000 2.635000 ;
        RECT 1.585000 1.835000 1.755000 2.635000 ;
        RECT 2.395000 1.835000 2.775000 2.635000 ;
        RECT 3.335000 1.835000 3.715000 2.635000 ;
        RECT 4.275000 1.835000 4.655000 2.635000 ;
        RECT 5.215000 1.485000 5.595000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 1.445000 1.745000 1.615000 ;
      RECT 0.095000 1.615000 0.425000 2.465000 ;
      RECT 0.175000 0.255000 0.345000 0.735000 ;
      RECT 0.175000 0.735000 1.745000 0.905000 ;
      RECT 0.985000 1.615000 1.365000 2.465000 ;
      RECT 1.115000 0.260000 1.285000 0.735000 ;
      RECT 1.570000 0.905000 1.745000 1.075000 ;
      RECT 1.570000 1.075000 4.495000 1.245000 ;
      RECT 1.570000 1.245000 1.745000 1.445000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_8


MACRO sky130_fd_sc_hdll__buf_16
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.50000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 2.735000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  4.016500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  3.335000 0.255000  3.635000 0.260000 ;
        RECT  3.335000 0.260000  3.715000 0.735000 ;
        RECT  3.335000 0.735000 11.135000 0.905000 ;
        RECT  3.335000 1.445000 11.135000 1.615000 ;
        RECT  3.335000 1.615000  3.715000 2.465000 ;
        RECT  4.275000 0.260000  4.655000 0.735000 ;
        RECT  4.275000 1.615000  4.655000 2.465000 ;
        RECT  4.405000 0.255000  4.575000 0.260000 ;
        RECT  5.215000 0.260000  5.595000 0.735000 ;
        RECT  5.215000 1.615000  5.595000 2.465000 ;
        RECT  5.345000 0.255000  5.515000 0.260000 ;
        RECT  6.155000 0.260000  6.535000 0.735000 ;
        RECT  6.155000 1.615000  6.535000 2.465000 ;
        RECT  7.095000 0.260000  7.475000 0.735000 ;
        RECT  7.095000 1.615000  7.475000 2.465000 ;
        RECT  8.035000 0.260000  8.415000 0.735000 ;
        RECT  8.035000 1.615000  8.415000 2.465000 ;
        RECT  8.975000 0.260000  9.355000 0.735000 ;
        RECT  8.975000 1.615000  9.355000 2.465000 ;
        RECT  9.915000 0.260000 10.295000 0.735000 ;
        RECT  9.915000 1.615000 10.295000 2.465000 ;
        RECT 10.635000 0.905000 11.135000 1.445000 ;
        RECT 10.860000 0.365000 11.135000 0.735000 ;
        RECT 10.860000 1.615000 11.135000 2.360000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.500000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.500000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.500000 0.085000 ;
      RECT  0.000000  2.635000 11.500000 2.805000 ;
      RECT  0.175000  0.085000  0.345000 0.905000 ;
      RECT  0.175000  1.445000  0.345000 2.635000 ;
      RECT  0.515000  0.260000  0.895000 0.735000 ;
      RECT  0.515000  0.735000  3.165000 0.905000 ;
      RECT  0.515000  1.445000  3.165000 1.615000 ;
      RECT  0.515000  1.615000  0.895000 2.465000 ;
      RECT  1.115000  0.085000  1.285000 0.565000 ;
      RECT  1.115000  1.835000  1.285000 2.635000 ;
      RECT  1.455000  0.260000  1.835000 0.735000 ;
      RECT  1.455000  1.615000  1.835000 2.465000 ;
      RECT  2.055000  0.085000  2.225000 0.565000 ;
      RECT  2.055000  1.835000  2.225000 2.635000 ;
      RECT  2.395000  0.260000  2.775000 0.735000 ;
      RECT  2.395000  1.615000  2.775000 2.465000 ;
      RECT  2.990000  0.905000  3.165000 1.075000 ;
      RECT  2.990000  1.075000 10.175000 1.275000 ;
      RECT  2.990000  1.275000  3.165000 1.445000 ;
      RECT  2.995000  0.085000  3.165000 0.565000 ;
      RECT  2.995000  1.835000  3.165000 2.635000 ;
      RECT  3.935000  0.085000  4.105000 0.565000 ;
      RECT  3.935000  1.835000  4.105000 2.635000 ;
      RECT  4.875000  0.085000  5.045000 0.565000 ;
      RECT  4.875000  1.835000  5.045000 2.635000 ;
      RECT  5.815000  0.085000  5.985000 0.565000 ;
      RECT  5.815000  1.835000  5.985000 2.635000 ;
      RECT  6.755000  0.085000  6.925000 0.565000 ;
      RECT  6.755000  1.835000  6.925000 2.635000 ;
      RECT  7.695000  0.085000  7.865000 0.565000 ;
      RECT  7.695000  1.835000  7.865000 2.635000 ;
      RECT  8.635000  0.085000  8.805000 0.565000 ;
      RECT  8.635000  1.835000  8.805000 2.635000 ;
      RECT  9.575000  0.085000  9.745000 0.565000 ;
      RECT  9.575000  1.835000  9.745000 2.635000 ;
      RECT 10.515000  0.085000 10.685000 0.565000 ;
      RECT 10.515000  1.835000 10.685000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_16


MACRO sky130_fd_sc_hdll__buf_12
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.280000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 1.075000 1.810000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.020500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 0.255000 2.695000 0.735000 ;
        RECT 2.525000 0.735000 7.395000 0.905000 ;
        RECT 2.525000 1.445000 7.395000 1.615000 ;
        RECT 2.525000 1.615000 2.695000 2.465000 ;
        RECT 3.465000 0.255000 3.635000 0.735000 ;
        RECT 3.465000 1.615000 3.635000 2.465000 ;
        RECT 4.405000 0.255000 4.575000 0.735000 ;
        RECT 4.405000 1.615000 4.575000 2.465000 ;
        RECT 5.210000 0.905000 7.395000 1.445000 ;
        RECT 5.345000 0.255000 5.515000 0.735000 ;
        RECT 5.345000 1.615000 5.515000 2.465000 ;
        RECT 6.285000 0.255000 6.455000 0.735000 ;
        RECT 6.285000 1.615000 6.455000 2.465000 ;
        RECT 7.225000 0.255000 7.395000 0.735000 ;
        RECT 7.225000 1.615000 7.395000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.280000 0.085000 ;
        RECT 0.095000  0.085000 0.425000 0.565000 ;
        RECT 0.985000  0.085000 1.365000 0.565000 ;
        RECT 1.925000  0.085000 2.305000 0.565000 ;
        RECT 2.865000  0.085000 3.245000 0.565000 ;
        RECT 3.805000  0.085000 4.185000 0.565000 ;
        RECT 4.745000  0.085000 5.125000 0.565000 ;
        RECT 5.685000  0.085000 6.065000 0.565000 ;
        RECT 6.625000  0.085000 7.005000 0.565000 ;
        RECT 7.565000  0.085000 7.945000 0.885000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.280000 2.805000 ;
        RECT 0.175000 1.835000 0.345000 2.635000 ;
        RECT 1.115000 1.835000 1.285000 2.635000 ;
        RECT 2.055000 1.835000 2.225000 2.635000 ;
        RECT 2.865000 1.835000 3.245000 2.635000 ;
        RECT 3.805000 1.835000 4.185000 2.635000 ;
        RECT 4.745000 1.835000 5.125000 2.635000 ;
        RECT 5.685000 1.835000 6.065000 2.635000 ;
        RECT 6.625000 1.835000 7.005000 2.635000 ;
        RECT 7.565000 1.485000 7.945000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515000 1.445000 2.215000 1.615000 ;
      RECT 0.515000 1.615000 0.895000 2.465000 ;
      RECT 0.645000 0.255000 0.815000 0.735000 ;
      RECT 0.645000 0.735000 2.215000 0.905000 ;
      RECT 1.455000 1.615000 1.835000 2.465000 ;
      RECT 1.585000 0.260000 1.755000 0.735000 ;
      RECT 2.040000 0.905000 2.215000 1.075000 ;
      RECT 2.040000 1.075000 4.965000 1.245000 ;
      RECT 2.040000 1.245000 2.215000 1.445000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_12


MACRO sky130_fd_sc_hdll__buf_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.470000 1.315000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 0.255000 1.285000 0.735000 ;
        RECT 1.115000 0.735000 2.225000 0.905000 ;
        RECT 1.115000 1.445000 2.225000 1.615000 ;
        RECT 1.115000 1.615000 1.285000 2.465000 ;
        RECT 1.920000 0.905000 2.225000 1.445000 ;
        RECT 2.055000 0.255000 2.225000 0.735000 ;
        RECT 2.055000 1.615000 2.225000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.220000 0.085000 ;
        RECT 0.525000  0.085000 0.815000 0.565000 ;
        RECT 1.455000  0.085000 1.835000 0.565000 ;
        RECT 2.395000  0.085000 2.775000 0.885000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.220000 2.805000 ;
        RECT 0.645000 1.835000 0.885000 2.635000 ;
        RECT 1.455000 1.835000 1.835000 2.635000 ;
        RECT 2.395000 1.485000 2.775000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 1.485000 0.860000 1.655000 ;
      RECT 0.095000 1.655000 0.425000 2.465000 ;
      RECT 0.175000 0.255000 0.345000 0.735000 ;
      RECT 0.175000 0.735000 0.860000 0.905000 ;
      RECT 0.690000 0.905000 0.860000 1.075000 ;
      RECT 0.690000 1.075000 1.240000 1.245000 ;
      RECT 0.690000 1.245000 0.860000 1.485000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_4


MACRO sky130_fd_sc_hdll__buf_6
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.280000 1.075000 1.265000 1.315000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.526500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845000 0.255000 2.015000 0.735000 ;
        RECT 1.845000 0.735000 3.895000 0.905000 ;
        RECT 1.845000 1.445000 3.895000 1.615000 ;
        RECT 1.845000 1.615000 2.015000 2.465000 ;
        RECT 2.410000 0.905000 3.895000 1.445000 ;
        RECT 2.785000 0.255000 2.955000 0.735000 ;
        RECT 2.785000 1.615000 2.955000 2.465000 ;
        RECT 3.725000 0.255000 3.895000 0.735000 ;
        RECT 3.725000 1.615000 3.895000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.600000 0.085000 ;
        RECT 0.435000  0.085000 0.605000 0.565000 ;
        RECT 1.375000  0.085000 1.545000 0.565000 ;
        RECT 2.185000  0.085000 2.565000 0.565000 ;
        RECT 3.125000  0.085000 3.505000 0.565000 ;
        RECT 4.065000  0.085000 4.445000 0.885000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.600000 2.805000 ;
        RECT 0.435000 1.485000 0.605000 2.635000 ;
        RECT 1.375000 1.835000 1.615000 2.635000 ;
        RECT 2.185000 1.835000 2.565000 2.635000 ;
        RECT 3.125000 1.835000 3.505000 2.635000 ;
        RECT 4.065000 1.485000 4.445000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.775000 0.255000 1.155000 0.735000 ;
      RECT 0.775000 0.735000 1.625000 0.905000 ;
      RECT 0.775000 1.485000 1.625000 1.655000 ;
      RECT 0.775000 1.655000 1.155000 2.465000 ;
      RECT 1.455000 0.905000 1.625000 1.075000 ;
      RECT 1.455000 1.075000 1.975000 1.245000 ;
      RECT 1.455000 1.245000 1.625000 1.485000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_6


MACRO sky130_fd_sc_hdll__buf_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.440000 1.355000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.703800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.270000 0.255000 1.695000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 2.300000 0.085000 ;
        RECT 0.610000  0.085000 0.940000 0.465000 ;
        RECT 1.865000  0.085000 2.125000 0.925000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 2.300000 2.805000 ;
        RECT 0.600000 1.875000 0.930000 2.635000 ;
        RECT 1.865000 1.485000 2.125000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.255000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 0.940000 0.805000 ;
      RECT 0.175000 1.535000 0.895000 1.705000 ;
      RECT 0.175000 1.705000 0.345000 2.465000 ;
      RECT 0.725000 0.805000 0.940000 0.995000 ;
      RECT 0.725000 0.995000 1.025000 1.325000 ;
      RECT 0.725000 1.325000 0.895000 1.535000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__buf_2


MACRO sky130_fd_sc_hdll__inputiso0n_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 0.590000 1.325000 ;
        RECT 0.100000 1.325000 0.365000 1.685000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 1.075000 1.275000 1.325000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.539000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595000 0.255000 2.205000 0.545000 ;
        RECT 1.745000 1.915000 2.205000 2.465000 ;
        RECT 1.955000 0.545000 2.205000 1.915000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.125000  0.355000 0.455000 0.715000 ;
      RECT 0.125000  0.715000 1.695000 0.905000 ;
      RECT 0.125000  1.965000 0.405000 2.635000 ;
      RECT 0.625000  1.575000 1.695000 1.745000 ;
      RECT 0.625000  1.745000 0.925000 2.295000 ;
      RECT 1.175000  0.085000 1.425000 0.545000 ;
      RECT 1.175000  1.915000 1.505000 2.635000 ;
      RECT 1.525000  0.905000 1.695000 1.575000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inputiso0n_1


MACRO sky130_fd_sc_hdll__o211ai_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 1.075000 4.915000 1.295000 ;
        RECT 4.465000 0.765000 4.915000 1.075000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.670000 1.075000 3.635000 1.355000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.215000 1.075000 2.210000 1.365000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.375000 1.970000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.114500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.670000 0.925000 1.540000 ;
        RECT 0.545000 1.540000 3.405000 1.710000 ;
        RECT 0.545000 1.710000 0.855000 2.465000 ;
        RECT 1.625000 1.710000 1.815000 2.465000 ;
        RECT 3.025000 1.710000 3.405000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.095000  0.255000 2.365000 0.445000 ;
      RECT 0.115000  2.175000 0.375000 2.635000 ;
      RECT 1.025000  1.915000 1.405000 2.635000 ;
      RECT 1.145000  0.445000 2.365000 0.465000 ;
      RECT 1.145000  0.465000 1.335000 0.890000 ;
      RECT 1.505000  0.635000 4.295000 0.845000 ;
      RECT 1.985000  1.915000 2.365000 2.635000 ;
      RECT 2.595000  0.085000 2.925000 0.445000 ;
      RECT 2.595000  2.100000 2.855000 2.295000 ;
      RECT 2.595000  2.295000 3.815000 2.465000 ;
      RECT 3.525000  0.085000 3.905000 0.445000 ;
      RECT 3.625000  1.525000 4.845000 1.695000 ;
      RECT 3.625000  1.695000 3.815000 2.295000 ;
      RECT 3.985000  1.865000 4.365000 2.635000 ;
      RECT 4.105000  0.515000 4.295000 0.635000 ;
      RECT 4.465000  0.085000 4.870000 0.445000 ;
      RECT 4.585000  1.695000 4.845000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211ai_2


MACRO sky130_fd_sc_hdll__o211ai_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.395000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 0.995000 1.080000 1.325000 ;
        RECT 0.565000 1.325000 0.825000 2.250000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 0.995000 1.745000 1.345000 ;
        RECT 1.495000 1.345000 1.745000 1.615000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.915000 1.020000 2.270000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.297000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.595000 1.325000 1.815000 ;
        RECT 0.995000 1.815000 2.675000 2.045000 ;
        RECT 0.995000 2.045000 1.325000 2.445000 ;
        RECT 1.725000 0.255000 2.675000 0.825000 ;
        RECT 2.075000 2.045000 2.675000 2.465000 ;
        RECT 2.440000 0.825000 2.675000 1.815000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  0.255000 0.400000 0.615000 ;
      RECT 0.095000  0.615000 1.450000 0.825000 ;
      RECT 0.095000  1.495000 0.395000 2.635000 ;
      RECT 0.570000  0.085000 0.900000 0.445000 ;
      RECT 1.070000  0.255000 1.450000 0.615000 ;
      RECT 1.540000  2.275000 1.870000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.590000 2.805000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211ai_1


MACRO sky130_fd_sc_hdll__o211ai_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.740000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.400000 1.075000 1.560000 1.330000 ;
        RECT 1.015000 1.330000 1.560000 1.515000 ;
        RECT 1.015000 1.515000 4.030000 1.685000 ;
        RECT 3.700000 0.995000 4.030000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.855000 1.075000 3.530000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.200000 0.995000 5.525000 1.410000 ;
        RECT 4.710000 1.410000 5.525000 1.515000 ;
        RECT 4.710000 1.515000 7.800000 1.685000 ;
        RECT 7.580000 0.995000 7.800000 1.515000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.970000 1.075000 7.140000 1.345000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.218500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 1.855000 8.480000 2.025000 ;
        RECT 1.955000 2.025000 3.820000 2.105000 ;
        RECT 4.495000 2.025000 8.480000 2.105000 ;
        RECT 5.830000 0.270000 7.485000 0.450000 ;
        RECT 7.265000 0.450000 7.485000 0.655000 ;
        RECT 7.265000 0.655000 8.160000 0.825000 ;
        RECT 7.980000 0.825000 8.160000 1.340000 ;
        RECT 7.980000 1.340000 8.480000 1.855000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.090000  1.665000 0.385000 2.635000 ;
      RECT 0.155000  0.535000 0.355000 0.625000 ;
      RECT 0.155000  0.625000 4.235000 0.795000 ;
      RECT 0.155000  0.795000 3.480000 0.905000 ;
      RECT 0.525000  0.085000 0.905000 0.445000 ;
      RECT 0.605000  1.860000 0.825000 1.935000 ;
      RECT 0.605000  1.935000 1.785000 2.105000 ;
      RECT 0.605000  2.105000 0.825000 2.190000 ;
      RECT 1.005000  2.275000 1.385000 2.635000 ;
      RECT 1.125000  0.425000 1.340000 0.625000 ;
      RECT 1.535000  0.085000 1.865000 0.455000 ;
      RECT 1.605000  2.105000 1.785000 2.275000 ;
      RECT 1.605000  2.275000 3.785000 2.465000 ;
      RECT 2.445000  0.085000 2.825000 0.445000 ;
      RECT 3.405000  0.085000 3.785000 0.445000 ;
      RECT 4.005000  0.255000 5.470000 0.455000 ;
      RECT 4.005000  0.455000 4.235000 0.625000 ;
      RECT 4.015000  2.195000 4.285000 2.635000 ;
      RECT 4.405000  0.635000 6.870000 0.815000 ;
      RECT 4.885000  2.275000 5.265000 2.635000 ;
      RECT 5.830000  2.275000 6.210000 2.635000 ;
      RECT 6.770000  2.275000 7.155000 2.635000 ;
      RECT 7.730000  0.310000 8.490000 0.480000 ;
      RECT 8.155000  2.275000 8.485000 2.635000 ;
      RECT 8.320000  0.480000 8.490000 0.595000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.170000  0.425000 1.340000 0.595000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.320000  0.425000 8.490000 0.595000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
    LAYER met1 ;
      RECT 1.110000 0.395000 1.400000 0.440000 ;
      RECT 1.110000 0.440000 8.550000 0.580000 ;
      RECT 1.110000 0.580000 1.400000 0.625000 ;
      RECT 8.260000 0.395000 8.550000 0.440000 ;
      RECT 8.260000 0.580000 8.550000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211ai_4


MACRO sky130_fd_sc_hdll__o21ba_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.540000 1.075000 6.355000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.180000 1.075000 5.320000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 0.935000 1.285000 ;
        RECT 0.605000 1.285000 0.935000 1.705000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.155000 0.255000 1.485000 0.725000 ;
        RECT 1.155000 0.725000 2.375000 0.910000 ;
        RECT 1.155000 0.910000 1.705000 1.445000 ;
        RECT 1.155000 1.445000 2.425000 1.705000 ;
        RECT 2.045000 0.255000 2.375000 0.725000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  0.265000 0.545000 0.855000 ;
      RECT 0.085000  0.855000 0.255000 1.455000 ;
      RECT 0.085000  1.455000 0.435000 1.875000 ;
      RECT 0.085000  1.875000 2.815000 2.045000 ;
      RECT 0.085000  2.045000 0.435000 2.465000 ;
      RECT 0.635000  2.215000 1.015000 2.635000 ;
      RECT 0.765000  0.085000 0.935000 0.905000 ;
      RECT 1.575000  2.215000 1.955000 2.635000 ;
      RECT 1.705000  0.085000 1.875000 0.555000 ;
      RECT 1.875000  1.080000 2.815000 1.250000 ;
      RECT 2.515000  2.215000 2.895000 2.635000 ;
      RECT 2.565000  0.085000 2.895000 0.475000 ;
      RECT 2.645000  0.645000 3.935000 0.895000 ;
      RECT 2.645000  0.895000 2.815000 1.080000 ;
      RECT 2.645000  1.445000 3.205000 1.615000 ;
      RECT 2.645000  1.615000 2.815000 1.875000 ;
      RECT 2.985000  1.075000 3.435000 1.245000 ;
      RECT 2.985000  1.245000 3.205000 1.445000 ;
      RECT 3.105000  0.255000 4.405000 0.475000 ;
      RECT 3.115000  1.795000 4.830000 1.965000 ;
      RECT 3.115000  1.965000 3.285000 2.465000 ;
      RECT 3.550000  2.135000 3.800000 2.635000 ;
      RECT 3.745000  0.895000 3.935000 1.795000 ;
      RECT 4.035000  2.135000 4.325000 2.295000 ;
      RECT 4.035000  2.295000 5.265000 2.465000 ;
      RECT 4.155000  0.475000 4.405000 0.725000 ;
      RECT 4.155000  0.725000 6.310000 0.905000 ;
      RECT 4.585000  1.445000 4.830000 1.795000 ;
      RECT 4.585000  1.965000 4.830000 2.125000 ;
      RECT 4.625000  0.085000 4.795000 0.555000 ;
      RECT 4.965000  0.255000 5.345000 0.725000 ;
      RECT 5.095000  1.455000 6.310000 1.665000 ;
      RECT 5.095000  1.665000 5.265000 2.295000 ;
      RECT 5.435000  1.835000 5.815000 2.635000 ;
      RECT 5.565000  0.085000 5.735000 0.555000 ;
      RECT 5.905000  0.265000 6.310000 0.725000 ;
      RECT 6.035000  1.665000 6.310000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ba_4


MACRO sky130_fd_sc_hdll__o21ba_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 1.075000 3.895000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.645000 1.075000 3.180000 1.285000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.825000 1.325000 ;
        RECT 0.605000 1.325000 0.825000 1.695000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.571700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 0.295000 1.380000 0.465000 ;
        RECT 0.995000 0.465000 1.235000 1.495000 ;
        RECT 0.995000 1.495000 1.455000 1.695000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.430000 0.345000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 0.395000 1.865000 ;
      RECT 0.085000  1.865000 2.085000 2.035000 ;
      RECT 0.520000  2.205000 0.960000 2.635000 ;
      RECT 0.645000  0.085000 0.825000 0.825000 ;
      RECT 1.405000  0.655000 2.470000 0.825000 ;
      RECT 1.405000  0.825000 1.575000 1.325000 ;
      RECT 1.520000  2.205000 2.380000 2.635000 ;
      RECT 1.560000  0.085000 1.925000 0.465000 ;
      RECT 1.915000  0.995000 2.085000 1.865000 ;
      RECT 2.140000  0.255000 2.470000 0.655000 ;
      RECT 2.255000  0.825000 2.470000 1.455000 ;
      RECT 2.255000  1.455000 2.925000 2.035000 ;
      RECT 2.600000  2.035000 2.925000 2.465000 ;
      RECT 2.695000  0.365000 2.945000 0.735000 ;
      RECT 2.695000  0.735000 3.890000 0.905000 ;
      RECT 3.165000  0.085000 3.335000 0.555000 ;
      RECT 3.450000  1.875000 3.830000 2.635000 ;
      RECT 3.555000  0.270000 3.890000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ba_2


MACRO sky130_fd_sc_hdll__o21ba_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.020000 1.075000 3.570000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.230000 1.075000 2.850000 1.285000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 0.995000 1.380000 1.325000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.450000 0.445000 0.825000 ;
        RECT 0.085000 0.825000 0.340000 1.480000 ;
        RECT 0.085000 1.480000 0.425000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.510000  0.995000 0.860000 1.325000 ;
      RECT 0.595000  2.205000 1.005000 2.635000 ;
      RECT 0.645000  1.325000 0.860000 1.865000 ;
      RECT 0.645000  1.865000 2.585000 2.035000 ;
      RECT 0.675000  0.085000 0.845000 0.825000 ;
      RECT 1.075000  1.525000 1.720000 1.695000 ;
      RECT 1.210000  0.450000 1.380000 0.655000 ;
      RECT 1.210000  0.655000 1.720000 0.825000 ;
      RECT 1.550000  0.825000 1.720000 1.525000 ;
      RECT 1.770000  2.215000 2.100000 2.635000 ;
      RECT 1.890000  0.255000 2.060000 1.455000 ;
      RECT 1.890000  1.455000 2.585000 1.865000 ;
      RECT 2.280000  0.255000 2.610000 0.735000 ;
      RECT 2.280000  0.735000 3.565000 0.905000 ;
      RECT 2.280000  2.035000 2.585000 2.465000 ;
      RECT 2.830000  0.085000 3.000000 0.555000 ;
      RECT 3.170000  1.535000 3.550000 2.635000 ;
      RECT 3.235000  0.270000 3.565000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ba_1


MACRO sky130_fd_sc_hdll__tapvpwrvgnd_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE WELLTAP ;
  SYMMETRY X Y R90 ;
  SIZE  0.460000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  1.470000 0.375000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__tapvpwrvgnd_1


MACRO sky130_fd_sc_hdll__or4_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 0.995000 2.210000 1.445000 ;
        RECT 1.940000 1.445000 2.475000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.380000 0.995000 1.760000 1.450000 ;
        RECT 1.500000 1.450000 1.760000 1.785000 ;
        RECT 1.500000 1.785000 1.870000 2.375000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.930000 0.995000 1.100000 1.620000 ;
        RECT 0.930000 1.620000 1.330000 2.375000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.755000 0.370000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.730000 1.455000 4.485000 1.625000 ;
        RECT 2.730000 1.625000 2.980000 2.465000 ;
        RECT 2.770000 0.255000 3.020000 0.725000 ;
        RECT 2.770000 0.725000 4.485000 0.905000 ;
        RECT 3.580000 0.255000 3.960000 0.725000 ;
        RECT 3.670000 1.625000 3.920000 2.465000 ;
        RECT 4.210000 0.905000 4.485000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.115000  1.495000 0.760000 1.665000 ;
      RECT 0.115000  1.665000 0.450000 2.450000 ;
      RECT 0.120000  0.085000 0.370000 0.585000 ;
      RECT 0.540000  0.655000 2.550000 0.825000 ;
      RECT 0.540000  0.825000 0.760000 1.495000 ;
      RECT 0.750000  0.305000 0.920000 0.655000 ;
      RECT 1.120000  0.085000 1.500000 0.485000 ;
      RECT 1.720000  0.305000 1.890000 0.655000 ;
      RECT 2.160000  0.085000 2.540000 0.485000 ;
      RECT 2.205000  1.795000 2.455000 2.635000 ;
      RECT 2.380000  0.825000 2.550000 1.075000 ;
      RECT 2.380000  1.075000 3.990000 1.245000 ;
      RECT 3.200000  1.795000 3.450000 2.635000 ;
      RECT 3.240000  0.085000 3.410000 0.555000 ;
      RECT 4.140000  1.795000 4.390000 2.635000 ;
      RECT 4.180000  0.085000 4.350000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4_4


MACRO sky130_fd_sc_hdll__or4_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 2.095000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 2.125000 1.895000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.660000 0.995000 1.355000 1.615000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.755000 0.440000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.703000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.805000 0.415000 3.075000 0.760000 ;
        RECT 2.805000 1.495000 3.075000 2.465000 ;
        RECT 2.905000 0.760000 3.075000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  1.495000 0.410000 1.785000 ;
      RECT 0.090000  1.785000 1.830000 1.955000 ;
      RECT 0.095000  0.085000 0.425000 0.585000 ;
      RECT 0.675000  0.305000 0.845000 0.655000 ;
      RECT 0.675000  0.655000 2.435000 0.825000 ;
      RECT 1.045000  0.085000 1.425000 0.485000 ;
      RECT 1.645000  0.305000 1.815000 0.655000 ;
      RECT 1.660000  1.495000 2.435000 1.665000 ;
      RECT 1.660000  1.665000 1.830000 1.785000 ;
      RECT 1.985000  0.085000 2.415000 0.485000 ;
      RECT 2.115000  1.835000 2.395000 2.635000 ;
      RECT 2.265000  0.825000 2.435000 0.995000 ;
      RECT 2.265000  0.995000 2.555000 1.325000 ;
      RECT 2.265000  1.325000 2.435000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4_1


MACRO sky130_fd_sc_hdll__or4_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 0.995000 2.095000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 2.125000 1.895000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.995000 1.305000 1.615000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.755000 0.435000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.802800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.820000 0.415000 3.125000 0.760000 ;
        RECT 2.820000 1.495000 3.125000 2.465000 ;
        RECT 2.890000 0.760000 3.125000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  1.495000 0.410000 1.785000 ;
      RECT 0.085000  1.785000 1.830000 1.955000 ;
      RECT 0.090000  0.085000 0.425000 0.585000 ;
      RECT 0.675000  0.305000 0.845000 0.655000 ;
      RECT 0.675000  0.655000 2.435000 0.825000 ;
      RECT 1.045000  0.085000 1.425000 0.485000 ;
      RECT 1.645000  0.305000 1.815000 0.655000 ;
      RECT 1.660000  1.495000 2.435000 1.665000 ;
      RECT 1.660000  1.665000 1.830000 1.785000 ;
      RECT 1.985000  0.085000 2.415000 0.485000 ;
      RECT 2.115000  1.835000 2.395000 2.635000 ;
      RECT 2.265000  0.825000 2.435000 0.995000 ;
      RECT 2.265000  0.995000 2.700000 1.325000 ;
      RECT 2.265000  1.325000 2.435000 1.495000 ;
      RECT 3.315000  0.085000 3.535000 1.000000 ;
      RECT 3.315000  1.455000 3.535000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4_2


MACRO sky130_fd_sc_hdll__and4b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.450000 1.675000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.675000 0.420000 2.155000 1.695000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 0.420000 2.615000 1.695000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 0.665000 3.075000 1.695000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.520000 0.295000 3.995000 0.805000 ;
        RECT 3.635000 1.495000 3.995000 2.465000 ;
        RECT 3.725000 0.805000 3.995000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.170000  0.255000 0.345000 0.655000 ;
      RECT 0.170000  0.655000 0.850000 0.825000 ;
      RECT 0.170000  1.845000 0.850000 2.015000 ;
      RECT 0.170000  2.015000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.895000 0.465000 ;
      RECT 0.515000  2.195000 0.895000 2.635000 ;
      RECT 0.680000  0.825000 0.850000 0.995000 ;
      RECT 0.680000  0.995000 1.025000 1.325000 ;
      RECT 0.680000  1.325000 0.850000 1.845000 ;
      RECT 1.140000  0.255000 1.370000 0.585000 ;
      RECT 1.200000  0.585000 1.370000 1.875000 ;
      RECT 1.200000  1.875000 3.415000 2.045000 ;
      RECT 1.200000  2.045000 1.370000 2.465000 ;
      RECT 1.655000  2.225000 2.375000 2.635000 ;
      RECT 2.630000  2.045000 2.800000 2.465000 ;
      RECT 2.955000  0.085000 3.350000 0.465000 ;
      RECT 3.060000  2.225000 3.390000 2.635000 ;
      RECT 3.245000  0.995000 3.535000 1.325000 ;
      RECT 3.245000  1.325000 3.415000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4b_1


MACRO sky130_fd_sc_hdll__and4b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 0.765000 0.840000 1.635000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.810000 0.735000 4.190000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.330000 0.755000 3.640000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.870000 0.995000 3.120000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 0.255000 1.340000 0.650000 ;
        RECT 1.030000 0.650000 2.280000 0.820000 ;
        RECT 1.030000 0.820000 1.360000 1.545000 ;
        RECT 1.030000 1.545000 2.360000 1.715000 ;
        RECT 2.110000 0.255000 2.280000 0.650000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.260000 1.915000 ;
      RECT 0.085000  1.915000 4.885000 2.085000 ;
      RECT 0.085000  2.085000 0.345000 2.465000 ;
      RECT 0.515000  2.255000 0.895000 2.635000 ;
      RECT 0.565000  0.085000 0.815000 0.545000 ;
      RECT 1.510000  0.085000 1.890000 0.470000 ;
      RECT 1.510000  2.255000 1.890000 2.635000 ;
      RECT 1.530000  0.995000 2.700000 1.325000 ;
      RECT 2.450000  2.255000 2.830000 2.635000 ;
      RECT 2.530000  1.325000 2.700000 1.545000 ;
      RECT 2.530000  1.545000 4.530000 1.715000 ;
      RECT 2.535000  0.085000 2.865000 0.445000 ;
      RECT 3.510000  2.255000 3.890000 2.635000 ;
      RECT 4.360000  0.640000 4.900000 0.810000 ;
      RECT 4.360000  0.810000 4.530000 1.545000 ;
      RECT 4.570000  2.255000 4.950000 2.635000 ;
      RECT 4.715000  0.995000 4.885000 1.915000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4b_4


MACRO sky130_fd_sc_hdll__and4b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.740000 0.335000 1.630000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 0.420000 2.155000 1.745000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 0.420000 2.615000 1.615000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 0.645000 3.115000 1.615000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.555700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.560000 0.255000 3.895000 0.640000 ;
        RECT 3.560000 0.640000 4.455000 0.825000 ;
        RECT 3.690000 1.535000 4.455000 1.665000 ;
        RECT 3.690000 1.665000 3.995000 2.465000 ;
        RECT 3.775000 0.825000 4.455000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.175000  1.830000 0.855000 2.000000 ;
      RECT 0.175000  2.000000 0.345000 2.465000 ;
      RECT 0.515000  2.195000 0.895000 2.635000 ;
      RECT 0.645000  0.255000 0.855000 0.585000 ;
      RECT 0.685000  0.585000 0.855000 0.995000 ;
      RECT 0.685000  0.995000 1.075000 1.325000 ;
      RECT 0.685000  1.325000 0.855000 1.830000 ;
      RECT 1.115000  1.660000 1.415000 1.915000 ;
      RECT 1.115000  1.915000 3.465000 1.965000 ;
      RECT 1.115000  1.965000 2.860000 2.085000 ;
      RECT 1.115000  2.085000 1.285000 2.465000 ;
      RECT 1.195000  0.255000 1.415000 0.585000 ;
      RECT 1.245000  0.585000 1.415000 1.660000 ;
      RECT 1.705000  2.255000 2.425000 2.635000 ;
      RECT 2.670000  2.085000 2.860000 2.465000 ;
      RECT 2.690000  1.795000 3.465000 1.915000 ;
      RECT 3.010000  0.085000 3.390000 0.465000 ;
      RECT 3.140000  2.195000 3.470000 2.635000 ;
      RECT 3.295000  0.995000 3.555000 1.325000 ;
      RECT 3.295000  1.325000 3.465000 1.795000 ;
      RECT 4.065000  0.085000 4.450000 0.465000 ;
      RECT 4.195000  1.835000 4.450000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4b_2


MACRO sky130_fd_sc_hdll__xnor3_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.200000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.495000 1.075000 8.215000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.735900 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.625000 0.995000 6.845000 1.445000 ;
        RECT 6.625000 1.445000 7.255000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.715000 1.075000 2.330000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.472000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.345000 1.440000 ;
        RECT 0.085000 1.440000 0.365000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.515000  0.085000 0.815000 0.525000 ;
      RECT 0.515000  0.695000 1.205000 0.865000 ;
      RECT 0.515000  0.865000 0.755000 1.330000 ;
      RECT 0.535000  1.330000 0.755000 1.875000 ;
      RECT 0.535000  1.875000 1.320000 2.045000 ;
      RECT 0.535000  2.215000 0.920000 2.635000 ;
      RECT 0.985000  0.255000 2.655000 0.425000 ;
      RECT 0.985000  0.425000 1.205000 0.695000 ;
      RECT 0.985000  1.535000 2.670000 1.705000 ;
      RECT 1.100000  2.045000 1.320000 2.235000 ;
      RECT 1.100000  2.235000 2.670000 2.405000 ;
      RECT 1.375000  0.595000 1.545000 1.535000 ;
      RECT 1.660000  1.895000 4.360000 2.065000 ;
      RECT 1.845000  0.625000 3.165000 0.795000 ;
      RECT 1.845000  0.795000 2.225000 0.905000 ;
      RECT 2.170000  0.425000 2.655000 0.455000 ;
      RECT 2.500000  0.995000 2.825000 1.325000 ;
      RECT 2.500000  1.325000 2.670000 1.535000 ;
      RECT 2.875000  0.285000 3.505000 0.455000 ;
      RECT 2.890000  1.525000 3.275000 1.695000 ;
      RECT 2.995000  0.795000 3.165000 1.375000 ;
      RECT 2.995000  1.375000 3.275000 1.525000 ;
      RECT 3.335000  0.455000 3.505000 1.035000 ;
      RECT 3.335000  1.035000 3.615000 1.205000 ;
      RECT 3.425000  2.235000 3.755000 2.635000 ;
      RECT 3.445000  1.205000 3.615000 1.895000 ;
      RECT 3.675000  0.085000 3.845000 0.865000 ;
      RECT 3.845000  1.445000 4.365000 1.715000 ;
      RECT 4.075000  0.415000 4.365000 1.445000 ;
      RECT 4.190000  2.065000 4.360000 2.275000 ;
      RECT 4.190000  2.275000 7.485000 2.445000 ;
      RECT 4.545000  0.265000 4.955000 0.485000 ;
      RECT 4.545000  0.485000 4.755000 0.595000 ;
      RECT 4.545000  0.595000 4.715000 2.105000 ;
      RECT 4.885000  0.720000 5.345000 0.825000 ;
      RECT 4.885000  0.825000 5.145000 0.890000 ;
      RECT 4.885000  0.890000 5.055000 2.275000 ;
      RECT 4.925000  0.655000 5.345000 0.720000 ;
      RECT 5.175000  0.320000 5.345000 0.655000 ;
      RECT 5.285000  1.445000 6.115000 1.615000 ;
      RECT 5.285000  1.615000 5.700000 2.045000 ;
      RECT 5.300000  0.995000 5.725000 1.270000 ;
      RECT 5.515000  0.630000 5.725000 0.995000 ;
      RECT 5.945000  0.255000 7.140000 0.425000 ;
      RECT 5.945000  0.425000 6.115000 1.445000 ;
      RECT 6.285000  0.595000 6.455000 1.935000 ;
      RECT 6.285000  1.935000 9.110000 2.105000 ;
      RECT 6.625000  0.425000 7.140000 0.465000 ;
      RECT 7.015000  0.730000 7.220000 0.945000 ;
      RECT 7.015000  0.945000 7.325000 1.275000 ;
      RECT 7.475000  1.495000 8.660000 1.705000 ;
      RECT 7.515000  0.295000 7.805000 0.735000 ;
      RECT 7.515000  0.735000 8.660000 0.750000 ;
      RECT 7.555000  0.750000 8.660000 0.905000 ;
      RECT 7.915000  2.275000 8.595000 2.635000 ;
      RECT 8.050000  0.085000 8.510000 0.565000 ;
      RECT 8.490000  0.905000 8.660000 0.995000 ;
      RECT 8.490000  0.995000 8.770000 1.325000 ;
      RECT 8.490000  1.325000 8.660000 1.495000 ;
      RECT 8.575000  1.875000 9.110000 1.935000 ;
      RECT 8.810000  0.255000 9.110000 0.585000 ;
      RECT 8.815000  2.105000 9.110000 2.465000 ;
      RECT 8.940000  0.585000 9.110000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.105000  1.445000 3.275000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.075000  0.765000 4.245000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.585000  0.425000 4.755000 0.595000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.555000  0.765000 5.725000 0.935000 ;
      RECT 5.555000  1.445000 5.725000 1.615000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.035000  0.765000 7.205000 0.935000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.545000  0.425000 7.715000 0.595000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 3.045000 1.415000 3.335000 1.460000 ;
      RECT 3.045000 1.460000 5.785000 1.600000 ;
      RECT 3.045000 1.600000 3.335000 1.645000 ;
      RECT 4.015000 0.735000 4.305000 0.780000 ;
      RECT 4.015000 0.780000 7.265000 0.920000 ;
      RECT 4.015000 0.920000 4.305000 0.965000 ;
      RECT 4.525000 0.395000 4.815000 0.440000 ;
      RECT 4.525000 0.440000 7.775000 0.580000 ;
      RECT 4.525000 0.580000 4.815000 0.625000 ;
      RECT 5.495000 0.735000 5.785000 0.780000 ;
      RECT 5.495000 0.920000 5.785000 0.965000 ;
      RECT 5.495000 1.415000 5.785000 1.460000 ;
      RECT 5.495000 1.600000 5.785000 1.645000 ;
      RECT 6.975000 0.735000 7.265000 0.780000 ;
      RECT 6.975000 0.920000 7.265000 0.965000 ;
      RECT 7.485000 0.395000 7.775000 0.440000 ;
      RECT 7.485000 0.580000 7.775000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor3_1


MACRO sky130_fd_sc_hdll__xnor3_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.660000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.055000 1.075000 8.695000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.735900 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.135000 0.995000 7.355000 1.445000 ;
        RECT 7.135000 1.445000 7.765000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225000 1.075000 2.840000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.550500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.350000 0.865000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.735000 ;
      RECT 0.085000  1.490000 0.375000 2.635000 ;
      RECT 1.035000  0.085000 1.325000 0.525000 ;
      RECT 1.045000  0.695000 1.715000 0.865000 ;
      RECT 1.045000  0.865000 1.265000 1.875000 ;
      RECT 1.045000  1.875000 1.830000 2.045000 ;
      RECT 1.045000  2.215000 1.430000 2.635000 ;
      RECT 1.495000  0.255000 3.165000 0.425000 ;
      RECT 1.495000  0.425000 1.715000 0.695000 ;
      RECT 1.495000  1.535000 3.180000 1.705000 ;
      RECT 1.610000  2.045000 1.830000 2.235000 ;
      RECT 1.610000  2.235000 3.180000 2.405000 ;
      RECT 1.885000  0.595000 2.055000 1.535000 ;
      RECT 2.170000  1.895000 4.870000 2.065000 ;
      RECT 2.355000  0.625000 3.675000 0.795000 ;
      RECT 2.355000  0.795000 2.735000 0.905000 ;
      RECT 2.680000  0.425000 3.165000 0.455000 ;
      RECT 3.010000  0.995000 3.335000 1.325000 ;
      RECT 3.010000  1.325000 3.180000 1.535000 ;
      RECT 3.385000  0.285000 4.015000 0.455000 ;
      RECT 3.400000  1.525000 3.785000 1.695000 ;
      RECT 3.505000  0.795000 3.675000 1.375000 ;
      RECT 3.505000  1.375000 3.785000 1.525000 ;
      RECT 3.845000  0.455000 4.015000 1.035000 ;
      RECT 3.845000  1.035000 4.125000 1.205000 ;
      RECT 3.935000  2.235000 4.265000 2.635000 ;
      RECT 3.955000  1.205000 4.125000 1.895000 ;
      RECT 4.185000  0.085000 4.355000 0.865000 ;
      RECT 4.355000  1.445000 4.875000 1.715000 ;
      RECT 4.585000  0.415000 4.875000 1.445000 ;
      RECT 4.700000  2.065000 4.870000 2.275000 ;
      RECT 4.700000  2.275000 7.995000 2.445000 ;
      RECT 5.055000  0.265000 5.465000 0.485000 ;
      RECT 5.055000  0.485000 5.265000 0.595000 ;
      RECT 5.055000  0.595000 5.225000 2.105000 ;
      RECT 5.395000  0.720000 5.855000 0.825000 ;
      RECT 5.395000  0.825000 5.655000 0.890000 ;
      RECT 5.395000  0.890000 5.565000 2.275000 ;
      RECT 5.435000  0.655000 5.855000 0.720000 ;
      RECT 5.685000  0.320000 5.855000 0.655000 ;
      RECT 5.795000  1.445000 6.625000 1.615000 ;
      RECT 5.795000  1.615000 6.210000 2.045000 ;
      RECT 5.810000  0.995000 6.235000 1.270000 ;
      RECT 6.025000  0.630000 6.235000 0.995000 ;
      RECT 6.455000  0.255000 7.650000 0.425000 ;
      RECT 6.455000  0.425000 6.625000 1.445000 ;
      RECT 6.795000  0.595000 6.965000 1.935000 ;
      RECT 6.795000  1.935000 9.485000 2.105000 ;
      RECT 7.135000  0.425000 7.650000 0.465000 ;
      RECT 7.525000  0.730000 7.730000 0.945000 ;
      RECT 7.525000  0.945000 7.835000 1.275000 ;
      RECT 7.985000  1.495000 9.035000 1.705000 ;
      RECT 8.025000  0.295000 8.315000 0.735000 ;
      RECT 8.025000  0.735000 9.035000 0.750000 ;
      RECT 8.065000  0.750000 9.035000 0.905000 ;
      RECT 8.455000  2.275000 8.790000 2.635000 ;
      RECT 8.535000  0.085000 8.705000 0.565000 ;
      RECT 8.865000  0.905000 9.035000 0.995000 ;
      RECT 8.865000  0.995000 9.145000 1.325000 ;
      RECT 8.865000  1.325000 9.035000 1.495000 ;
      RECT 8.950000  1.875000 9.485000 1.935000 ;
      RECT 9.185000  0.255000 9.485000 0.585000 ;
      RECT 9.190000  2.105000 9.485000 2.465000 ;
      RECT 9.315000  0.585000 9.485000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.615000  1.445000 3.785000 1.615000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.585000  0.765000 4.755000 0.935000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.095000  0.425000 5.265000 0.595000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.065000  0.765000 6.235000 0.935000 ;
      RECT 6.065000  1.445000 6.235000 1.615000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.545000  0.765000 7.715000 0.935000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.055000  0.425000 8.225000 0.595000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 3.555000 1.415000 3.845000 1.460000 ;
      RECT 3.555000 1.460000 6.295000 1.600000 ;
      RECT 3.555000 1.600000 3.845000 1.645000 ;
      RECT 4.525000 0.735000 4.815000 0.780000 ;
      RECT 4.525000 0.780000 7.775000 0.920000 ;
      RECT 4.525000 0.920000 4.815000 0.965000 ;
      RECT 5.035000 0.395000 5.325000 0.440000 ;
      RECT 5.035000 0.440000 8.285000 0.580000 ;
      RECT 5.035000 0.580000 5.325000 0.625000 ;
      RECT 6.005000 0.735000 6.295000 0.780000 ;
      RECT 6.005000 0.920000 6.295000 0.965000 ;
      RECT 6.005000 1.415000 6.295000 1.460000 ;
      RECT 6.005000 1.600000 6.295000 1.645000 ;
      RECT 7.485000 0.735000 7.775000 0.780000 ;
      RECT 7.485000 0.920000 7.775000 0.965000 ;
      RECT 7.995000 0.395000 8.285000 0.440000 ;
      RECT 7.995000 0.580000 8.285000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor3_2


MACRO sky130_fd_sc_hdll__xnor3_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.58000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.075000 1.075000 9.535000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.735900 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.155000 0.995000 8.375000 1.445000 ;
        RECT 8.155000 1.445000 8.785000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.245000 1.075000 3.860000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.375000 0.925000 0.995000 ;
        RECT 0.625000 0.995000 1.860000 1.325000 ;
        RECT 0.625000 1.325000 1.005000 2.425000 ;
        RECT 1.565000 0.350000 1.875000 0.925000 ;
        RECT 1.565000 0.925000 1.860000 0.995000 ;
        RECT 1.565000 1.325000 1.860000 1.440000 ;
        RECT 1.565000 1.440000 1.895000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.285000  0.085000  0.455000 0.735000 ;
      RECT  0.285000  1.490000  0.455000 2.635000 ;
      RECT  1.225000  0.085000  1.395000 0.735000 ;
      RECT  1.225000  1.495000  1.395000 2.635000 ;
      RECT  2.030000  0.995000  2.285000 1.325000 ;
      RECT  2.045000  0.085000  2.345000 0.525000 ;
      RECT  2.060000  0.695000  2.735000 0.865000 ;
      RECT  2.060000  0.865000  2.285000 0.995000 ;
      RECT  2.065000  1.325000  2.285000 1.875000 ;
      RECT  2.065000  1.875000  2.850000 2.045000 ;
      RECT  2.065000  2.215000  2.450000 2.635000 ;
      RECT  2.515000  0.255000  4.185000 0.425000 ;
      RECT  2.515000  0.425000  2.735000 0.695000 ;
      RECT  2.515000  1.535000  4.200000 1.705000 ;
      RECT  2.630000  2.045000  2.850000 2.235000 ;
      RECT  2.630000  2.235000  4.200000 2.405000 ;
      RECT  2.905000  0.595000  3.075000 1.535000 ;
      RECT  3.190000  1.895000  5.890000 2.065000 ;
      RECT  3.375000  0.625000  4.695000 0.795000 ;
      RECT  3.375000  0.795000  3.755000 0.905000 ;
      RECT  3.700000  0.425000  4.185000 0.455000 ;
      RECT  4.030000  0.995000  4.355000 1.325000 ;
      RECT  4.030000  1.325000  4.200000 1.535000 ;
      RECT  4.405000  0.285000  5.035000 0.455000 ;
      RECT  4.420000  1.525000  4.805000 1.695000 ;
      RECT  4.525000  0.795000  4.695000 1.375000 ;
      RECT  4.525000  1.375000  4.805000 1.525000 ;
      RECT  4.865000  0.455000  5.035000 1.035000 ;
      RECT  4.865000  1.035000  5.145000 1.205000 ;
      RECT  4.955000  2.235000  5.285000 2.635000 ;
      RECT  4.975000  1.205000  5.145000 1.895000 ;
      RECT  5.205000  0.085000  5.375000 0.865000 ;
      RECT  5.375000  1.445000  5.895000 1.715000 ;
      RECT  5.605000  0.415000  5.895000 1.445000 ;
      RECT  5.720000  2.065000  5.890000 2.275000 ;
      RECT  5.720000  2.275000  9.015000 2.445000 ;
      RECT  6.075000  0.265000  6.520000 0.485000 ;
      RECT  6.075000  0.485000  6.245000 2.105000 ;
      RECT  6.415000  0.655000  6.875000 0.825000 ;
      RECT  6.415000  0.825000  6.585000 2.275000 ;
      RECT  6.705000  0.320000  6.875000 0.655000 ;
      RECT  6.815000  1.445000  7.645000 1.615000 ;
      RECT  6.815000  1.615000  7.230000 2.045000 ;
      RECT  6.830000  0.995000  7.255000 1.270000 ;
      RECT  7.045000  0.630000  7.255000 0.995000 ;
      RECT  7.475000  0.255000  8.670000 0.425000 ;
      RECT  7.475000  0.425000  7.645000 1.445000 ;
      RECT  7.815000  0.595000  7.985000 1.935000 ;
      RECT  7.815000  1.935000 10.325000 2.105000 ;
      RECT  8.155000  0.425000  8.670000 0.465000 ;
      RECT  8.545000  0.730000  8.750000 0.945000 ;
      RECT  8.545000  0.945000  8.855000 1.275000 ;
      RECT  9.005000  1.495000  9.875000 1.705000 ;
      RECT  9.045000  0.295000  9.335000 0.735000 ;
      RECT  9.045000  0.735000  9.875000 0.750000 ;
      RECT  9.085000  0.750000  9.875000 0.905000 ;
      RECT  9.425000  2.275000  9.810000 2.635000 ;
      RECT  9.555000  0.085000  9.725000 0.565000 ;
      RECT  9.705000  0.905000  9.875000 0.995000 ;
      RECT  9.705000  0.995000  9.985000 1.325000 ;
      RECT  9.705000  1.325000  9.875000 1.495000 ;
      RECT  9.790000  1.875000 10.325000 1.935000 ;
      RECT 10.025000  0.255000 10.325000 0.585000 ;
      RECT 10.030000  2.105000 10.325000 2.465000 ;
      RECT 10.155000  0.585000 10.325000 1.875000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.635000  1.445000  4.805000 1.615000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.605000  0.765000  5.775000 0.935000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.075000  0.425000  6.245000 0.595000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.085000  0.765000  7.255000 0.935000 ;
      RECT  7.085000  1.445000  7.255000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.565000  0.765000  8.735000 0.935000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.075000  0.425000  9.245000 0.595000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 4.575000 1.415000 4.865000 1.460000 ;
      RECT 4.575000 1.460000 7.315000 1.600000 ;
      RECT 4.575000 1.600000 4.865000 1.645000 ;
      RECT 5.545000 0.735000 5.835000 0.780000 ;
      RECT 5.545000 0.780000 8.795000 0.920000 ;
      RECT 5.545000 0.920000 5.835000 0.965000 ;
      RECT 6.015000 0.395000 6.315000 0.440000 ;
      RECT 6.015000 0.440000 9.305000 0.580000 ;
      RECT 6.015000 0.580000 6.315000 0.625000 ;
      RECT 7.025000 0.735000 7.315000 0.780000 ;
      RECT 7.025000 0.920000 7.315000 0.965000 ;
      RECT 7.025000 1.415000 7.315000 1.460000 ;
      RECT 7.025000 1.600000 7.315000 1.645000 ;
      RECT 8.505000 0.735000 8.795000 0.780000 ;
      RECT 8.505000 0.920000 8.795000 0.965000 ;
      RECT 9.015000 0.395000 9.305000 0.440000 ;
      RECT 9.015000 0.580000 9.305000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor3_4


MACRO sky130_fd_sc_hdll__or2_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.900000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.415000 1.075000 1.085000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.075000 2.025000 1.275000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.862000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 0.255000 3.285000 0.725000 ;
        RECT 2.985000 0.725000 6.335000 0.905000 ;
        RECT 2.985000 1.495000 6.335000 1.665000 ;
        RECT 2.985000 1.665000 3.315000 2.465000 ;
        RECT 3.925000 1.665000 4.255000 2.465000 ;
        RECT 3.955000 0.255000 4.225000 0.725000 ;
        RECT 4.865000 1.665000 5.195000 2.465000 ;
        RECT 4.895000 0.255000 5.165000 0.725000 ;
        RECT 5.805000 1.665000 6.135000 2.465000 ;
        RECT 5.835000 0.255000 6.105000 0.725000 ;
        RECT 5.935000 0.905000 6.335000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.090000  1.455000 1.355000 1.665000 ;
      RECT 0.090000  1.665000 0.415000 2.465000 ;
      RECT 0.145000  0.085000 0.415000 0.905000 ;
      RECT 0.585000  0.255000 0.915000 0.725000 ;
      RECT 0.585000  0.725000 1.855000 0.735000 ;
      RECT 0.585000  0.735000 2.375000 0.905000 ;
      RECT 0.585000  1.835000 0.915000 2.635000 ;
      RECT 1.085000  0.085000 1.355000 0.555000 ;
      RECT 1.085000  1.665000 1.355000 2.295000 ;
      RECT 1.085000  2.295000 2.325000 2.465000 ;
      RECT 1.525000  0.255000 1.855000 0.725000 ;
      RECT 1.525000  1.445000 2.375000 1.665000 ;
      RECT 1.525000  1.665000 1.855000 2.125000 ;
      RECT 2.025000  0.085000 2.815000 0.555000 ;
      RECT 2.025000  1.835000 2.325000 2.295000 ;
      RECT 2.195000  0.905000 2.375000 1.075000 ;
      RECT 2.195000  1.075000 5.525000 1.275000 ;
      RECT 2.195000  1.275000 2.375000 1.445000 ;
      RECT 2.545000  0.555000 2.815000 0.905000 ;
      RECT 2.545000  1.495000 2.815000 2.635000 ;
      RECT 3.455000  0.085000 3.785000 0.555000 ;
      RECT 3.485000  1.835000 3.755000 2.635000 ;
      RECT 4.395000  0.085000 4.725000 0.555000 ;
      RECT 4.425000  1.835000 4.695000 2.635000 ;
      RECT 5.335000  0.085000 5.665000 0.555000 ;
      RECT 5.365000  1.835000 5.635000 2.635000 ;
      RECT 6.275000  0.085000 6.605000 0.555000 ;
      RECT 6.305000  1.835000 6.575000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2_8


MACRO sky130_fd_sc_hdll__or2_6
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.415000 1.075000 1.085000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.075000 2.025000 1.275000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.396500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 0.255000 3.285000 0.725000 ;
        RECT 2.985000 0.725000 5.415000 0.905000 ;
        RECT 2.985000 1.495000 5.415000 1.665000 ;
        RECT 2.985000 1.665000 3.315000 2.465000 ;
        RECT 3.925000 1.665000 4.255000 2.465000 ;
        RECT 3.955000 0.255000 4.225000 0.725000 ;
        RECT 4.865000 1.665000 5.195000 2.465000 ;
        RECT 4.895000 0.255000 5.165000 0.725000 ;
        RECT 5.015000 0.905000 5.415000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.090000  1.455000 1.355000 1.665000 ;
      RECT 0.090000  1.665000 0.415000 2.465000 ;
      RECT 0.145000  0.085000 0.415000 0.905000 ;
      RECT 0.585000  0.255000 0.915000 0.725000 ;
      RECT 0.585000  0.725000 1.855000 0.735000 ;
      RECT 0.585000  0.735000 2.375000 0.905000 ;
      RECT 0.585000  1.835000 0.915000 2.635000 ;
      RECT 1.085000  0.085000 1.355000 0.555000 ;
      RECT 1.085000  1.665000 1.355000 2.295000 ;
      RECT 1.085000  2.295000 2.325000 2.465000 ;
      RECT 1.525000  0.255000 1.855000 0.725000 ;
      RECT 1.525000  1.445000 2.375000 1.665000 ;
      RECT 1.525000  1.665000 1.855000 2.125000 ;
      RECT 2.025000  0.085000 2.815000 0.555000 ;
      RECT 2.025000  1.835000 2.325000 2.295000 ;
      RECT 2.195000  0.905000 2.375000 1.075000 ;
      RECT 2.195000  1.075000 4.845000 1.275000 ;
      RECT 2.195000  1.275000 2.375000 1.445000 ;
      RECT 2.545000  0.555000 2.815000 0.905000 ;
      RECT 2.545000  1.495000 2.815000 2.635000 ;
      RECT 3.455000  0.085000 3.785000 0.555000 ;
      RECT 3.485000  1.835000 3.755000 2.635000 ;
      RECT 4.395000  0.085000 4.725000 0.555000 ;
      RECT 4.425000  1.835000 4.695000 2.635000 ;
      RECT 5.335000  0.085000 5.665000 0.555000 ;
      RECT 5.365000  1.835000 5.635000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2_6


MACRO sky130_fd_sc_hdll__or2_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.915000 0.765000 1.375000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.765000 0.345000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.540000 1.835000 2.415000 2.005000 ;
        RECT 1.540000 2.005000 1.920000 2.465000 ;
        RECT 1.670000 0.385000 1.840000 0.655000 ;
        RECT 1.670000 0.655000 2.415000 0.825000 ;
        RECT 1.935000 0.825000 2.415000 1.835000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.105000  0.085000 0.345000 0.595000 ;
      RECT 0.155000  1.495000 1.765000 1.665000 ;
      RECT 0.155000  1.665000 0.515000 1.840000 ;
      RECT 0.515000  0.255000 0.855000 0.595000 ;
      RECT 0.515000  0.595000 0.745000 1.495000 ;
      RECT 1.135000  0.085000 1.450000 0.595000 ;
      RECT 1.200000  1.835000 1.370000 2.635000 ;
      RECT 1.545000  0.995000 1.765000 1.495000 ;
      RECT 2.010000  0.085000 2.390000 0.485000 ;
      RECT 2.140000  2.175000 2.310000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2_2


MACRO sky130_fd_sc_hdll__or2_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.765000 1.285000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.440000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.551500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 0.255000 2.215000 0.825000 ;
        RECT 1.645000 1.845000 2.215000 2.465000 ;
        RECT 1.915000 0.825000 2.215000 1.845000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.110000  0.085000 0.350000 0.595000 ;
      RECT 0.120000  1.495000 1.745000 1.665000 ;
      RECT 0.120000  1.665000 0.510000 1.840000 ;
      RECT 0.610000  0.265000 0.850000 0.595000 ;
      RECT 0.610000  0.595000 0.780000 1.495000 ;
      RECT 1.095000  1.835000 1.425000 2.635000 ;
      RECT 1.130000  0.085000 1.345000 0.595000 ;
      RECT 1.525000  0.995000 1.745000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2_1


MACRO sky130_fd_sc_hdll__or2_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.915000 0.995000 1.340000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.765000 0.345000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.590000 0.265000 1.970000 0.735000 ;
        RECT 1.590000 0.735000 3.170000 0.905000 ;
        RECT 1.590000 1.835000 2.910000 2.005000 ;
        RECT 1.590000 2.005000 1.970000 2.465000 ;
        RECT 2.530000 0.265000 2.910000 0.735000 ;
        RECT 2.530000 1.495000 3.170000 1.665000 ;
        RECT 2.530000 1.665000 2.910000 1.835000 ;
        RECT 2.530000 2.005000 2.910000 2.465000 ;
        RECT 2.825000 0.905000 3.170000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.105000  0.085000 0.345000 0.595000 ;
      RECT 0.155000  1.495000 1.765000 1.665000 ;
      RECT 0.155000  1.665000 0.515000 2.465000 ;
      RECT 0.515000  0.290000 0.895000 0.825000 ;
      RECT 0.515000  0.825000 0.745000 1.495000 ;
      RECT 1.160000  0.085000 1.330000 0.825000 ;
      RECT 1.160000  1.835000 1.330000 2.635000 ;
      RECT 1.510000  1.075000 2.620000 1.245000 ;
      RECT 1.510000  1.245000 1.765000 1.495000 ;
      RECT 2.140000  0.085000 2.310000 0.565000 ;
      RECT 2.140000  2.175000 2.310000 2.635000 ;
      RECT 3.080000  0.085000 3.250000 0.565000 ;
      RECT 3.080000  1.835000 3.250000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2_4


MACRO sky130_fd_sc_hdll__sdfsbp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  14.72000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855000 1.720000 3.335000 1.970000 ;
        RECT 3.155000 1.055000 3.815000 1.590000 ;
        RECT 3.155000 1.590000 3.335000 1.720000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 0.765000 1.425000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.065000 0.275000 14.625000 0.825000 ;
        RECT 14.065000 1.495000 14.625000 2.450000 ;
        RECT 14.270000 0.825000 14.625000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.471500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.550000 0.255000 12.930000 2.465000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.365000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.467400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.570000 1.075000 0.860000 1.120000 ;
        RECT 0.570000 1.120000 2.875000 1.260000 ;
        RECT 0.570000 1.260000 0.860000 1.305000 ;
        RECT 2.585000 1.075000 2.875000 1.120000 ;
        RECT 2.585000 1.260000 2.875000 1.305000 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.385000 1.415000 7.725000 1.460000 ;
        RECT 7.385000 1.460000 9.965000 1.600000 ;
        RECT 7.385000 1.600000 7.725000 1.645000 ;
        RECT 9.675000 1.415000 9.965000 1.460000 ;
        RECT 9.675000 1.600000 9.965000 1.645000 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.720000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.720000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.720000 0.085000 ;
      RECT  0.000000  2.635000 14.720000 2.805000 ;
      RECT  0.085000  0.085000  0.430000 0.595000 ;
      RECT  0.085000  1.845000  1.205000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.815000 2.635000 ;
      RECT  0.550000  0.765000  0.860000 1.675000 ;
      RECT  0.975000  0.280000  1.845000 0.560000 ;
      RECT  1.035000  2.025000  1.205000 2.255000 ;
      RECT  1.035000  2.255000  2.245000 2.465000 ;
      RECT  1.395000  1.870000  1.845000 2.075000 ;
      RECT  1.655000  0.560000  1.845000 1.870000 ;
      RECT  2.025000  0.085000  2.205000 0.545000 ;
      RECT  2.065000  0.715000  2.715000 0.905000 ;
      RECT  2.065000  0.905000  2.400000 1.770000 ;
      RECT  2.065000  1.770000  2.685000 2.085000 ;
      RECT  2.460000  0.255000  2.715000 0.715000 ;
      RECT  2.470000  2.085000  2.685000 2.465000 ;
      RECT  2.570000  1.075000  2.950000 1.550000 ;
      RECT  2.940000  0.085000  3.280000 0.555000 ;
      RECT  2.940000  2.140000  3.280000 2.635000 ;
      RECT  3.505000  1.775000  4.295000 1.955000 ;
      RECT  3.505000  1.955000  3.675000 2.325000 ;
      RECT  3.520000  0.255000  3.705000 0.715000 ;
      RECT  3.520000  0.715000  4.295000 0.885000 ;
      RECT  3.845000  2.275000  4.225000 2.635000 ;
      RECT  3.930000  0.085000  4.240000 0.545000 ;
      RECT  4.035000  0.885000  4.295000 1.775000 ;
      RECT  4.445000  2.135000  4.790000 2.465000 ;
      RECT  4.460000  0.255000  4.685000 0.585000 ;
      RECT  4.515000  0.585000  4.685000 1.090000 ;
      RECT  4.515000  1.090000  4.840000 1.420000 ;
      RECT  4.515000  1.420000  4.790000 2.135000 ;
      RECT  4.855000  0.255000  5.180000 0.920000 ;
      RECT  4.960000  1.590000  5.180000 2.465000 ;
      RECT  5.010000  0.920000  5.180000 1.590000 ;
      RECT  5.400000  0.255000  5.890000 1.225000 ;
      RECT  5.400000  1.225000  8.360000 1.275000 ;
      RECT  5.430000  2.135000  6.205000 2.465000 ;
      RECT  5.485000  1.275000  6.935000 1.395000 ;
      RECT  5.605000  1.575000  5.865000 1.955000 ;
      RECT  6.035000  1.395000  6.205000 2.135000 ;
      RECT  6.060000  0.085000  6.595000 0.465000 ;
      RECT  6.060000  0.635000  7.085000 0.805000 ;
      RECT  6.060000  0.805000  6.475000 1.015000 ;
      RECT  6.425000  1.575000  6.595000 1.935000 ;
      RECT  6.425000  1.935000  7.365000 2.105000 ;
      RECT  6.445000  2.275000  6.775000 2.635000 ;
      RECT  6.750000  0.975000  8.360000 1.225000 ;
      RECT  6.775000  0.255000  7.085000 0.635000 ;
      RECT  7.100000  2.105000  7.365000 2.450000 ;
      RECT  7.190000  1.445000  7.725000 1.765000 ;
      RECT  7.540000  0.085000  8.275000 0.690000 ;
      RECT  7.655000  2.125000  8.710000 2.635000 ;
      RECT  7.910000  1.495000  8.755000 1.955000 ;
      RECT  7.950000  1.275000  8.360000 1.325000 ;
      RECT  8.535000  0.695000  9.890000 0.895000 ;
      RECT  8.535000  0.895000  8.755000 1.495000 ;
      RECT  8.880000  2.125000  9.735000 2.460000 ;
      RECT  9.115000  1.075000  9.395000 1.905000 ;
      RECT  9.160000  0.275000 10.775000 0.445000 ;
      RECT  9.565000  1.895000 11.465000 2.065000 ;
      RECT  9.565000  2.065000  9.735000 2.125000 ;
      RECT  9.610000  0.895000  9.890000 1.245000 ;
      RECT  9.685000  1.415000  9.960000 1.525000 ;
      RECT  9.685000  1.525000 11.075000 1.725000 ;
      RECT 10.045000  2.235000 10.425000 2.635000 ;
      RECT 10.140000  0.855000 10.365000 1.185000 ;
      RECT 10.140000  1.185000 11.945000 1.355000 ;
      RECT 10.605000  0.445000 10.775000 0.845000 ;
      RECT 10.605000  0.845000 11.545000 1.015000 ;
      RECT 10.645000  2.065000 10.860000 2.450000 ;
      RECT 11.135000  2.235000 11.465000 2.635000 ;
      RECT 11.220000  0.085000 11.390000 0.545000 ;
      RECT 11.245000  1.525000 11.465000 1.895000 ;
      RECT 11.560000  0.255000 11.945000 0.540000 ;
      RECT 11.685000  1.355000 11.945000 2.465000 ;
      RECT 11.765000  0.540000 11.945000 1.185000 ;
      RECT 12.170000  0.085000 12.380000 0.885000 ;
      RECT 12.170000  1.485000 12.380000 2.635000 ;
      RECT 13.160000  0.255000 13.370000 0.995000 ;
      RECT 13.160000  0.995000 14.050000 1.325000 ;
      RECT 13.160000  1.325000 13.370000 2.465000 ;
      RECT 13.690000  0.085000 13.895000 0.825000 ;
      RECT 13.725000  1.575000 13.895000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.630000  1.105000  0.800000 1.275000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.675000  1.445000  1.845000 1.615000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.645000  1.105000  2.815000 1.275000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.125000  1.785000  4.295000 1.955000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.585000  1.105000  4.755000 1.275000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.010000  1.445000  5.180000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.605000  1.785000  5.775000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.445000  1.445000  7.615000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.205000  1.785000  8.375000 1.955000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.225000  1.105000  9.395000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.735000  1.445000  9.905000 1.615000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
    LAYER met1 ;
      RECT 1.615000 1.415000 1.955000 1.460000 ;
      RECT 1.615000 1.460000 5.240000 1.600000 ;
      RECT 1.615000 1.600000 1.955000 1.645000 ;
      RECT 4.065000 1.755000 4.405000 1.800000 ;
      RECT 4.065000 1.800000 8.435000 1.940000 ;
      RECT 4.065000 1.940000 4.405000 1.985000 ;
      RECT 4.525000 1.075000 4.815000 1.120000 ;
      RECT 4.525000 1.120000 9.455000 1.260000 ;
      RECT 4.525000 1.260000 4.815000 1.305000 ;
      RECT 4.950000 1.415000 5.240000 1.460000 ;
      RECT 4.950000 1.600000 5.240000 1.645000 ;
      RECT 5.545000 1.755000 5.885000 1.800000 ;
      RECT 5.545000 1.940000 5.885000 1.985000 ;
      RECT 8.145000 1.755000 8.435000 1.800000 ;
      RECT 8.145000 1.940000 8.435000 1.985000 ;
      RECT 9.115000 1.075000 9.455000 1.120000 ;
      RECT 9.115000 1.260000 9.455000 1.305000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfsbp_1


MACRO sky130_fd_sc_hdll__sdfsbp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  15.64000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855000 1.720000 3.335000 1.970000 ;
        RECT 3.155000 1.055000 3.815000 1.590000 ;
        RECT 3.155000 1.590000 3.335000 1.720000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 0.765000 1.425000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.700000 0.275000 15.080000 0.825000 ;
        RECT 14.700000 1.495000 15.080000 2.450000 ;
        RECT 14.805000 0.825000 15.080000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.555000 0.255000 13.000000 2.465000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.365000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.467400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.570000 1.075000 0.860000 1.120000 ;
        RECT 0.570000 1.120000 2.875000 1.260000 ;
        RECT 0.570000 1.260000 0.860000 1.305000 ;
        RECT 2.585000 1.075000 2.875000 1.120000 ;
        RECT 2.585000 1.260000 2.875000 1.305000 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.385000 1.415000 7.725000 1.460000 ;
        RECT 7.385000 1.460000 9.965000 1.600000 ;
        RECT 7.385000 1.600000 7.725000 1.645000 ;
        RECT 9.675000 1.415000 9.965000 1.460000 ;
        RECT 9.675000 1.600000 9.965000 1.645000 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.640000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 15.640000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.640000 0.085000 ;
      RECT  0.000000  2.635000 15.640000 2.805000 ;
      RECT  0.085000  0.085000  0.430000 0.595000 ;
      RECT  0.085000  1.845000  1.205000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.815000 2.635000 ;
      RECT  0.550000  0.765000  0.860000 1.675000 ;
      RECT  0.975000  0.280000  1.845000 0.560000 ;
      RECT  1.035000  2.025000  1.205000 2.255000 ;
      RECT  1.035000  2.255000  2.245000 2.465000 ;
      RECT  1.395000  1.870000  1.845000 2.075000 ;
      RECT  1.655000  0.560000  1.845000 1.870000 ;
      RECT  2.025000  0.085000  2.205000 0.545000 ;
      RECT  2.065000  0.715000  2.715000 0.905000 ;
      RECT  2.065000  0.905000  2.400000 1.770000 ;
      RECT  2.065000  1.770000  2.685000 2.085000 ;
      RECT  2.460000  0.255000  2.715000 0.715000 ;
      RECT  2.470000  2.085000  2.685000 2.465000 ;
      RECT  2.570000  1.075000  2.950000 1.550000 ;
      RECT  2.940000  0.085000  3.280000 0.555000 ;
      RECT  2.940000  2.140000  3.280000 2.635000 ;
      RECT  3.505000  1.775000  4.295000 1.955000 ;
      RECT  3.505000  1.955000  3.675000 2.325000 ;
      RECT  3.520000  0.255000  3.705000 0.715000 ;
      RECT  3.520000  0.715000  4.295000 0.885000 ;
      RECT  3.845000  2.275000  4.225000 2.635000 ;
      RECT  3.930000  0.085000  4.240000 0.545000 ;
      RECT  4.035000  0.885000  4.295000 1.775000 ;
      RECT  4.445000  2.135000  4.790000 2.465000 ;
      RECT  4.460000  0.255000  4.685000 0.585000 ;
      RECT  4.515000  0.585000  4.685000 1.090000 ;
      RECT  4.515000  1.090000  4.840000 1.420000 ;
      RECT  4.515000  1.420000  4.790000 2.135000 ;
      RECT  4.855000  0.255000  5.180000 0.920000 ;
      RECT  4.960000  1.590000  5.180000 2.465000 ;
      RECT  5.010000  0.920000  5.180000 1.590000 ;
      RECT  5.400000  0.255000  5.890000 1.225000 ;
      RECT  5.400000  1.225000  8.360000 1.275000 ;
      RECT  5.430000  2.135000  6.205000 2.465000 ;
      RECT  5.485000  1.275000  6.935000 1.395000 ;
      RECT  5.605000  1.575000  5.865000 1.955000 ;
      RECT  6.035000  1.395000  6.205000 2.135000 ;
      RECT  6.060000  0.085000  6.595000 0.465000 ;
      RECT  6.060000  0.635000  7.085000 0.805000 ;
      RECT  6.060000  0.805000  6.475000 1.015000 ;
      RECT  6.425000  1.575000  6.595000 1.935000 ;
      RECT  6.425000  1.935000  7.365000 2.105000 ;
      RECT  6.445000  2.275000  6.775000 2.635000 ;
      RECT  6.750000  0.975000  8.360000 1.225000 ;
      RECT  6.775000  0.255000  7.085000 0.635000 ;
      RECT  7.100000  2.105000  7.365000 2.450000 ;
      RECT  7.190000  1.445000  7.725000 1.765000 ;
      RECT  7.540000  0.085000  8.275000 0.690000 ;
      RECT  7.655000  2.125000  8.710000 2.635000 ;
      RECT  7.910000  1.495000  8.755000 1.955000 ;
      RECT  7.950000  1.275000  8.360000 1.325000 ;
      RECT  8.535000  0.695000  9.890000 0.895000 ;
      RECT  8.535000  0.895000  8.755000 1.495000 ;
      RECT  8.880000  2.125000  9.735000 2.460000 ;
      RECT  9.115000  1.075000  9.395000 1.905000 ;
      RECT  9.160000  0.275000 10.775000 0.445000 ;
      RECT  9.565000  1.895000 11.465000 2.065000 ;
      RECT  9.565000  2.065000  9.735000 2.125000 ;
      RECT  9.610000  0.895000  9.890000 1.245000 ;
      RECT  9.685000  1.415000  9.960000 1.525000 ;
      RECT  9.685000  1.525000 11.075000 1.725000 ;
      RECT 10.045000  2.235000 10.425000 2.635000 ;
      RECT 10.140000  0.855000 10.365000 1.185000 ;
      RECT 10.140000  1.185000 11.945000 1.355000 ;
      RECT 10.605000  0.445000 10.775000 0.845000 ;
      RECT 10.605000  0.845000 11.545000 1.015000 ;
      RECT 10.645000  2.065000 10.860000 2.450000 ;
      RECT 11.135000  2.235000 11.465000 2.635000 ;
      RECT 11.220000  0.085000 11.390000 0.545000 ;
      RECT 11.245000  1.525000 11.465000 1.895000 ;
      RECT 11.560000  0.255000 11.945000 0.540000 ;
      RECT 11.685000  1.355000 11.945000 2.465000 ;
      RECT 11.765000  0.540000 11.945000 1.185000 ;
      RECT 12.170000  0.085000 12.380000 0.885000 ;
      RECT 12.170000  1.485000 12.380000 2.635000 ;
      RECT 13.215000  0.085000 13.505000 0.885000 ;
      RECT 13.215000  1.485000 13.505000 2.635000 ;
      RECT 13.720000  0.255000 13.905000 0.995000 ;
      RECT 13.720000  0.995000 14.585000 1.325000 ;
      RECT 13.720000  1.325000 13.905000 2.465000 ;
      RECT 14.075000  0.085000 14.480000 0.825000 ;
      RECT 14.075000  1.635000 14.480000 2.635000 ;
      RECT 15.250000  0.085000 15.515000 0.885000 ;
      RECT 15.250000  1.485000 15.515000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.630000  1.105000  0.800000 1.275000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.675000  1.445000  1.845000 1.615000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.645000  1.105000  2.815000 1.275000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.125000  1.785000  4.295000 1.955000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.585000  1.105000  4.755000 1.275000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.010000  1.445000  5.180000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.605000  1.785000  5.775000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.445000  1.445000  7.615000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.205000  1.785000  8.375000 1.955000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.225000  1.105000  9.395000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.735000  1.445000  9.905000 1.615000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
    LAYER met1 ;
      RECT 1.615000 1.415000 1.955000 1.460000 ;
      RECT 1.615000 1.460000 5.240000 1.600000 ;
      RECT 1.615000 1.600000 1.955000 1.645000 ;
      RECT 4.065000 1.755000 4.405000 1.800000 ;
      RECT 4.065000 1.800000 8.435000 1.940000 ;
      RECT 4.065000 1.940000 4.405000 1.985000 ;
      RECT 4.525000 1.075000 4.815000 1.120000 ;
      RECT 4.525000 1.120000 9.455000 1.260000 ;
      RECT 4.525000 1.260000 4.815000 1.305000 ;
      RECT 4.950000 1.415000 5.240000 1.460000 ;
      RECT 4.950000 1.600000 5.240000 1.645000 ;
      RECT 5.545000 1.755000 5.885000 1.800000 ;
      RECT 5.545000 1.940000 5.885000 1.985000 ;
      RECT 8.145000 1.755000 8.435000 1.800000 ;
      RECT 8.145000 1.940000 8.435000 1.985000 ;
      RECT 9.115000 1.075000 9.455000 1.120000 ;
      RECT 9.115000 1.260000 9.455000 1.305000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfsbp_2


MACRO sky130_fd_sc_hdll__nand4bb_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.070000 0.940000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.070000 0.330000 1.615000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.240000 1.075000 4.950000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.315000 1.075000 6.295000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.368000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.185000 0.655000 2.630000 1.445000 ;
        RECT 2.185000 1.445000 5.875000 1.665000 ;
        RECT 2.185000 1.665000 2.485000 2.465000 ;
        RECT 3.125000 1.665000 3.505000 2.465000 ;
        RECT 3.495000 1.075000 4.045000 1.445000 ;
        RECT 4.555000 1.665000 4.935000 2.465000 ;
        RECT 5.495000 1.665000 5.875000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.730000 ;
      RECT 0.085000  0.730000 1.330000 0.900000 ;
      RECT 0.085000  1.785000 1.330000 1.980000 ;
      RECT 0.085000  1.980000 0.370000 2.440000 ;
      RECT 0.515000  0.085000 0.815000 0.545000 ;
      RECT 0.540000  2.195000 0.815000 2.635000 ;
      RECT 0.985000  0.255000 1.675000 0.560000 ;
      RECT 0.985000  2.150000 1.675000 2.465000 ;
      RECT 1.160000  0.900000 1.330000 1.785000 ;
      RECT 1.500000  0.560000 1.675000 2.150000 ;
      RECT 1.845000  0.255000 3.975000 0.485000 ;
      RECT 1.845000  0.485000 2.015000 0.585000 ;
      RECT 1.845000  1.495000 2.015000 2.635000 ;
      RECT 2.655000  1.835000 2.955000 2.635000 ;
      RECT 2.945000  1.075000 3.325000 1.275000 ;
      RECT 3.125000  0.655000 4.935000 0.905000 ;
      RECT 3.725000  1.835000 4.385000 2.635000 ;
      RECT 4.165000  0.255000 5.405000 0.485000 ;
      RECT 5.155000  0.485000 5.405000 0.735000 ;
      RECT 5.155000  0.735000 6.345000 0.905000 ;
      RECT 5.155000  1.835000 5.325000 2.635000 ;
      RECT 5.625000  0.085000 5.795000 0.565000 ;
      RECT 5.965000  0.255000 6.345000 0.735000 ;
      RECT 6.095000  1.445000 6.345000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.160000  1.105000 1.330000 1.275000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.155000  1.105000 3.325000 1.275000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 1.100000 1.075000 3.385000 1.305000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4bb_2


MACRO sky130_fd_sc_hdll__nand4bb_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.300000 0.725000 3.710000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.075000 0.825000 1.655000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 0.735000 1.760000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.075000 1.325000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.901500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.155000 1.495000 2.680000 1.665000 ;
        RECT 1.155000 1.665000 1.485000 2.465000 ;
        RECT 2.190000 1.665000 2.680000 2.005000 ;
        RECT 2.190000 2.005000 2.580000 2.465000 ;
        RECT 2.410000 0.255000 3.000000 0.825000 ;
        RECT 2.410000 0.825000 2.680000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.485000 0.425000 0.715000 ;
      RECT 0.085000  0.715000 1.220000 0.905000 ;
      RECT 0.085000  0.905000 0.260000 2.065000 ;
      RECT 0.085000  2.065000 0.425000 2.465000 ;
      RECT 0.645000  0.085000 0.880000 0.545000 ;
      RECT 0.645000  1.835000 0.975000 2.635000 ;
      RECT 1.050000  0.365000 2.240000 0.555000 ;
      RECT 1.050000  0.555000 1.220000 0.715000 ;
      RECT 1.695000  1.835000 2.015000 2.635000 ;
      RECT 1.990000  0.555000 2.240000 1.325000 ;
      RECT 2.750000  2.175000 3.520000 2.635000 ;
      RECT 2.850000  0.995000 3.125000 1.835000 ;
      RECT 2.850000  1.835000 4.055000 2.005000 ;
      RECT 3.190000  0.085000 3.540000 0.545000 ;
      RECT 3.710000  0.255000 4.055000 0.545000 ;
      RECT 3.740000  2.005000 4.055000 2.465000 ;
      RECT 3.885000  0.545000 4.055000 1.835000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4bb_1


MACRO sky130_fd_sc_hdll__nand4bb_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.58000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.995000 0.330000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 0.995000 1.025000 1.615000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.045000 1.075000 7.985000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.395000 1.075000 10.340000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.736000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.355000 0.655000 4.015000 0.905000 ;
        RECT 2.355000 1.445000 9.865000 1.665000 ;
        RECT 2.355000 1.665000 2.655000 2.465000 ;
        RECT 3.295000 1.665000 3.675000 2.465000 ;
        RECT 3.665000 0.905000 4.015000 1.445000 ;
        RECT 4.235000 1.665000 4.615000 2.465000 ;
        RECT 5.175000 1.665000 5.555000 2.465000 ;
        RECT 6.665000 1.665000 7.045000 2.465000 ;
        RECT 7.605000 1.665000 7.985000 2.465000 ;
        RECT 8.545000 1.665000 8.925000 2.465000 ;
        RECT 9.485000 1.665000 9.865000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.085000  0.255000  0.345000 0.635000 ;
      RECT  0.085000  0.635000  1.505000 0.805000 ;
      RECT  0.085000  1.785000  1.505000 1.980000 ;
      RECT  0.085000  1.980000  0.370000 2.440000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.540000  2.195000  0.815000 2.635000 ;
      RECT  0.985000  2.150000  1.845000 2.465000 ;
      RECT  1.115000  0.255000  1.845000 0.465000 ;
      RECT  1.195000  0.805000  1.505000 1.785000 ;
      RECT  1.675000  0.465000  1.845000 1.075000 ;
      RECT  1.675000  1.075000  2.025000 1.305000 ;
      RECT  1.675000  1.305000  1.845000 2.150000 ;
      RECT  2.015000  0.255000  6.025000 0.485000 ;
      RECT  2.015000  0.485000  2.185000 0.905000 ;
      RECT  2.015000  1.495000  2.185000 2.635000 ;
      RECT  2.355000  1.075000  3.200000 1.245000 ;
      RECT  2.825000  1.835000  3.125000 2.635000 ;
      RECT  3.895000  1.835000  4.065000 2.635000 ;
      RECT  4.185000  1.075000  5.555000 1.275000 ;
      RECT  4.235000  0.655000  8.010000 0.905000 ;
      RECT  4.835000  1.835000  5.005000 2.635000 ;
      RECT  5.825000  1.835000  6.465000 2.635000 ;
      RECT  6.265000  0.255000  8.375000 0.485000 ;
      RECT  7.265000  1.835000  7.435000 2.635000 ;
      RECT  8.205000  0.485000  8.375000 0.655000 ;
      RECT  8.205000  0.655000 10.285000 0.825000 ;
      RECT  8.205000  1.835000  8.375000 2.635000 ;
      RECT  8.595000  0.085000  8.925000 0.485000 ;
      RECT  9.145000  1.835000  9.315000 2.635000 ;
      RECT  9.535000  0.085000  9.865000 0.485000 ;
      RECT 10.085000  1.445000 10.360000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.795000  1.105000  1.965000 1.275000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.330000  1.105000  4.500000 1.275000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 1.735000 1.075000 2.025000 1.120000 ;
      RECT 1.735000 1.120000 4.575000 1.260000 ;
      RECT 1.735000 1.260000 2.025000 1.305000 ;
      RECT 4.235000 1.075000 4.575000 1.120000 ;
      RECT 4.235000 1.260000 4.575000 1.305000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4bb_4


MACRO sky130_fd_sc_hdll__muxb8to1_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  24.84000 BY  5.440000 ;
  SITE unithd ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.655000 1.055000 6.045000 1.325000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.655000 4.115000 6.045000 4.385000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.375000 1.055000 7.765000 1.325000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.375000 4.115000 7.765000 4.385000 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.075000 1.055000 18.465000 1.325000 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.075000 4.115000 18.465000 4.385000 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.795000 1.055000 20.185000 1.325000 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.795000 4.115000 20.185000 4.385000 ;
    END
  END D[7]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.680000 1.325000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 4.115000 0.680000 4.445000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.740000 0.995000 12.335000 1.325000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.740000 4.115000 12.335000 4.445000 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.505000 0.995000 13.100000 1.325000 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.505000 4.115000 13.100000 4.445000 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.160000 0.995000 24.755000 1.325000 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.160000 4.115000 24.755000 4.445000 ;
    END
  END S[7]
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  2.225000 1.755000  2.515000 1.800000 ;
        RECT  2.225000 1.800000 22.615000 1.940000 ;
        RECT  2.225000 1.940000  2.515000 1.985000 ;
        RECT  2.225000 3.455000  2.515000 3.500000 ;
        RECT  2.225000 3.500000 22.615000 3.640000 ;
        RECT  2.225000 3.640000  2.515000 3.685000 ;
        RECT  3.165000 1.755000  3.455000 1.800000 ;
        RECT  3.165000 1.940000  3.455000 1.985000 ;
        RECT  3.165000 3.455000  3.455000 3.500000 ;
        RECT  3.165000 3.640000  3.455000 3.685000 ;
        RECT  8.965000 1.755000  9.255000 1.800000 ;
        RECT  8.965000 1.940000  9.255000 1.985000 ;
        RECT  8.965000 3.455000  9.255000 3.500000 ;
        RECT  8.965000 3.640000  9.255000 3.685000 ;
        RECT  9.905000 1.755000 10.195000 1.800000 ;
        RECT  9.905000 1.940000 10.195000 1.985000 ;
        RECT  9.905000 3.455000 10.195000 3.500000 ;
        RECT  9.905000 3.640000 10.195000 3.685000 ;
        RECT 14.645000 1.755000 14.935000 1.800000 ;
        RECT 14.645000 1.940000 14.935000 1.985000 ;
        RECT 14.645000 3.455000 14.935000 3.500000 ;
        RECT 14.645000 3.640000 14.935000 3.685000 ;
        RECT 15.585000 1.755000 15.875000 1.800000 ;
        RECT 15.585000 1.940000 15.875000 1.985000 ;
        RECT 15.585000 3.455000 15.875000 3.500000 ;
        RECT 15.585000 3.640000 15.875000 3.685000 ;
        RECT 21.385000 1.755000 21.675000 1.800000 ;
        RECT 21.385000 1.940000 21.675000 1.985000 ;
        RECT 21.385000 3.455000 21.675000 3.500000 ;
        RECT 21.385000 3.640000 21.675000 3.685000 ;
        RECT 22.325000 1.755000 22.615000 1.800000 ;
        RECT 22.325000 1.940000 22.615000 1.985000 ;
        RECT 22.325000 3.455000 22.615000 3.500000 ;
        RECT 22.325000 3.640000 22.615000 3.685000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 24.840000 0.240000 ;
        RECT 0.000000  5.200000 24.840000 5.680000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 24.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 24.840000 0.085000 ;
      RECT  0.000000  2.635000  2.035000 2.805000 ;
      RECT  0.000000  5.355000 24.840000 5.525000 ;
      RECT  0.220000  1.605000  0.520000 2.635000 ;
      RECT  0.220000  2.805000  0.520000 3.835000 ;
      RECT  0.270000  0.085000  0.560000 0.610000 ;
      RECT  0.270000  4.830000  0.560000 5.355000 ;
      RECT  0.690000  1.605000  1.020000 2.465000 ;
      RECT  0.690000  2.975000  1.020000 3.835000 ;
      RECT  0.770000  0.280000  1.020000 0.825000 ;
      RECT  0.770000  4.615000  1.020000 5.160000 ;
      RECT  0.850000  0.825000  1.020000 1.065000 ;
      RECT  0.850000  1.065000  2.035000 1.395000 ;
      RECT  0.850000  1.395000  1.020000 1.605000 ;
      RECT  0.850000  3.835000  1.020000 4.045000 ;
      RECT  0.850000  4.045000  2.035000 4.375000 ;
      RECT  0.850000  4.375000  1.020000 4.615000 ;
      RECT  1.190000  0.085000  1.480000 0.610000 ;
      RECT  1.190000  4.830000  1.480000 5.355000 ;
      RECT  1.215000  1.605000  1.490000 2.635000 ;
      RECT  1.215000  2.805000  1.490000 3.835000 ;
      RECT  1.735000  1.565000  2.035000 2.465000 ;
      RECT  1.735000  2.975000  2.035000 3.875000 ;
      RECT  1.985000  0.255000  4.015000 0.425000 ;
      RECT  1.985000  0.425000  2.235000 0.770000 ;
      RECT  1.985000  4.670000  2.235000 5.015000 ;
      RECT  1.985000  5.015000  4.015000 5.185000 ;
      RECT  2.205000  1.065000  3.475000 1.365000 ;
      RECT  2.205000  1.365000  2.535000 4.075000 ;
      RECT  2.205000  4.075000  3.475000 4.375000 ;
      RECT  2.405000  0.595000  2.735000 1.065000 ;
      RECT  2.405000  4.375000  2.735000 4.845000 ;
      RECT  2.705000  1.535000  2.975000 2.465000 ;
      RECT  2.705000  2.975000  2.975000 3.905000 ;
      RECT  2.905000  0.425000  3.075000 0.770000 ;
      RECT  2.905000  4.670000  3.075000 5.015000 ;
      RECT  3.145000  1.365000  3.475000 4.075000 ;
      RECT  3.245000  0.595000  3.575000 0.885000 ;
      RECT  3.245000  0.885000  3.475000 1.065000 ;
      RECT  3.245000  4.375000  3.475000 4.555000 ;
      RECT  3.245000  4.555000  3.575000 4.845000 ;
      RECT  3.645000  1.495000  5.875000 1.665000 ;
      RECT  3.645000  1.665000  3.945000 2.465000 ;
      RECT  3.645000  2.635000  8.775000 2.805000 ;
      RECT  3.645000  2.975000  3.945000 3.775000 ;
      RECT  3.645000  3.775000  5.875000 3.945000 ;
      RECT  3.745000  0.425000  4.015000 0.715000 ;
      RECT  3.745000  0.715000  5.875000 0.885000 ;
      RECT  3.745000  4.555000  5.875000 4.725000 ;
      RECT  3.745000  4.725000  4.015000 5.015000 ;
      RECT  4.165000  1.835000  4.435000 2.635000 ;
      RECT  4.165000  2.805000  4.435000 3.605000 ;
      RECT  4.185000  0.085000  4.435000 0.545000 ;
      RECT  4.185000  4.895000  4.435000 5.355000 ;
      RECT  4.605000  0.255000  4.935000 0.715000 ;
      RECT  4.605000  1.665000  4.935000 2.465000 ;
      RECT  4.605000  2.975000  4.935000 3.775000 ;
      RECT  4.605000  4.725000  4.935000 5.185000 ;
      RECT  5.105000  0.085000  5.375000 0.545000 ;
      RECT  5.105000  1.835000  5.375000 2.635000 ;
      RECT  5.105000  2.805000  5.375000 3.605000 ;
      RECT  5.105000  4.895000  5.375000 5.355000 ;
      RECT  5.545000  0.255000  5.875000 0.715000 ;
      RECT  5.545000  1.665000  5.875000 2.465000 ;
      RECT  5.545000  2.975000  5.875000 3.775000 ;
      RECT  5.545000  4.725000  5.875000 5.185000 ;
      RECT  6.045000  0.085000  6.375000 0.885000 ;
      RECT  6.045000  1.495000  6.375000 2.635000 ;
      RECT  6.045000  2.805000  6.375000 3.945000 ;
      RECT  6.045000  4.555000  6.375000 5.355000 ;
      RECT  6.545000  0.255000  6.875000 0.715000 ;
      RECT  6.545000  0.715000  8.675000 0.885000 ;
      RECT  6.545000  1.495000  8.775000 1.665000 ;
      RECT  6.545000  1.665000  6.875000 2.465000 ;
      RECT  6.545000  2.975000  6.875000 3.775000 ;
      RECT  6.545000  3.775000  8.775000 3.945000 ;
      RECT  6.545000  4.555000  8.675000 4.725000 ;
      RECT  6.545000  4.725000  6.875000 5.185000 ;
      RECT  7.045000  0.085000  7.315000 0.545000 ;
      RECT  7.045000  1.835000  7.315000 2.635000 ;
      RECT  7.045000  2.805000  7.315000 3.605000 ;
      RECT  7.045000  4.895000  7.315000 5.355000 ;
      RECT  7.485000  0.255000  7.815000 0.715000 ;
      RECT  7.485000  1.665000  7.815000 2.465000 ;
      RECT  7.485000  2.975000  7.815000 3.775000 ;
      RECT  7.485000  4.725000  7.815000 5.185000 ;
      RECT  7.985000  0.085000  8.235000 0.545000 ;
      RECT  7.985000  1.835000  8.255000 2.635000 ;
      RECT  7.985000  2.805000  8.255000 3.605000 ;
      RECT  7.985000  4.895000  8.235000 5.355000 ;
      RECT  8.405000  0.255000 10.435000 0.425000 ;
      RECT  8.405000  0.425000  8.675000 0.715000 ;
      RECT  8.405000  4.725000  8.675000 5.015000 ;
      RECT  8.405000  5.015000 10.435000 5.185000 ;
      RECT  8.475000  1.665000  8.775000 2.465000 ;
      RECT  8.475000  2.975000  8.775000 3.775000 ;
      RECT  8.845000  0.595000  9.175000 0.885000 ;
      RECT  8.845000  4.555000  9.175000 4.845000 ;
      RECT  8.945000  0.885000  9.175000 1.065000 ;
      RECT  8.945000  1.065000 10.215000 1.365000 ;
      RECT  8.945000  1.365000  9.275000 4.075000 ;
      RECT  8.945000  4.075000 10.215000 4.375000 ;
      RECT  8.945000  4.375000  9.175000 4.555000 ;
      RECT  9.345000  0.425000  9.515000 0.770000 ;
      RECT  9.345000  4.670000  9.515000 5.015000 ;
      RECT  9.445000  1.535000  9.715000 2.465000 ;
      RECT  9.445000  2.975000  9.715000 3.905000 ;
      RECT  9.685000  0.595000 10.015000 1.065000 ;
      RECT  9.685000  4.375000 10.015000 4.845000 ;
      RECT  9.885000  1.365000 10.215000 4.075000 ;
      RECT 10.185000  0.425000 10.435000 0.770000 ;
      RECT 10.185000  4.670000 10.435000 5.015000 ;
      RECT 10.385000  1.065000 11.570000 1.395000 ;
      RECT 10.385000  1.565000 10.685000 2.465000 ;
      RECT 10.385000  2.635000 14.455000 2.805000 ;
      RECT 10.385000  2.975000 10.685000 3.875000 ;
      RECT 10.385000  4.045000 11.570000 4.375000 ;
      RECT 10.930000  1.605000 11.205000 2.635000 ;
      RECT 10.930000  2.805000 11.205000 3.835000 ;
      RECT 10.940000  0.085000 11.230000 0.610000 ;
      RECT 10.940000  4.830000 11.230000 5.355000 ;
      RECT 11.400000  0.280000 11.650000 0.825000 ;
      RECT 11.400000  0.825000 11.570000 1.065000 ;
      RECT 11.400000  1.395000 11.570000 1.605000 ;
      RECT 11.400000  1.605000 11.730000 2.465000 ;
      RECT 11.400000  2.975000 11.730000 3.835000 ;
      RECT 11.400000  3.835000 11.570000 4.045000 ;
      RECT 11.400000  4.375000 11.570000 4.615000 ;
      RECT 11.400000  4.615000 11.650000 5.160000 ;
      RECT 11.860000  0.085000 12.150000 0.610000 ;
      RECT 11.860000  4.830000 12.150000 5.355000 ;
      RECT 11.900000  1.605000 12.200000 2.635000 ;
      RECT 11.900000  2.805000 12.200000 3.835000 ;
      RECT 12.640000  1.605000 12.940000 2.635000 ;
      RECT 12.640000  2.805000 12.940000 3.835000 ;
      RECT 12.690000  0.085000 12.980000 0.610000 ;
      RECT 12.690000  4.830000 12.980000 5.355000 ;
      RECT 13.110000  1.605000 13.440000 2.465000 ;
      RECT 13.110000  2.975000 13.440000 3.835000 ;
      RECT 13.190000  0.280000 13.440000 0.825000 ;
      RECT 13.190000  4.615000 13.440000 5.160000 ;
      RECT 13.270000  0.825000 13.440000 1.065000 ;
      RECT 13.270000  1.065000 14.455000 1.395000 ;
      RECT 13.270000  1.395000 13.440000 1.605000 ;
      RECT 13.270000  3.835000 13.440000 4.045000 ;
      RECT 13.270000  4.045000 14.455000 4.375000 ;
      RECT 13.270000  4.375000 13.440000 4.615000 ;
      RECT 13.610000  0.085000 13.900000 0.610000 ;
      RECT 13.610000  4.830000 13.900000 5.355000 ;
      RECT 13.635000  1.605000 13.910000 2.635000 ;
      RECT 13.635000  2.805000 13.910000 3.835000 ;
      RECT 14.155000  1.565000 14.455000 2.465000 ;
      RECT 14.155000  2.975000 14.455000 3.875000 ;
      RECT 14.405000  0.255000 16.435000 0.425000 ;
      RECT 14.405000  0.425000 14.655000 0.770000 ;
      RECT 14.405000  4.670000 14.655000 5.015000 ;
      RECT 14.405000  5.015000 16.435000 5.185000 ;
      RECT 14.625000  1.065000 15.895000 1.365000 ;
      RECT 14.625000  1.365000 14.955000 4.075000 ;
      RECT 14.625000  4.075000 15.895000 4.375000 ;
      RECT 14.825000  0.595000 15.155000 1.065000 ;
      RECT 14.825000  4.375000 15.155000 4.845000 ;
      RECT 15.125000  1.535000 15.395000 2.465000 ;
      RECT 15.125000  2.975000 15.395000 3.905000 ;
      RECT 15.325000  0.425000 15.495000 0.770000 ;
      RECT 15.325000  4.670000 15.495000 5.015000 ;
      RECT 15.565000  1.365000 15.895000 4.075000 ;
      RECT 15.665000  0.595000 15.995000 0.885000 ;
      RECT 15.665000  0.885000 15.895000 1.065000 ;
      RECT 15.665000  4.375000 15.895000 4.555000 ;
      RECT 15.665000  4.555000 15.995000 4.845000 ;
      RECT 16.065000  1.495000 18.295000 1.665000 ;
      RECT 16.065000  1.665000 16.365000 2.465000 ;
      RECT 16.065000  2.635000 21.195000 2.805000 ;
      RECT 16.065000  2.975000 16.365000 3.775000 ;
      RECT 16.065000  3.775000 18.295000 3.945000 ;
      RECT 16.165000  0.425000 16.435000 0.715000 ;
      RECT 16.165000  0.715000 18.295000 0.885000 ;
      RECT 16.165000  4.555000 18.295000 4.725000 ;
      RECT 16.165000  4.725000 16.435000 5.015000 ;
      RECT 16.585000  1.835000 16.855000 2.635000 ;
      RECT 16.585000  2.805000 16.855000 3.605000 ;
      RECT 16.605000  0.085000 16.855000 0.545000 ;
      RECT 16.605000  4.895000 16.855000 5.355000 ;
      RECT 17.025000  0.255000 17.355000 0.715000 ;
      RECT 17.025000  1.665000 17.355000 2.465000 ;
      RECT 17.025000  2.975000 17.355000 3.775000 ;
      RECT 17.025000  4.725000 17.355000 5.185000 ;
      RECT 17.525000  0.085000 17.795000 0.545000 ;
      RECT 17.525000  1.835000 17.795000 2.635000 ;
      RECT 17.525000  2.805000 17.795000 3.605000 ;
      RECT 17.525000  4.895000 17.795000 5.355000 ;
      RECT 17.965000  0.255000 18.295000 0.715000 ;
      RECT 17.965000  1.665000 18.295000 2.465000 ;
      RECT 17.965000  2.975000 18.295000 3.775000 ;
      RECT 17.965000  4.725000 18.295000 5.185000 ;
      RECT 18.465000  0.085000 18.795000 0.885000 ;
      RECT 18.465000  1.495000 18.795000 2.635000 ;
      RECT 18.465000  2.805000 18.795000 3.945000 ;
      RECT 18.465000  4.555000 18.795000 5.355000 ;
      RECT 18.965000  0.255000 19.295000 0.715000 ;
      RECT 18.965000  0.715000 21.095000 0.885000 ;
      RECT 18.965000  1.495000 21.195000 1.665000 ;
      RECT 18.965000  1.665000 19.295000 2.465000 ;
      RECT 18.965000  2.975000 19.295000 3.775000 ;
      RECT 18.965000  3.775000 21.195000 3.945000 ;
      RECT 18.965000  4.555000 21.095000 4.725000 ;
      RECT 18.965000  4.725000 19.295000 5.185000 ;
      RECT 19.465000  0.085000 19.735000 0.545000 ;
      RECT 19.465000  1.835000 19.735000 2.635000 ;
      RECT 19.465000  2.805000 19.735000 3.605000 ;
      RECT 19.465000  4.895000 19.735000 5.355000 ;
      RECT 19.905000  0.255000 20.235000 0.715000 ;
      RECT 19.905000  1.665000 20.235000 2.465000 ;
      RECT 19.905000  2.975000 20.235000 3.775000 ;
      RECT 19.905000  4.725000 20.235000 5.185000 ;
      RECT 20.405000  0.085000 20.655000 0.545000 ;
      RECT 20.405000  1.835000 20.675000 2.635000 ;
      RECT 20.405000  2.805000 20.675000 3.605000 ;
      RECT 20.405000  4.895000 20.655000 5.355000 ;
      RECT 20.825000  0.255000 22.855000 0.425000 ;
      RECT 20.825000  0.425000 21.095000 0.715000 ;
      RECT 20.825000  4.725000 21.095000 5.015000 ;
      RECT 20.825000  5.015000 22.855000 5.185000 ;
      RECT 20.895000  1.665000 21.195000 2.465000 ;
      RECT 20.895000  2.975000 21.195000 3.775000 ;
      RECT 21.265000  0.595000 21.595000 0.885000 ;
      RECT 21.265000  4.555000 21.595000 4.845000 ;
      RECT 21.365000  0.885000 21.595000 1.065000 ;
      RECT 21.365000  1.065000 22.635000 1.365000 ;
      RECT 21.365000  1.365000 21.695000 4.075000 ;
      RECT 21.365000  4.075000 22.635000 4.375000 ;
      RECT 21.365000  4.375000 21.595000 4.555000 ;
      RECT 21.765000  0.425000 21.935000 0.770000 ;
      RECT 21.765000  4.670000 21.935000 5.015000 ;
      RECT 21.865000  1.535000 22.135000 2.465000 ;
      RECT 21.865000  2.975000 22.135000 3.905000 ;
      RECT 22.105000  0.595000 22.435000 1.065000 ;
      RECT 22.105000  4.375000 22.435000 4.845000 ;
      RECT 22.305000  1.365000 22.635000 4.075000 ;
      RECT 22.605000  0.425000 22.855000 0.770000 ;
      RECT 22.605000  4.670000 22.855000 5.015000 ;
      RECT 22.805000  1.065000 23.990000 1.395000 ;
      RECT 22.805000  1.565000 23.105000 2.465000 ;
      RECT 22.805000  2.635000 24.840000 2.805000 ;
      RECT 22.805000  2.975000 23.105000 3.875000 ;
      RECT 22.805000  4.045000 23.990000 4.375000 ;
      RECT 23.350000  1.605000 23.625000 2.635000 ;
      RECT 23.350000  2.805000 23.625000 3.835000 ;
      RECT 23.360000  0.085000 23.650000 0.610000 ;
      RECT 23.360000  4.830000 23.650000 5.355000 ;
      RECT 23.820000  0.280000 24.070000 0.825000 ;
      RECT 23.820000  0.825000 23.990000 1.065000 ;
      RECT 23.820000  1.395000 23.990000 1.605000 ;
      RECT 23.820000  1.605000 24.150000 2.465000 ;
      RECT 23.820000  2.975000 24.150000 3.835000 ;
      RECT 23.820000  3.835000 23.990000 4.045000 ;
      RECT 23.820000  4.375000 23.990000 4.615000 ;
      RECT 23.820000  4.615000 24.070000 5.160000 ;
      RECT 24.280000  0.085000 24.570000 0.610000 ;
      RECT 24.280000  4.830000 24.570000 5.355000 ;
      RECT 24.320000  1.605000 24.620000 2.635000 ;
      RECT 24.320000  2.805000 24.620000 3.835000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.145000  5.355000  0.315000 5.525000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.605000  5.355000  0.775000 5.525000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.065000  5.355000  1.235000 5.525000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.525000  5.355000  1.695000 5.525000 ;
      RECT  1.805000  2.140000  1.975000 2.310000 ;
      RECT  1.805000  3.130000  1.975000 3.300000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  5.355000  2.155000 5.525000 ;
      RECT  2.285000  1.785000  2.455000 1.955000 ;
      RECT  2.285000  3.485000  2.455000 3.655000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  5.355000  2.615000 5.525000 ;
      RECT  2.755000  2.140000  2.925000 2.310000 ;
      RECT  2.755000  3.130000  2.925000 3.300000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  5.355000  3.075000 5.525000 ;
      RECT  3.225000  1.785000  3.395000 1.955000 ;
      RECT  3.225000  3.485000  3.395000 3.655000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  5.355000  3.535000 5.525000 ;
      RECT  3.705000  2.140000  3.875000 2.310000 ;
      RECT  3.705000  3.130000  3.875000 3.300000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  3.825000  5.355000  3.995000 5.525000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.285000  5.355000  4.455000 5.525000 ;
      RECT  4.685000  2.140000  4.855000 2.310000 ;
      RECT  4.685000  3.130000  4.855000 3.300000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.745000  5.355000  4.915000 5.525000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.205000  5.355000  5.375000 5.525000 ;
      RECT  5.625000  2.140000  5.795000 2.310000 ;
      RECT  5.625000  3.130000  5.795000 3.300000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.665000  5.355000  5.835000 5.525000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.125000  5.355000  6.295000 5.525000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.585000  5.355000  6.755000 5.525000 ;
      RECT  6.625000  2.140000  6.795000 2.310000 ;
      RECT  6.625000  3.130000  6.795000 3.300000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.045000  5.355000  7.215000 5.525000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.505000  5.355000  7.675000 5.525000 ;
      RECT  7.565000  2.140000  7.735000 2.310000 ;
      RECT  7.565000  3.130000  7.735000 3.300000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  7.965000  5.355000  8.135000 5.525000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.425000  5.355000  8.595000 5.525000 ;
      RECT  8.545000  2.140000  8.715000 2.310000 ;
      RECT  8.545000  3.130000  8.715000 3.300000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  5.355000  9.055000 5.525000 ;
      RECT  9.025000  1.785000  9.195000 1.955000 ;
      RECT  9.025000  3.485000  9.195000 3.655000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  5.355000  9.515000 5.525000 ;
      RECT  9.495000  2.140000  9.665000 2.310000 ;
      RECT  9.495000  3.130000  9.665000 3.300000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  5.355000  9.975000 5.525000 ;
      RECT  9.965000  1.785000 10.135000 1.955000 ;
      RECT  9.965000  3.485000 10.135000 3.655000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  5.355000 10.435000 5.525000 ;
      RECT 10.445000  2.140000 10.615000 2.310000 ;
      RECT 10.445000  3.130000 10.615000 3.300000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.725000  5.355000 10.895000 5.525000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.185000  5.355000 11.355000 5.525000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 11.645000  5.355000 11.815000 5.525000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.105000  5.355000 12.275000 5.525000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 12.565000  5.355000 12.735000 5.525000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.025000  5.355000 13.195000 5.525000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.485000  5.355000 13.655000 5.525000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 13.945000  5.355000 14.115000 5.525000 ;
      RECT 14.225000  2.140000 14.395000 2.310000 ;
      RECT 14.225000  3.130000 14.395000 3.300000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  5.355000 14.575000 5.525000 ;
      RECT 14.705000  1.785000 14.875000 1.955000 ;
      RECT 14.705000  3.485000 14.875000 3.655000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  5.355000 15.035000 5.525000 ;
      RECT 15.175000  2.140000 15.345000 2.310000 ;
      RECT 15.175000  3.130000 15.345000 3.300000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  5.355000 15.495000 5.525000 ;
      RECT 15.645000  1.785000 15.815000 1.955000 ;
      RECT 15.645000  3.485000 15.815000 3.655000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  5.355000 15.955000 5.525000 ;
      RECT 16.125000  2.140000 16.295000 2.310000 ;
      RECT 16.125000  3.130000 16.295000 3.300000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.245000  5.355000 16.415000 5.525000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
      RECT 16.705000  5.355000 16.875000 5.525000 ;
      RECT 17.105000  2.140000 17.275000 2.310000 ;
      RECT 17.105000  3.130000 17.275000 3.300000 ;
      RECT 17.165000 -0.085000 17.335000 0.085000 ;
      RECT 17.165000  2.635000 17.335000 2.805000 ;
      RECT 17.165000  5.355000 17.335000 5.525000 ;
      RECT 17.625000 -0.085000 17.795000 0.085000 ;
      RECT 17.625000  2.635000 17.795000 2.805000 ;
      RECT 17.625000  5.355000 17.795000 5.525000 ;
      RECT 18.045000  2.140000 18.215000 2.310000 ;
      RECT 18.045000  3.130000 18.215000 3.300000 ;
      RECT 18.085000 -0.085000 18.255000 0.085000 ;
      RECT 18.085000  2.635000 18.255000 2.805000 ;
      RECT 18.085000  5.355000 18.255000 5.525000 ;
      RECT 18.545000 -0.085000 18.715000 0.085000 ;
      RECT 18.545000  2.635000 18.715000 2.805000 ;
      RECT 18.545000  5.355000 18.715000 5.525000 ;
      RECT 19.005000 -0.085000 19.175000 0.085000 ;
      RECT 19.005000  2.635000 19.175000 2.805000 ;
      RECT 19.005000  5.355000 19.175000 5.525000 ;
      RECT 19.045000  2.140000 19.215000 2.310000 ;
      RECT 19.045000  3.130000 19.215000 3.300000 ;
      RECT 19.465000 -0.085000 19.635000 0.085000 ;
      RECT 19.465000  2.635000 19.635000 2.805000 ;
      RECT 19.465000  5.355000 19.635000 5.525000 ;
      RECT 19.925000 -0.085000 20.095000 0.085000 ;
      RECT 19.925000  2.635000 20.095000 2.805000 ;
      RECT 19.925000  5.355000 20.095000 5.525000 ;
      RECT 19.985000  2.140000 20.155000 2.310000 ;
      RECT 19.985000  3.130000 20.155000 3.300000 ;
      RECT 20.385000 -0.085000 20.555000 0.085000 ;
      RECT 20.385000  2.635000 20.555000 2.805000 ;
      RECT 20.385000  5.355000 20.555000 5.525000 ;
      RECT 20.845000 -0.085000 21.015000 0.085000 ;
      RECT 20.845000  2.635000 21.015000 2.805000 ;
      RECT 20.845000  5.355000 21.015000 5.525000 ;
      RECT 20.965000  2.140000 21.135000 2.310000 ;
      RECT 20.965000  3.130000 21.135000 3.300000 ;
      RECT 21.305000 -0.085000 21.475000 0.085000 ;
      RECT 21.305000  5.355000 21.475000 5.525000 ;
      RECT 21.445000  1.785000 21.615000 1.955000 ;
      RECT 21.445000  3.485000 21.615000 3.655000 ;
      RECT 21.765000 -0.085000 21.935000 0.085000 ;
      RECT 21.765000  5.355000 21.935000 5.525000 ;
      RECT 21.915000  2.140000 22.085000 2.310000 ;
      RECT 21.915000  3.130000 22.085000 3.300000 ;
      RECT 22.225000 -0.085000 22.395000 0.085000 ;
      RECT 22.225000  5.355000 22.395000 5.525000 ;
      RECT 22.385000  1.785000 22.555000 1.955000 ;
      RECT 22.385000  3.485000 22.555000 3.655000 ;
      RECT 22.685000 -0.085000 22.855000 0.085000 ;
      RECT 22.685000  5.355000 22.855000 5.525000 ;
      RECT 22.865000  2.140000 23.035000 2.310000 ;
      RECT 22.865000  3.130000 23.035000 3.300000 ;
      RECT 23.145000 -0.085000 23.315000 0.085000 ;
      RECT 23.145000  2.635000 23.315000 2.805000 ;
      RECT 23.145000  5.355000 23.315000 5.525000 ;
      RECT 23.605000 -0.085000 23.775000 0.085000 ;
      RECT 23.605000  2.635000 23.775000 2.805000 ;
      RECT 23.605000  5.355000 23.775000 5.525000 ;
      RECT 24.065000 -0.085000 24.235000 0.085000 ;
      RECT 24.065000  2.635000 24.235000 2.805000 ;
      RECT 24.065000  5.355000 24.235000 5.525000 ;
      RECT 24.525000 -0.085000 24.695000 0.085000 ;
      RECT 24.525000  2.635000 24.695000 2.805000 ;
      RECT 24.525000  5.355000 24.695000 5.525000 ;
    LAYER met1 ;
      RECT  1.745000 2.110000  2.035000 2.155000 ;
      RECT  1.745000 2.155000  5.855000 2.295000 ;
      RECT  1.745000 2.295000  2.035000 2.340000 ;
      RECT  1.745000 3.100000  2.035000 3.145000 ;
      RECT  1.745000 3.145000  5.855000 3.285000 ;
      RECT  1.745000 3.285000  2.035000 3.330000 ;
      RECT  2.695000 2.110000  2.985000 2.155000 ;
      RECT  2.695000 2.295000  2.985000 2.340000 ;
      RECT  2.695000 3.100000  2.985000 3.145000 ;
      RECT  2.695000 3.285000  2.985000 3.330000 ;
      RECT  3.645000 2.110000  3.935000 2.155000 ;
      RECT  3.645000 2.295000  3.935000 2.340000 ;
      RECT  3.645000 3.100000  3.935000 3.145000 ;
      RECT  3.645000 3.285000  3.935000 3.330000 ;
      RECT  4.625000 2.110000  4.915000 2.155000 ;
      RECT  4.625000 2.295000  4.915000 2.340000 ;
      RECT  4.625000 3.100000  4.915000 3.145000 ;
      RECT  4.625000 3.285000  4.915000 3.330000 ;
      RECT  5.565000 2.110000  5.855000 2.155000 ;
      RECT  5.565000 2.295000  5.855000 2.340000 ;
      RECT  5.565000 3.100000  5.855000 3.145000 ;
      RECT  5.565000 3.285000  5.855000 3.330000 ;
      RECT  6.565000 2.110000  6.855000 2.155000 ;
      RECT  6.565000 2.155000 10.675000 2.295000 ;
      RECT  6.565000 2.295000  6.855000 2.340000 ;
      RECT  6.565000 3.100000  6.855000 3.145000 ;
      RECT  6.565000 3.145000 10.675000 3.285000 ;
      RECT  6.565000 3.285000  6.855000 3.330000 ;
      RECT  7.505000 2.110000  7.795000 2.155000 ;
      RECT  7.505000 2.295000  7.795000 2.340000 ;
      RECT  7.505000 3.100000  7.795000 3.145000 ;
      RECT  7.505000 3.285000  7.795000 3.330000 ;
      RECT  8.485000 2.110000  8.775000 2.155000 ;
      RECT  8.485000 2.295000  8.775000 2.340000 ;
      RECT  8.485000 3.100000  8.775000 3.145000 ;
      RECT  8.485000 3.285000  8.775000 3.330000 ;
      RECT  9.435000 2.110000  9.725000 2.155000 ;
      RECT  9.435000 2.295000  9.725000 2.340000 ;
      RECT  9.435000 3.100000  9.725000 3.145000 ;
      RECT  9.435000 3.285000  9.725000 3.330000 ;
      RECT 10.385000 2.110000 10.675000 2.155000 ;
      RECT 10.385000 2.295000 10.675000 2.340000 ;
      RECT 10.385000 3.100000 10.675000 3.145000 ;
      RECT 10.385000 3.285000 10.675000 3.330000 ;
      RECT 14.165000 2.110000 14.455000 2.155000 ;
      RECT 14.165000 2.155000 18.275000 2.295000 ;
      RECT 14.165000 2.295000 14.455000 2.340000 ;
      RECT 14.165000 3.100000 14.455000 3.145000 ;
      RECT 14.165000 3.145000 18.275000 3.285000 ;
      RECT 14.165000 3.285000 14.455000 3.330000 ;
      RECT 15.115000 2.110000 15.405000 2.155000 ;
      RECT 15.115000 2.295000 15.405000 2.340000 ;
      RECT 15.115000 3.100000 15.405000 3.145000 ;
      RECT 15.115000 3.285000 15.405000 3.330000 ;
      RECT 16.065000 2.110000 16.355000 2.155000 ;
      RECT 16.065000 2.295000 16.355000 2.340000 ;
      RECT 16.065000 3.100000 16.355000 3.145000 ;
      RECT 16.065000 3.285000 16.355000 3.330000 ;
      RECT 17.045000 2.110000 17.335000 2.155000 ;
      RECT 17.045000 2.295000 17.335000 2.340000 ;
      RECT 17.045000 3.100000 17.335000 3.145000 ;
      RECT 17.045000 3.285000 17.335000 3.330000 ;
      RECT 17.985000 2.110000 18.275000 2.155000 ;
      RECT 17.985000 2.295000 18.275000 2.340000 ;
      RECT 17.985000 3.100000 18.275000 3.145000 ;
      RECT 17.985000 3.285000 18.275000 3.330000 ;
      RECT 18.985000 2.110000 19.275000 2.155000 ;
      RECT 18.985000 2.155000 23.095000 2.295000 ;
      RECT 18.985000 2.295000 19.275000 2.340000 ;
      RECT 18.985000 3.100000 19.275000 3.145000 ;
      RECT 18.985000 3.145000 23.095000 3.285000 ;
      RECT 18.985000 3.285000 19.275000 3.330000 ;
      RECT 19.925000 2.110000 20.215000 2.155000 ;
      RECT 19.925000 2.295000 20.215000 2.340000 ;
      RECT 19.925000 3.100000 20.215000 3.145000 ;
      RECT 19.925000 3.285000 20.215000 3.330000 ;
      RECT 20.905000 2.110000 21.195000 2.155000 ;
      RECT 20.905000 2.295000 21.195000 2.340000 ;
      RECT 20.905000 3.100000 21.195000 3.145000 ;
      RECT 20.905000 3.285000 21.195000 3.330000 ;
      RECT 21.855000 2.110000 22.145000 2.155000 ;
      RECT 21.855000 2.295000 22.145000 2.340000 ;
      RECT 21.855000 3.100000 22.145000 3.145000 ;
      RECT 21.855000 3.285000 22.145000 3.330000 ;
      RECT 22.805000 2.110000 23.095000 2.155000 ;
      RECT 22.805000 2.295000 23.095000 2.340000 ;
      RECT 22.805000 3.100000 23.095000 3.145000 ;
      RECT 22.805000 3.285000 23.095000 3.330000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb8to1_4


MACRO sky130_fd_sc_hdll__muxb8to1_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  17.02000 BY  2.720000 ;
  SITE unithd ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.335000 1.055000 0.730000 1.325000 ;
        RECT 0.560000 0.395000 0.835000 0.625000 ;
        RECT 0.560000 0.625000 0.730000 1.055000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 0.395000 4.040000 0.625000 ;
        RECT 3.870000 0.625000 4.040000 1.055000 ;
        RECT 3.870000 1.055000 4.265000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 1.055000 4.870000 1.325000 ;
        RECT 4.700000 0.395000 4.975000 0.625000 ;
        RECT 4.700000 0.625000 4.870000 1.055000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.905000 0.395000 8.180000 0.625000 ;
        RECT 8.010000 0.625000 8.180000 1.055000 ;
        RECT 8.010000 1.055000 8.405000 1.325000 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.615000 1.055000 9.010000 1.325000 ;
        RECT 8.840000 0.395000 9.115000 0.625000 ;
        RECT 8.840000 0.625000 9.010000 1.055000 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.045000 0.395000 12.320000 0.625000 ;
        RECT 12.150000 0.625000 12.320000 1.055000 ;
        RECT 12.150000 1.055000 12.545000 1.325000 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755000 1.055000 13.150000 1.325000 ;
        RECT 12.980000 0.395000 13.255000 0.625000 ;
        RECT 12.980000 0.625000 13.150000 1.055000 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.185000 0.395000 16.460000 0.625000 ;
        RECT 16.290000 0.625000 16.460000 1.055000 ;
        RECT 16.290000 1.055000 16.685000 1.325000 ;
    END
  END D[7]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 0.945000 2.205000 1.295000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.395000 0.945000 2.795000 1.295000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.945000 0.945000 6.345000 1.295000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 0.945000 6.935000 1.295000 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.085000 0.945000 10.485000 1.295000 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.675000 0.945000 11.075000 1.295000 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.225000 0.945000 14.625000 1.295000 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.815000 0.945000 15.215000 1.295000 ;
    END
  END S[7]
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  1.005000 1.755000  1.295000 1.800000 ;
        RECT  1.005000 1.800000 16.015000 1.940000 ;
        RECT  1.005000 1.940000  1.295000 1.985000 ;
        RECT  3.305000 1.755000  3.595000 1.800000 ;
        RECT  3.305000 1.940000  3.595000 1.985000 ;
        RECT  5.145000 1.755000  5.435000 1.800000 ;
        RECT  5.145000 1.940000  5.435000 1.985000 ;
        RECT  7.445000 1.755000  7.735000 1.800000 ;
        RECT  7.445000 1.940000  7.735000 1.985000 ;
        RECT  9.285000 1.755000  9.575000 1.800000 ;
        RECT  9.285000 1.940000  9.575000 1.985000 ;
        RECT 11.585000 1.755000 11.875000 1.800000 ;
        RECT 11.585000 1.940000 11.875000 1.985000 ;
        RECT 13.425000 1.755000 13.715000 1.800000 ;
        RECT 13.425000 1.940000 13.715000 1.985000 ;
        RECT 15.725000 1.755000 16.015000 1.800000 ;
        RECT 15.725000 1.940000 16.015000 1.985000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 17.020000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 17.020000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 17.020000 0.085000 ;
      RECT  0.000000  2.635000 17.020000 2.805000 ;
      RECT  0.095000  1.495000  0.425000 2.635000 ;
      RECT  0.130000  0.085000  0.390000 0.885000 ;
      RECT  0.900000  0.835000  1.290000 1.005000 ;
      RECT  0.900000  1.005000  1.070000 1.755000 ;
      RECT  0.900000  1.755000  1.295000 1.805000 ;
      RECT  0.900000  1.805000  1.420000 1.985000 ;
      RECT  1.045000  0.330000  1.290000 0.835000 ;
      RECT  1.090000  1.985000  1.420000 2.465000 ;
      RECT  1.240000  1.175000  1.630000 1.465000 ;
      RECT  1.240000  1.465000  1.940000 1.505000 ;
      RECT  1.460000  0.585000  1.900000 0.755000 ;
      RECT  1.460000  0.755000  1.630000 1.175000 ;
      RECT  1.460000  1.505000  1.940000 1.635000 ;
      RECT  1.610000  1.635000  1.940000 2.465000 ;
      RECT  1.650000  0.330000  1.900000 0.585000 ;
      RECT  2.135000  0.085000  2.465000 0.660000 ;
      RECT  2.135000  1.465000  2.465000 2.635000 ;
      RECT  2.660000  1.465000  3.360000 1.505000 ;
      RECT  2.660000  1.505000  3.140000 1.635000 ;
      RECT  2.660000  1.635000  2.990000 2.465000 ;
      RECT  2.700000  0.330000  2.950000 0.585000 ;
      RECT  2.700000  0.585000  3.140000 0.755000 ;
      RECT  2.970000  0.755000  3.140000 1.175000 ;
      RECT  2.970000  1.175000  3.360000 1.465000 ;
      RECT  3.180000  1.805000  3.700000 1.985000 ;
      RECT  3.180000  1.985000  3.510000 2.465000 ;
      RECT  3.305000  1.755000  3.700000 1.805000 ;
      RECT  3.310000  0.330000  3.555000 0.835000 ;
      RECT  3.310000  0.835000  3.700000 1.005000 ;
      RECT  3.530000  1.005000  3.700000 1.755000 ;
      RECT  4.175000  1.495000  4.565000 2.635000 ;
      RECT  4.210000  0.085000  4.530000 0.885000 ;
      RECT  5.040000  0.835000  5.430000 1.005000 ;
      RECT  5.040000  1.005000  5.210000 1.755000 ;
      RECT  5.040000  1.755000  5.435000 1.805000 ;
      RECT  5.040000  1.805000  5.560000 1.985000 ;
      RECT  5.185000  0.330000  5.430000 0.835000 ;
      RECT  5.230000  1.985000  5.560000 2.465000 ;
      RECT  5.380000  1.175000  5.770000 1.465000 ;
      RECT  5.380000  1.465000  6.080000 1.505000 ;
      RECT  5.600000  0.585000  6.040000 0.755000 ;
      RECT  5.600000  0.755000  5.770000 1.175000 ;
      RECT  5.600000  1.505000  6.080000 1.635000 ;
      RECT  5.750000  1.635000  6.080000 2.465000 ;
      RECT  5.790000  0.330000  6.040000 0.585000 ;
      RECT  6.275000  0.085000  6.605000 0.660000 ;
      RECT  6.275000  1.465000  6.605000 2.635000 ;
      RECT  6.800000  1.465000  7.500000 1.505000 ;
      RECT  6.800000  1.505000  7.280000 1.635000 ;
      RECT  6.800000  1.635000  7.130000 2.465000 ;
      RECT  6.840000  0.330000  7.090000 0.585000 ;
      RECT  6.840000  0.585000  7.280000 0.755000 ;
      RECT  7.110000  0.755000  7.280000 1.175000 ;
      RECT  7.110000  1.175000  7.500000 1.465000 ;
      RECT  7.320000  1.805000  7.840000 1.985000 ;
      RECT  7.320000  1.985000  7.650000 2.465000 ;
      RECT  7.445000  1.755000  7.840000 1.805000 ;
      RECT  7.450000  0.330000  7.695000 0.835000 ;
      RECT  7.450000  0.835000  7.840000 1.005000 ;
      RECT  7.670000  1.005000  7.840000 1.755000 ;
      RECT  8.315000  1.495000  8.705000 2.635000 ;
      RECT  8.350000  0.085000  8.670000 0.885000 ;
      RECT  9.180000  0.835000  9.570000 1.005000 ;
      RECT  9.180000  1.005000  9.350000 1.755000 ;
      RECT  9.180000  1.755000  9.575000 1.805000 ;
      RECT  9.180000  1.805000  9.700000 1.985000 ;
      RECT  9.325000  0.330000  9.570000 0.835000 ;
      RECT  9.370000  1.985000  9.700000 2.465000 ;
      RECT  9.520000  1.175000  9.910000 1.465000 ;
      RECT  9.520000  1.465000 10.220000 1.505000 ;
      RECT  9.740000  0.585000 10.180000 0.755000 ;
      RECT  9.740000  0.755000  9.910000 1.175000 ;
      RECT  9.740000  1.505000 10.220000 1.635000 ;
      RECT  9.890000  1.635000 10.220000 2.465000 ;
      RECT  9.930000  0.330000 10.180000 0.585000 ;
      RECT 10.415000  0.085000 10.745000 0.660000 ;
      RECT 10.415000  1.465000 10.745000 2.635000 ;
      RECT 10.940000  1.465000 11.640000 1.505000 ;
      RECT 10.940000  1.505000 11.420000 1.635000 ;
      RECT 10.940000  1.635000 11.270000 2.465000 ;
      RECT 10.980000  0.330000 11.230000 0.585000 ;
      RECT 10.980000  0.585000 11.420000 0.755000 ;
      RECT 11.250000  0.755000 11.420000 1.175000 ;
      RECT 11.250000  1.175000 11.640000 1.465000 ;
      RECT 11.460000  1.805000 11.980000 1.985000 ;
      RECT 11.460000  1.985000 11.790000 2.465000 ;
      RECT 11.585000  1.755000 11.980000 1.805000 ;
      RECT 11.590000  0.330000 11.835000 0.835000 ;
      RECT 11.590000  0.835000 11.980000 1.005000 ;
      RECT 11.810000  1.005000 11.980000 1.755000 ;
      RECT 12.455000  1.495000 12.845000 2.635000 ;
      RECT 12.490000  0.085000 12.810000 0.885000 ;
      RECT 13.320000  0.835000 13.710000 1.005000 ;
      RECT 13.320000  1.005000 13.490000 1.755000 ;
      RECT 13.320000  1.755000 13.715000 1.805000 ;
      RECT 13.320000  1.805000 13.840000 1.985000 ;
      RECT 13.465000  0.330000 13.710000 0.835000 ;
      RECT 13.510000  1.985000 13.840000 2.465000 ;
      RECT 13.660000  1.175000 14.050000 1.465000 ;
      RECT 13.660000  1.465000 14.360000 1.505000 ;
      RECT 13.880000  0.585000 14.320000 0.755000 ;
      RECT 13.880000  0.755000 14.050000 1.175000 ;
      RECT 13.880000  1.505000 14.360000 1.635000 ;
      RECT 14.030000  1.635000 14.360000 2.465000 ;
      RECT 14.070000  0.330000 14.320000 0.585000 ;
      RECT 14.555000  0.085000 14.885000 0.660000 ;
      RECT 14.555000  1.465000 14.885000 2.635000 ;
      RECT 15.080000  1.465000 15.780000 1.505000 ;
      RECT 15.080000  1.505000 15.560000 1.635000 ;
      RECT 15.080000  1.635000 15.410000 2.465000 ;
      RECT 15.120000  0.330000 15.370000 0.585000 ;
      RECT 15.120000  0.585000 15.560000 0.755000 ;
      RECT 15.390000  0.755000 15.560000 1.175000 ;
      RECT 15.390000  1.175000 15.780000 1.465000 ;
      RECT 15.600000  1.805000 16.120000 1.985000 ;
      RECT 15.600000  1.985000 15.930000 2.465000 ;
      RECT 15.725000  1.755000 16.120000 1.805000 ;
      RECT 15.730000  0.330000 15.975000 0.835000 ;
      RECT 15.730000  0.835000 16.120000 1.005000 ;
      RECT 15.950000  1.005000 16.120000 1.755000 ;
      RECT 16.595000  1.495000 16.925000 2.635000 ;
      RECT 16.630000  0.085000 16.890000 0.885000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  1.785000  1.235000 1.955000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  1.785000  3.535000 1.955000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  1.785000  7.675000 1.955000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  1.785000  9.515000 1.955000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  1.785000 11.815000 1.955000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  1.785000 13.655000 1.955000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  1.785000 15.955000 1.955000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb8to1_1


MACRO sky130_fd_sc_hdll__muxb8to1_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  25.76000 BY  2.720000 ;
  SITE unithd ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.055000 0.915000 1.325000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.525000 1.055000 6.345000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 1.055000 7.355000 1.325000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.965000 1.055000 12.785000 1.325000 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.975000 1.055000 13.795000 1.325000 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.405000 1.055000 19.225000 1.325000 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.415000 1.055000 20.235000 1.325000 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.845000 1.055000 25.665000 1.325000 ;
    END
  END D[7]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 1.025000 3.125000 1.295000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.025000 3.650000 1.295000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.230000 1.025000 9.565000 1.295000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.755000 1.025000 10.090000 1.295000 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.670000 1.025000 16.005000 1.295000 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.195000 1.025000 16.530000 1.295000 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.110000 1.025000 22.445000 1.295000 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.635000 1.025000 22.970000 1.295000 ;
    END
  END S[7]
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  1.465000 1.755000  1.755000 1.800000 ;
        RECT  1.465000 1.800000 24.295000 1.940000 ;
        RECT  1.465000 1.940000  1.755000 1.985000 ;
        RECT  4.685000 1.755000  4.975000 1.800000 ;
        RECT  4.685000 1.940000  4.975000 1.985000 ;
        RECT  7.905000 1.755000  8.195000 1.800000 ;
        RECT  7.905000 1.940000  8.195000 1.985000 ;
        RECT 11.125000 1.755000 11.415000 1.800000 ;
        RECT 11.125000 1.940000 11.415000 1.985000 ;
        RECT 14.345000 1.755000 14.635000 1.800000 ;
        RECT 14.345000 1.940000 14.635000 1.985000 ;
        RECT 17.565000 1.755000 17.855000 1.800000 ;
        RECT 17.565000 1.940000 17.855000 1.985000 ;
        RECT 20.785000 1.755000 21.075000 1.800000 ;
        RECT 20.785000 1.940000 21.075000 1.985000 ;
        RECT 24.005000 1.755000 24.295000 1.800000 ;
        RECT 24.005000 1.940000 24.295000 1.985000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 25.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 25.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 25.760000 0.085000 ;
      RECT  0.000000  2.635000 25.760000 2.805000 ;
      RECT  0.095000  1.495000  1.285000 1.665000 ;
      RECT  0.095000  1.665000  0.395000 2.210000 ;
      RECT  0.095000  2.210000  0.425000 2.465000 ;
      RECT  0.145000  0.255000  0.475000 0.715000 ;
      RECT  0.145000  0.715000  1.335000 0.885000 ;
      RECT  0.565000  1.835000  0.895000 2.105000 ;
      RECT  0.595000  2.105000  0.895000 2.635000 ;
      RECT  0.645000  0.085000  0.860000 0.545000 ;
      RECT  1.030000  0.255000  2.175000 0.425000 ;
      RECT  1.030000  0.425000  1.335000 0.715000 ;
      RECT  1.030000  0.885000  1.335000 0.925000 ;
      RECT  1.115000  1.665000  1.285000 2.295000 ;
      RECT  1.115000  2.295000  2.280000 2.465000 ;
      RECT  1.465000  1.755000  1.895000 2.125000 ;
      RECT  1.505000  0.595000  1.835000 0.885000 ;
      RECT  1.585000  0.885000  1.755000 1.755000 ;
      RECT  2.005000  0.425000  2.175000 0.770000 ;
      RECT  2.100000  1.205000  2.515000 1.305000 ;
      RECT  2.100000  1.305000  2.620000 1.465000 ;
      RECT  2.100000  1.465000  2.880000 1.475000 ;
      RECT  2.110000  1.645000  2.280000 2.295000 ;
      RECT  2.345000  0.585000  2.925000 0.755000 ;
      RECT  2.345000  0.755000  2.515000 1.205000 ;
      RECT  2.450000  1.475000  2.880000 1.635000 ;
      RECT  2.550000  1.635000  2.880000 2.465000 ;
      RECT  2.675000  0.330000  2.925000 0.585000 ;
      RECT  3.055000  1.465000  3.385000 2.635000 ;
      RECT  3.095000  0.085000  3.345000 0.660000 ;
      RECT  3.515000  0.330000  3.765000 0.585000 ;
      RECT  3.515000  0.585000  4.095000 0.755000 ;
      RECT  3.560000  1.465000  4.340000 1.475000 ;
      RECT  3.560000  1.475000  3.990000 1.635000 ;
      RECT  3.560000  1.635000  3.890000 2.465000 ;
      RECT  3.820000  1.305000  4.340000 1.465000 ;
      RECT  3.925000  0.755000  4.095000 1.205000 ;
      RECT  3.925000  1.205000  4.340000 1.305000 ;
      RECT  4.160000  1.645000  4.330000 2.295000 ;
      RECT  4.160000  2.295000  5.325000 2.465000 ;
      RECT  4.265000  0.255000  5.410000 0.425000 ;
      RECT  4.265000  0.425000  4.435000 0.770000 ;
      RECT  4.545000  1.755000  4.975000 2.125000 ;
      RECT  4.605000  0.595000  4.935000 0.885000 ;
      RECT  4.685000  0.885000  4.855000 1.755000 ;
      RECT  5.105000  0.425000  5.410000 0.715000 ;
      RECT  5.105000  0.715000  6.295000 0.885000 ;
      RECT  5.105000  0.885000  5.410000 0.925000 ;
      RECT  5.155000  1.495000  6.345000 1.665000 ;
      RECT  5.155000  1.665000  5.325000 2.295000 ;
      RECT  5.545000  1.835000  5.875000 2.105000 ;
      RECT  5.545000  2.105000  5.845000 2.635000 ;
      RECT  5.580000  0.085000  5.795000 0.545000 ;
      RECT  5.965000  0.255000  6.295000 0.715000 ;
      RECT  6.015000  2.210000  6.345000 2.465000 ;
      RECT  6.045000  1.665000  6.345000 2.210000 ;
      RECT  6.535000  1.495000  7.725000 1.665000 ;
      RECT  6.535000  1.665000  6.835000 2.210000 ;
      RECT  6.535000  2.210000  6.865000 2.465000 ;
      RECT  6.585000  0.255000  6.915000 0.715000 ;
      RECT  6.585000  0.715000  7.775000 0.885000 ;
      RECT  7.005000  1.835000  7.335000 2.105000 ;
      RECT  7.035000  2.105000  7.335000 2.635000 ;
      RECT  7.085000  0.085000  7.300000 0.545000 ;
      RECT  7.470000  0.255000  8.615000 0.425000 ;
      RECT  7.470000  0.425000  7.775000 0.715000 ;
      RECT  7.470000  0.885000  7.775000 0.925000 ;
      RECT  7.555000  1.665000  7.725000 2.295000 ;
      RECT  7.555000  2.295000  8.720000 2.465000 ;
      RECT  7.905000  1.755000  8.335000 2.125000 ;
      RECT  7.945000  0.595000  8.275000 0.885000 ;
      RECT  8.025000  0.885000  8.195000 1.755000 ;
      RECT  8.445000  0.425000  8.615000 0.770000 ;
      RECT  8.540000  1.205000  8.955000 1.305000 ;
      RECT  8.540000  1.305000  9.060000 1.465000 ;
      RECT  8.540000  1.465000  9.320000 1.475000 ;
      RECT  8.550000  1.645000  8.720000 2.295000 ;
      RECT  8.785000  0.585000  9.365000 0.755000 ;
      RECT  8.785000  0.755000  8.955000 1.205000 ;
      RECT  8.890000  1.475000  9.320000 1.635000 ;
      RECT  8.990000  1.635000  9.320000 2.465000 ;
      RECT  9.115000  0.330000  9.365000 0.585000 ;
      RECT  9.495000  1.465000  9.825000 2.635000 ;
      RECT  9.535000  0.085000  9.785000 0.660000 ;
      RECT  9.955000  0.330000 10.205000 0.585000 ;
      RECT  9.955000  0.585000 10.535000 0.755000 ;
      RECT 10.000000  1.465000 10.780000 1.475000 ;
      RECT 10.000000  1.475000 10.430000 1.635000 ;
      RECT 10.000000  1.635000 10.330000 2.465000 ;
      RECT 10.260000  1.305000 10.780000 1.465000 ;
      RECT 10.365000  0.755000 10.535000 1.205000 ;
      RECT 10.365000  1.205000 10.780000 1.305000 ;
      RECT 10.600000  1.645000 10.770000 2.295000 ;
      RECT 10.600000  2.295000 11.765000 2.465000 ;
      RECT 10.705000  0.255000 11.850000 0.425000 ;
      RECT 10.705000  0.425000 10.875000 0.770000 ;
      RECT 10.985000  1.755000 11.415000 2.125000 ;
      RECT 11.045000  0.595000 11.375000 0.885000 ;
      RECT 11.125000  0.885000 11.295000 1.755000 ;
      RECT 11.545000  0.425000 11.850000 0.715000 ;
      RECT 11.545000  0.715000 12.735000 0.885000 ;
      RECT 11.545000  0.885000 11.850000 0.925000 ;
      RECT 11.595000  1.495000 12.785000 1.665000 ;
      RECT 11.595000  1.665000 11.765000 2.295000 ;
      RECT 11.985000  1.835000 12.315000 2.105000 ;
      RECT 11.985000  2.105000 12.285000 2.635000 ;
      RECT 12.020000  0.085000 12.235000 0.545000 ;
      RECT 12.405000  0.255000 12.735000 0.715000 ;
      RECT 12.455000  2.210000 12.785000 2.465000 ;
      RECT 12.485000  1.665000 12.785000 2.210000 ;
      RECT 12.975000  1.495000 14.165000 1.665000 ;
      RECT 12.975000  1.665000 13.275000 2.210000 ;
      RECT 12.975000  2.210000 13.305000 2.465000 ;
      RECT 13.025000  0.255000 13.355000 0.715000 ;
      RECT 13.025000  0.715000 14.215000 0.885000 ;
      RECT 13.445000  1.835000 13.775000 2.105000 ;
      RECT 13.475000  2.105000 13.775000 2.635000 ;
      RECT 13.525000  0.085000 13.740000 0.545000 ;
      RECT 13.910000  0.255000 15.055000 0.425000 ;
      RECT 13.910000  0.425000 14.215000 0.715000 ;
      RECT 13.910000  0.885000 14.215000 0.925000 ;
      RECT 13.995000  1.665000 14.165000 2.295000 ;
      RECT 13.995000  2.295000 15.160000 2.465000 ;
      RECT 14.345000  1.755000 14.775000 2.125000 ;
      RECT 14.385000  0.595000 14.715000 0.885000 ;
      RECT 14.465000  0.885000 14.635000 1.755000 ;
      RECT 14.885000  0.425000 15.055000 0.770000 ;
      RECT 14.980000  1.205000 15.395000 1.305000 ;
      RECT 14.980000  1.305000 15.500000 1.465000 ;
      RECT 14.980000  1.465000 15.760000 1.475000 ;
      RECT 14.990000  1.645000 15.160000 2.295000 ;
      RECT 15.225000  0.585000 15.805000 0.755000 ;
      RECT 15.225000  0.755000 15.395000 1.205000 ;
      RECT 15.330000  1.475000 15.760000 1.635000 ;
      RECT 15.430000  1.635000 15.760000 2.465000 ;
      RECT 15.555000  0.330000 15.805000 0.585000 ;
      RECT 15.935000  1.465000 16.265000 2.635000 ;
      RECT 15.975000  0.085000 16.225000 0.660000 ;
      RECT 16.395000  0.330000 16.645000 0.585000 ;
      RECT 16.395000  0.585000 16.975000 0.755000 ;
      RECT 16.440000  1.465000 17.220000 1.475000 ;
      RECT 16.440000  1.475000 16.870000 1.635000 ;
      RECT 16.440000  1.635000 16.770000 2.465000 ;
      RECT 16.700000  1.305000 17.220000 1.465000 ;
      RECT 16.805000  0.755000 16.975000 1.205000 ;
      RECT 16.805000  1.205000 17.220000 1.305000 ;
      RECT 17.040000  1.645000 17.210000 2.295000 ;
      RECT 17.040000  2.295000 18.205000 2.465000 ;
      RECT 17.145000  0.255000 18.290000 0.425000 ;
      RECT 17.145000  0.425000 17.315000 0.770000 ;
      RECT 17.425000  1.755000 17.855000 2.125000 ;
      RECT 17.485000  0.595000 17.815000 0.885000 ;
      RECT 17.565000  0.885000 17.735000 1.755000 ;
      RECT 17.985000  0.425000 18.290000 0.715000 ;
      RECT 17.985000  0.715000 19.175000 0.885000 ;
      RECT 17.985000  0.885000 18.290000 0.925000 ;
      RECT 18.035000  1.495000 19.225000 1.665000 ;
      RECT 18.035000  1.665000 18.205000 2.295000 ;
      RECT 18.425000  1.835000 18.755000 2.105000 ;
      RECT 18.425000  2.105000 18.725000 2.635000 ;
      RECT 18.460000  0.085000 18.675000 0.545000 ;
      RECT 18.845000  0.255000 19.175000 0.715000 ;
      RECT 18.895000  2.210000 19.225000 2.465000 ;
      RECT 18.925000  1.665000 19.225000 2.210000 ;
      RECT 19.415000  1.495000 20.605000 1.665000 ;
      RECT 19.415000  1.665000 19.715000 2.210000 ;
      RECT 19.415000  2.210000 19.745000 2.465000 ;
      RECT 19.465000  0.255000 19.795000 0.715000 ;
      RECT 19.465000  0.715000 20.655000 0.885000 ;
      RECT 19.885000  1.835000 20.215000 2.105000 ;
      RECT 19.915000  2.105000 20.215000 2.635000 ;
      RECT 19.965000  0.085000 20.180000 0.545000 ;
      RECT 20.350000  0.255000 21.495000 0.425000 ;
      RECT 20.350000  0.425000 20.655000 0.715000 ;
      RECT 20.350000  0.885000 20.655000 0.925000 ;
      RECT 20.435000  1.665000 20.605000 2.295000 ;
      RECT 20.435000  2.295000 21.600000 2.465000 ;
      RECT 20.785000  1.755000 21.215000 2.125000 ;
      RECT 20.825000  0.595000 21.155000 0.885000 ;
      RECT 20.905000  0.885000 21.075000 1.755000 ;
      RECT 21.325000  0.425000 21.495000 0.770000 ;
      RECT 21.420000  1.205000 21.835000 1.305000 ;
      RECT 21.420000  1.305000 21.940000 1.465000 ;
      RECT 21.420000  1.465000 22.200000 1.475000 ;
      RECT 21.430000  1.645000 21.600000 2.295000 ;
      RECT 21.665000  0.585000 22.245000 0.755000 ;
      RECT 21.665000  0.755000 21.835000 1.205000 ;
      RECT 21.770000  1.475000 22.200000 1.635000 ;
      RECT 21.870000  1.635000 22.200000 2.465000 ;
      RECT 21.995000  0.330000 22.245000 0.585000 ;
      RECT 22.375000  1.465000 22.705000 2.635000 ;
      RECT 22.415000  0.085000 22.665000 0.660000 ;
      RECT 22.835000  0.330000 23.085000 0.585000 ;
      RECT 22.835000  0.585000 23.415000 0.755000 ;
      RECT 22.880000  1.465000 23.660000 1.475000 ;
      RECT 22.880000  1.475000 23.310000 1.635000 ;
      RECT 22.880000  1.635000 23.210000 2.465000 ;
      RECT 23.140000  1.305000 23.660000 1.465000 ;
      RECT 23.245000  0.755000 23.415000 1.205000 ;
      RECT 23.245000  1.205000 23.660000 1.305000 ;
      RECT 23.480000  1.645000 23.650000 2.295000 ;
      RECT 23.480000  2.295000 24.645000 2.465000 ;
      RECT 23.585000  0.255000 24.730000 0.425000 ;
      RECT 23.585000  0.425000 23.755000 0.770000 ;
      RECT 23.865000  1.755000 24.295000 2.125000 ;
      RECT 23.925000  0.595000 24.255000 0.885000 ;
      RECT 24.005000  0.885000 24.175000 1.755000 ;
      RECT 24.425000  0.425000 24.730000 0.715000 ;
      RECT 24.425000  0.715000 25.615000 0.885000 ;
      RECT 24.425000  0.885000 24.730000 0.925000 ;
      RECT 24.475000  1.495000 25.665000 1.665000 ;
      RECT 24.475000  1.665000 24.645000 2.295000 ;
      RECT 24.865000  1.835000 25.195000 2.105000 ;
      RECT 24.865000  2.105000 25.165000 2.635000 ;
      RECT 24.900000  0.085000 25.115000 0.545000 ;
      RECT 25.285000  0.255000 25.615000 0.715000 ;
      RECT 25.335000  2.210000 25.665000 2.465000 ;
      RECT 25.365000  1.665000 25.665000 2.210000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.785000  1.695000 1.955000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.785000  4.915000 1.955000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  1.785000  8.135000 1.955000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  1.785000 11.355000 1.955000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  1.785000 14.575000 1.955000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
      RECT 17.165000 -0.085000 17.335000 0.085000 ;
      RECT 17.165000  2.635000 17.335000 2.805000 ;
      RECT 17.625000 -0.085000 17.795000 0.085000 ;
      RECT 17.625000  1.785000 17.795000 1.955000 ;
      RECT 17.625000  2.635000 17.795000 2.805000 ;
      RECT 18.085000 -0.085000 18.255000 0.085000 ;
      RECT 18.085000  2.635000 18.255000 2.805000 ;
      RECT 18.545000 -0.085000 18.715000 0.085000 ;
      RECT 18.545000  2.635000 18.715000 2.805000 ;
      RECT 19.005000 -0.085000 19.175000 0.085000 ;
      RECT 19.005000  2.635000 19.175000 2.805000 ;
      RECT 19.465000 -0.085000 19.635000 0.085000 ;
      RECT 19.465000  2.635000 19.635000 2.805000 ;
      RECT 19.925000 -0.085000 20.095000 0.085000 ;
      RECT 19.925000  2.635000 20.095000 2.805000 ;
      RECT 20.385000 -0.085000 20.555000 0.085000 ;
      RECT 20.385000  2.635000 20.555000 2.805000 ;
      RECT 20.845000 -0.085000 21.015000 0.085000 ;
      RECT 20.845000  1.785000 21.015000 1.955000 ;
      RECT 20.845000  2.635000 21.015000 2.805000 ;
      RECT 21.305000 -0.085000 21.475000 0.085000 ;
      RECT 21.305000  2.635000 21.475000 2.805000 ;
      RECT 21.765000 -0.085000 21.935000 0.085000 ;
      RECT 21.765000  2.635000 21.935000 2.805000 ;
      RECT 22.225000 -0.085000 22.395000 0.085000 ;
      RECT 22.225000 -0.085000 22.395000 0.085000 ;
      RECT 22.225000  2.635000 22.395000 2.805000 ;
      RECT 22.225000  2.635000 22.395000 2.805000 ;
      RECT 22.685000 -0.085000 22.855000 0.085000 ;
      RECT 22.685000 -0.085000 22.855000 0.085000 ;
      RECT 22.685000  2.635000 22.855000 2.805000 ;
      RECT 22.685000  2.635000 22.855000 2.805000 ;
      RECT 23.145000 -0.085000 23.315000 0.085000 ;
      RECT 23.145000  2.635000 23.315000 2.805000 ;
      RECT 23.605000 -0.085000 23.775000 0.085000 ;
      RECT 23.605000  2.635000 23.775000 2.805000 ;
      RECT 24.065000 -0.085000 24.235000 0.085000 ;
      RECT 24.065000  1.785000 24.235000 1.955000 ;
      RECT 24.065000  2.635000 24.235000 2.805000 ;
      RECT 24.525000 -0.085000 24.695000 0.085000 ;
      RECT 24.525000  2.635000 24.695000 2.805000 ;
      RECT 24.985000 -0.085000 25.155000 0.085000 ;
      RECT 24.985000  2.635000 25.155000 2.805000 ;
      RECT 25.445000 -0.085000 25.615000 0.085000 ;
      RECT 25.445000  2.635000 25.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb8to1_2


MACRO sky130_fd_sc_hdll__a32o_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875000 0.415000 3.145000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 0.425000 3.650000 1.625000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 0.995000 4.505000 1.630000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.235000 1.075000 2.670000 1.245000 ;
        RECT 2.445000 1.245000 2.670000 1.615000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.745000 1.630000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.748000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.655000 0.895000 0.825000 ;
        RECT 0.135000 0.825000 0.345000 1.785000 ;
        RECT 0.135000 1.785000 1.285000 1.955000 ;
        RECT 0.135000 1.955000 0.345000 2.465000 ;
        RECT 1.115000 1.955000 1.285000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.465000 ;
      RECT 0.515000  2.125000 0.895000 2.635000 ;
      RECT 0.535000  0.995000 0.755000 1.445000 ;
      RECT 0.535000  1.445000 2.275000 1.615000 ;
      RECT 0.985000  0.085000 1.740000 0.445000 ;
      RECT 1.635000  1.785000 1.805000 2.295000 ;
      RECT 1.635000  2.295000 2.745000 2.465000 ;
      RECT 1.800000  0.675000 2.705000 0.845000 ;
      RECT 1.800000  0.845000 2.040000 1.445000 ;
      RECT 2.025000  1.615000 2.275000 1.945000 ;
      RECT 2.025000  1.945000 2.355000 2.115000 ;
      RECT 2.405000  0.295000 2.705000 0.675000 ;
      RECT 2.575000  1.795000 3.845000 1.965000 ;
      RECT 2.575000  1.965000 2.745000 2.295000 ;
      RECT 2.915000  2.140000 3.295000 2.635000 ;
      RECT 3.675000  1.965000 3.845000 2.465000 ;
      RECT 4.015000  0.085000 4.400000 0.805000 ;
      RECT 4.015000  1.915000 4.400000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32o_2


MACRO sky130_fd_sc_hdll__a32o_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.260000 0.955000 2.665000 1.325000 ;
        RECT 2.380000 0.665000 2.665000 0.955000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.665000 1.950000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 0.995000 1.355000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.835000 0.660000 3.135000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.430000 0.995000 4.030000 1.325000 ;
        RECT 3.790000 1.325000 4.030000 1.615000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.554500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.300000 0.425000 0.560000 ;
        RECT 0.090000 0.560000 0.345000 1.915000 ;
        RECT 0.090000 1.915000 0.425000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.570000  0.995000 0.845000 1.325000 ;
      RECT 0.595000  0.085000 0.975000 0.485000 ;
      RECT 0.675000  0.655000 1.315000 0.825000 ;
      RECT 0.675000  0.825000 0.845000 0.995000 ;
      RECT 0.675000  1.325000 0.845000 1.495000 ;
      RECT 0.675000  1.495000 3.325000 1.665000 ;
      RECT 0.725000  1.835000 1.055000 2.635000 ;
      RECT 1.145000  0.315000 2.910000 0.485000 ;
      RECT 1.145000  0.485000 1.315000 0.655000 ;
      RECT 1.350000  1.875000 2.875000 2.045000 ;
      RECT 1.350000  2.045000 1.635000 2.465000 ;
      RECT 1.940000  2.215000 2.270000 2.635000 ;
      RECT 2.545000  2.045000 2.875000 2.295000 ;
      RECT 2.545000  2.295000 3.895000 2.465000 ;
      RECT 3.155000  1.665000 3.325000 2.125000 ;
      RECT 3.505000  0.085000 3.885000 0.805000 ;
      RECT 3.635000  1.795000 3.895000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32o_1


MACRO sky130_fd_sc_hdll__a32o_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.280000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.680000 1.075000 5.575000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.635000 1.075000 4.430000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.410000 1.075000 3.405000 1.295000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.120000 1.075000 7.140000 1.625000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.440000 1.075000 8.170000 1.295000 ;
        RECT 7.440000 1.295000 7.635000 1.635000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.635000 1.755000 0.805000 ;
        RECT 0.120000 0.805000 0.340000 1.495000 ;
        RECT 0.120000 1.495000 1.755000 1.665000 ;
        RECT 0.645000 0.255000 0.815000 0.635000 ;
        RECT 0.645000 1.665000 0.815000 2.465000 ;
        RECT 1.585000 0.255000 1.755000 0.635000 ;
        RECT 1.585000 1.665000 1.755000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.095000  1.915000 0.425000 2.635000 ;
      RECT 0.620000  0.995000 2.170000 1.325000 ;
      RECT 0.985000  0.085000 1.365000 0.465000 ;
      RECT 0.985000  1.915000 1.365000 2.635000 ;
      RECT 1.925000  0.085000 2.305000 0.465000 ;
      RECT 1.925000  1.915000 2.305000 2.635000 ;
      RECT 1.950000  1.325000 2.170000 1.495000 ;
      RECT 1.950000  1.495000 5.950000 1.665000 ;
      RECT 2.525000  0.255000 2.695000 0.655000 ;
      RECT 2.525000  0.655000 4.235000 0.825000 ;
      RECT 2.525000  1.915000 5.565000 2.085000 ;
      RECT 2.525000  2.085000 2.695000 2.465000 ;
      RECT 2.865000  0.085000 3.245000 0.465000 ;
      RECT 2.865000  2.255000 3.245000 2.635000 ;
      RECT 3.435000  0.295000 5.645000 0.465000 ;
      RECT 3.515000  2.085000 3.685000 2.465000 ;
      RECT 3.855000  2.255000 4.235000 2.635000 ;
      RECT 4.455000  2.085000 4.625000 2.465000 ;
      RECT 4.795000  0.635000 6.735000 0.805000 ;
      RECT 4.795000  2.255000 5.175000 2.635000 ;
      RECT 5.395000  2.085000 5.565000 2.255000 ;
      RECT 5.395000  2.255000 8.185000 2.425000 ;
      RECT 5.780000  0.805000 5.950000 1.495000 ;
      RECT 5.780000  1.665000 5.950000 1.905000 ;
      RECT 5.780000  1.905000 6.510000 1.915000 ;
      RECT 5.780000  1.915000 7.715000 2.075000 ;
      RECT 5.930000  0.295000 7.165000 0.465000 ;
      RECT 6.445000  2.075000 7.715000 2.085000 ;
      RECT 6.995000  0.255000 7.165000 0.295000 ;
      RECT 6.995000  0.465000 7.165000 0.645000 ;
      RECT 6.995000  0.645000 8.105000 0.815000 ;
      RECT 7.335000  0.085000 7.715000 0.465000 ;
      RECT 7.935000  0.255000 8.105000 0.645000 ;
      RECT 7.935000  1.755000 8.185000 2.255000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32o_4


MACRO sky130_fd_sc_hdll__o32ai_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.395000 0.995000 2.990000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.915000 0.995000 2.205000 2.465000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 0.995000 1.745000 1.615000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.685000 0.360000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.920000 0.995000 1.305000 1.615000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.758800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 0.655000 0.895000 0.825000 ;
        RECT 0.530000 0.825000 0.750000 1.785000 ;
        RECT 0.530000 1.785000 1.530000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.255000 1.440000 0.485000 ;
      RECT 0.090000  1.495000 0.360000 2.635000 ;
      RECT 1.065000  0.485000 1.440000 0.655000 ;
      RECT 1.065000  0.655000 2.555000 0.825000 ;
      RECT 1.645000  0.085000 1.975000 0.485000 ;
      RECT 2.385000  0.375000 2.555000 0.655000 ;
      RECT 2.725000  0.085000 3.095000 0.825000 ;
      RECT 2.785000  1.495000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o32ai_1


MACRO sky130_fd_sc_hdll__o32ai_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.04000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.090000 1.075000 10.925000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.520000 1.075000 8.010000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.170000 1.075000 5.980000 1.275000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.075000 3.940000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.835000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.655000 3.730000 0.905000 ;
        RECT 0.515000 1.495000 6.130000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.085000 ;
        RECT 1.455000 1.665000 1.850000 2.085000 ;
        RECT 2.055000 0.905000 2.235000 1.495000 ;
        RECT 4.860000 1.665000 5.190000 2.085000 ;
        RECT 5.750000 1.665000 6.130000 2.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.090000  0.255000  4.200000 0.465000 ;
      RECT  0.090000  0.465000  0.345000 0.905000 ;
      RECT  0.090000  1.495000  0.345000 2.255000 ;
      RECT  0.090000  2.255000  2.240000 2.465000 ;
      RECT  1.115000  1.835000  1.285000 2.255000 ;
      RECT  2.070000  1.835000  4.200000 2.005000 ;
      RECT  2.070000  2.005000  2.240000 2.255000 ;
      RECT  2.410000  2.175000  2.790000 2.635000 ;
      RECT  3.010000  2.005000  3.180000 2.425000 ;
      RECT  3.350000  2.175000  3.730000 2.635000 ;
      RECT  3.950000  0.465000  4.200000 0.735000 ;
      RECT  3.950000  0.735000 10.925000 0.905000 ;
      RECT  3.950000  2.005000  4.200000 2.465000 ;
      RECT  4.390000  1.835000  4.640000 2.255000 ;
      RECT  4.390000  2.255000  8.480000 2.465000 ;
      RECT  4.420000  0.085000  4.590000 0.545000 ;
      RECT  4.760000  0.255000  5.140000 0.735000 ;
      RECT  5.360000  0.085000  5.690000 0.545000 ;
      RECT  5.410000  1.835000  5.580000 2.255000 ;
      RECT  5.910000  0.255000  6.580000 0.735000 ;
      RECT  6.350000  1.835000  6.520000 2.255000 ;
      RECT  6.690000  1.495000 10.410000 1.665000 ;
      RECT  6.690000  1.665000  7.070000 2.085000 ;
      RECT  6.820000  0.085000  6.990000 0.545000 ;
      RECT  7.160000  0.255000  7.540000 0.735000 ;
      RECT  7.290000  1.835000  7.460000 2.255000 ;
      RECT  7.630000  1.665000  8.010000 2.085000 ;
      RECT  7.760000  0.085000  7.930000 0.545000 ;
      RECT  8.100000  0.255000  8.840000 0.735000 ;
      RECT  8.230000  1.835000  8.480000 2.255000 ;
      RECT  8.670000  1.835000  8.920000 2.635000 ;
      RECT  9.090000  1.665000  9.470000 2.465000 ;
      RECT  9.220000  0.085000  9.390000 0.545000 ;
      RECT  9.560000  0.255000  9.940000 0.735000 ;
      RECT  9.690000  1.835000  9.860000 2.635000 ;
      RECT 10.030000  1.665000 10.410000 2.465000 ;
      RECT 10.160000  0.085000 10.375000 0.545000 ;
      RECT 10.545000  0.255000 10.925000 0.735000 ;
      RECT 10.675000  1.495000 10.925000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o32ai_4


MACRO sky130_fd_sc_hdll__o32ai_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.200000 1.075000 6.295000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.720000 1.075000 4.930000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.655000 1.075000 3.365000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.815000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.895000 1.325000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.061000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.655000 2.245000 0.905000 ;
        RECT 0.515000 1.495000 3.405000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.095000 ;
        RECT 1.985000 0.905000 2.245000 1.105000 ;
        RECT 1.985000 1.105000 2.370000 1.495000 ;
        RECT 3.025000 1.665000 3.405000 2.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.090000  0.255000 2.655000 0.485000 ;
      RECT 0.090000  0.485000 0.345000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.295000 ;
      RECT 0.090000  2.295000 1.365000 2.465000 ;
      RECT 1.115000  1.835000 2.305000 2.005000 ;
      RECT 1.115000  2.005000 1.365000 2.295000 ;
      RECT 1.585000  2.175000 1.755000 2.635000 ;
      RECT 1.925000  2.005000 2.305000 2.455000 ;
      RECT 2.485000  0.485000 2.655000 0.715000 ;
      RECT 2.485000  0.715000 6.305000 0.905000 ;
      RECT 2.585000  1.835000 2.835000 2.255000 ;
      RECT 2.585000  2.255000 4.835000 2.445000 ;
      RECT 2.870000  0.085000 3.250000 0.545000 ;
      RECT 3.435000  0.255000 3.815000 0.715000 ;
      RECT 3.625000  1.495000 3.795000 2.255000 ;
      RECT 4.015000  1.495000 5.825000 1.665000 ;
      RECT 4.015000  1.665000 4.345000 2.085000 ;
      RECT 4.035000  0.085000 4.205000 0.545000 ;
      RECT 4.505000  0.255000 5.175000 0.715000 ;
      RECT 4.585000  1.835000 4.835000 2.255000 ;
      RECT 5.070000  1.835000 5.275000 2.635000 ;
      RECT 5.355000  0.085000 5.735000 0.545000 ;
      RECT 5.495000  1.665000 5.825000 2.460000 ;
      RECT 5.975000  0.255000 6.305000 0.715000 ;
      RECT 6.045000  1.495000 6.265000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o32ai_2


MACRO sky130_fd_sc_hdll__clkinv_12
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.200000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  3.996000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.035000 7.925000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.290400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.695000 8.655000 0.865000 ;
        RECT 0.115000 0.865000 0.285000 1.460000 ;
        RECT 0.115000 1.460000 8.655000 1.630000 ;
        RECT 0.595000 1.630000 0.865000 2.465000 ;
        RECT 1.535000 1.630000 1.805000 2.465000 ;
        RECT 2.005000 0.255000 2.275000 0.695000 ;
        RECT 2.475000 1.630000 2.745000 2.465000 ;
        RECT 2.945000 0.255000 3.215000 0.695000 ;
        RECT 3.415000 1.630000 3.685000 2.465000 ;
        RECT 3.885000 0.255000 4.155000 0.695000 ;
        RECT 4.355000 1.630000 4.625000 2.465000 ;
        RECT 4.825000 0.255000 5.095000 0.695000 ;
        RECT 5.295000 1.630000 5.565000 2.465000 ;
        RECT 5.765000 0.255000 6.035000 0.695000 ;
        RECT 6.235000 1.630000 6.505000 2.465000 ;
        RECT 6.705000 0.255000 6.975000 0.695000 ;
        RECT 7.175000 1.630000 7.445000 2.465000 ;
        RECT 8.100000 0.865000 8.655000 1.460000 ;
        RECT 8.115000 1.630000 8.385000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.095000  1.800000 0.425000 2.635000 ;
      RECT 1.035000  1.800000 1.365000 2.635000 ;
      RECT 1.165000  0.085000 1.835000 0.525000 ;
      RECT 1.975000  1.800000 2.305000 2.635000 ;
      RECT 2.445000  0.085000 2.775000 0.525000 ;
      RECT 2.915000  1.800000 3.245000 2.635000 ;
      RECT 3.385000  0.085000 3.715000 0.525000 ;
      RECT 3.855000  1.800000 4.185000 2.635000 ;
      RECT 4.325000  0.085000 4.655000 0.525000 ;
      RECT 4.795000  1.800000 5.125000 2.635000 ;
      RECT 5.265000  0.085000 5.595000 0.525000 ;
      RECT 5.735000  1.800000 6.065000 2.635000 ;
      RECT 6.205000  0.085000 6.535000 0.525000 ;
      RECT 6.675000  1.800000 7.005000 2.635000 ;
      RECT 7.145000  0.085000 7.815000 0.525000 ;
      RECT 7.615000  1.800000 7.945000 2.635000 ;
      RECT 8.555000  1.800000 8.885000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_12


MACRO sky130_fd_sc_hdll__clkinv_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.332000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.065000 2.910000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.177200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.725000 3.570000 0.895000 ;
        RECT 0.105000 0.895000 0.275000 1.460000 ;
        RECT 0.105000 1.460000 3.570000 1.630000 ;
        RECT 0.655000 1.630000 0.910000 2.435000 ;
        RECT 1.130000 0.280000 1.390000 0.725000 ;
        RECT 1.615000 1.630000 1.870000 2.435000 ;
        RECT 2.090000 0.280000 2.345000 0.725000 ;
        RECT 2.570000 1.630000 2.830000 2.435000 ;
        RECT 3.270000 0.895000 3.570000 1.460000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  1.800000 0.430000 2.635000 ;
      RECT 0.565000  0.085000 0.910000 0.555000 ;
      RECT 1.130000  1.800000 1.390000 2.635000 ;
      RECT 1.610000  0.085000 1.870000 0.555000 ;
      RECT 2.090000  1.800000 2.350000 2.635000 ;
      RECT 2.565000  0.085000 2.865000 0.555000 ;
      RECT 3.050000  1.800000 3.435000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_4


MACRO sky130_fd_sc_hdll__clkinv_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.666000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.065000 1.335000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.728600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.460000 2.155000 1.630000 ;
        RECT 0.155000 1.630000 0.410000 2.435000 ;
        RECT 1.110000 1.630000 1.370000 2.435000 ;
        RECT 1.125000 0.280000 1.350000 0.725000 ;
        RECT 1.125000 0.725000 2.155000 0.895000 ;
        RECT 1.520000 0.895000 2.155000 1.460000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.560000  0.085000 0.905000 0.610000 ;
      RECT 0.630000  1.800000 0.890000 2.635000 ;
      RECT 1.520000  0.085000 1.900000 0.555000 ;
      RECT 1.605000  1.800000 1.860000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_2


MACRO sky130_fd_sc_hdll__clkinv_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  1.840000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.365400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.375000 0.325000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.375900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.890000 0.760000 ;
        RECT 0.515000 0.760000 1.395000 1.290000 ;
        RECT 0.515000 1.290000 0.895000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  1.665000 0.345000 2.635000 ;
      RECT 1.115000  0.085000 1.395000 0.590000 ;
      RECT 1.115000  1.665000 1.395000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_1


MACRO sky130_fd_sc_hdll__clkinv_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.664000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.035000 5.565000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.386400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.695000 6.330000 0.865000 ;
        RECT 0.115000 0.865000 0.285000 1.460000 ;
        RECT 0.115000 1.460000 6.330000 1.630000 ;
        RECT 0.615000 1.630000 0.855000 2.435000 ;
        RECT 1.555000 1.630000 1.795000 2.435000 ;
        RECT 1.685000 0.280000 1.875000 0.695000 ;
        RECT 2.495000 1.630000 2.745000 2.435000 ;
        RECT 2.645000 0.280000 2.835000 0.695000 ;
        RECT 3.430000 1.630000 3.675000 2.435000 ;
        RECT 3.605000 0.280000 3.795000 0.695000 ;
        RECT 4.420000 1.630000 4.725000 2.435000 ;
        RECT 4.665000 0.280000 4.855000 0.695000 ;
        RECT 5.465000 1.630000 5.705000 2.435000 ;
        RECT 6.060000 0.865000 6.330000 1.460000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.135000  1.800000 0.395000 2.635000 ;
      RECT 1.075000  1.800000 1.335000 2.635000 ;
      RECT 1.135000  0.085000 1.465000 0.525000 ;
      RECT 2.015000  1.800000 2.275000 2.635000 ;
      RECT 2.095000  0.085000 2.425000 0.525000 ;
      RECT 2.965000  1.800000 3.210000 2.635000 ;
      RECT 3.055000  0.085000 3.435000 0.525000 ;
      RECT 3.895000  1.800000 4.200000 2.635000 ;
      RECT 4.015000  0.085000 4.445000 0.525000 ;
      RECT 4.945000  1.800000 5.245000 2.635000 ;
      RECT 5.075000  0.085000 5.505000 0.525000 ;
      RECT 5.925000  1.800000 6.180000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_8


MACRO sky130_fd_sc_hdll__clkinv_16
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  12.42000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  5.328000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.345000 0.895000 2.355000 1.275000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.928900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.625000 1.455000 11.630000 1.665000 ;
        RECT  0.625000 1.665000  0.880000 2.465000 ;
        RECT  1.585000 1.665000  1.840000 2.450000 ;
        RECT  2.575000 0.280000  2.800000 1.415000 ;
        RECT  2.575000 1.415000  9.705000 1.455000 ;
        RECT  2.575000 1.665000  2.800000 2.465000 ;
        RECT  3.505000 0.280000  3.760000 1.415000 ;
        RECT  3.505000 1.665000  3.760000 2.450000 ;
        RECT  4.465000 0.280000  4.705000 1.415000 ;
        RECT  4.465000 1.665000  4.705000 2.450000 ;
        RECT  5.455000 0.280000  5.805000 1.415000 ;
        RECT  5.455000 1.665000  5.830000 2.450000 ;
        RECT  6.575000 0.280000  6.825000 1.415000 ;
        RECT  6.575000 1.665000  6.825000 2.450000 ;
        RECT  7.535000 0.280000  7.785000 1.415000 ;
        RECT  7.535000 1.665000  7.785000 2.450000 ;
        RECT  8.495000 0.280000  8.745000 1.415000 ;
        RECT  8.495000 1.665000  8.745000 2.450000 ;
        RECT  9.455000 0.280000  9.705000 1.415000 ;
        RECT  9.455000 1.665000  9.705000 2.450000 ;
        RECT 10.415000 1.665000 10.655000 2.450000 ;
        RECT 11.375000 1.665000 11.630000 2.450000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.140000  1.495000  0.405000 2.635000 ;
      RECT  1.100000  1.835000  1.360000 2.635000 ;
      RECT  2.055000  0.085000  2.325000 0.610000 ;
      RECT  2.065000  1.835000  2.320000 2.635000 ;
      RECT  3.020000  0.085000  3.285000 0.610000 ;
      RECT  3.020000  1.835000  3.280000 2.635000 ;
      RECT  3.980000  0.085000  4.245000 0.610000 ;
      RECT  3.985000  1.835000  4.240000 2.635000 ;
      RECT  4.965000  0.085000  5.230000 0.610000 ;
      RECT  4.965000  1.835000  5.220000 2.635000 ;
      RECT  6.090000  0.085000  6.355000 0.610000 ;
      RECT  6.090000  1.835000  6.345000 2.120000 ;
      RECT  6.090000  2.120000  6.350000 2.635000 ;
      RECT  7.050000  0.085000  7.275000 0.610000 ;
      RECT  7.055000  1.835000  7.310000 2.635000 ;
      RECT  8.010000  0.085000  8.275000 0.610000 ;
      RECT  8.015000  1.835000  8.270000 2.635000 ;
      RECT  8.970000  0.085000  9.235000 0.610000 ;
      RECT  8.975000  1.835000  9.230000 2.635000 ;
      RECT  9.930000  0.085000 10.195000 0.610000 ;
      RECT  9.930000  0.895000 11.910000 1.275000 ;
      RECT  9.935000  1.835000 10.190000 2.635000 ;
      RECT 10.895000  1.835000 11.150000 2.635000 ;
      RECT 11.850000  1.835000 12.110000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.675000  1.105000  1.845000 1.275000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.185000  1.105000  2.355000 1.275000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.395000  1.105000 10.565000 1.275000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.905000  1.105000 11.075000 1.275000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
    LAYER met1 ;
      RECT  1.615000 1.075000  2.415000 1.120000 ;
      RECT  1.615000 1.120000 11.135000 1.260000 ;
      RECT  1.615000 1.260000  2.415000 1.305000 ;
      RECT 10.285000 1.075000 11.135000 1.120000 ;
      RECT 10.285000 1.260000 11.135000 1.305000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_16


MACRO sky130_fd_sc_hdll__and3_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.470000 1.245000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 2.125000 1.520000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.305000 1.315000 0.750000 ;
        RECT 1.065000 0.750000 1.625000 1.245000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.255000 2.430000 0.715000 ;
        RECT 2.170000 1.795000 2.620000 2.465000 ;
        RECT 2.260000 0.715000 2.430000 0.925000 ;
        RECT 2.260000 0.925000 2.925000 1.445000 ;
        RECT 2.260000 1.445000 2.620000 1.795000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  2.130000 0.765000 2.635000 ;
      RECT 0.100000  1.425000 2.040000 1.595000 ;
      RECT 0.100000  1.595000 0.355000 1.960000 ;
      RECT 0.105000  0.305000 0.895000 0.570000 ;
      RECT 0.525000  1.765000 0.905000 1.955000 ;
      RECT 0.525000  1.955000 0.765000 2.130000 ;
      RECT 0.690000  0.570000 0.895000 1.425000 ;
      RECT 1.180000  1.595000 1.480000 1.890000 ;
      RECT 1.485000  0.085000 1.815000 0.580000 ;
      RECT 1.705000  1.790000 1.920000 2.635000 ;
      RECT 1.810000  0.995000 2.040000 1.425000 ;
      RECT 2.695000  0.085000 2.970000 0.745000 ;
      RECT 2.790000  1.625000 3.050000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3_2


MACRO sky130_fd_sc_hdll__and3_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.995000 0.875000 1.340000 ;
        RECT 0.115000 1.340000 0.330000 2.335000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 0.745000 1.355000 1.340000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 2.050000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.061500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.650000 0.515000 2.840000 0.615000 ;
        RECT 2.650000 0.615000 4.490000 0.845000 ;
        RECT 2.650000 1.535000 4.490000 1.760000 ;
        RECT 2.650000 1.760000 2.840000 2.465000 ;
        RECT 3.610000 0.255000 3.800000 0.615000 ;
        RECT 3.610000 1.760000 4.490000 1.765000 ;
        RECT 3.610000 1.765000 3.800000 2.465000 ;
        RECT 4.210000 0.845000 4.490000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.465000  0.255000 1.825000 0.445000 ;
      RECT 0.465000  0.445000 0.800000 0.805000 ;
      RECT 0.500000  1.580000 2.430000 1.750000 ;
      RECT 0.500000  1.750000 0.680000 2.465000 ;
      RECT 0.895000  1.935000 1.395000 2.635000 ;
      RECT 1.620000  1.750000 1.800000 2.465000 ;
      RECT 1.635000  0.445000 1.825000 0.615000 ;
      RECT 1.635000  0.615000 2.430000 0.805000 ;
      RECT 2.055000  0.085000 2.385000 0.445000 ;
      RECT 2.060000  1.935000 2.390000 2.635000 ;
      RECT 2.220000  0.805000 2.430000 1.020000 ;
      RECT 2.220000  1.020000 3.905000 1.355000 ;
      RECT 2.220000  1.355000 2.430000 1.580000 ;
      RECT 3.010000  0.085000 3.390000 0.445000 ;
      RECT 3.010000  1.935000 3.390000 2.635000 ;
      RECT 3.970000  0.085000 4.350000 0.445000 ;
      RECT 3.970000  1.935000 4.350000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3_4


MACRO sky130_fd_sc_hdll__and3_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.635000 0.685000 1.020000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.915000 2.125000 1.495000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.390000 0.305000 1.760000 1.200000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385000 1.765000 2.660000 2.465000 ;
        RECT 2.400000 0.255000 2.660000 0.735000 ;
        RECT 2.490000 0.735000 2.660000 1.765000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.295000 1.075000 0.465000 ;
      RECT 0.085000  1.190000 1.075000 1.360000 ;
      RECT 0.085000  1.360000 0.345000 1.810000 ;
      RECT 0.085000  1.980000 0.750000 2.080000 ;
      RECT 0.085000  2.080000 0.740000 2.635000 ;
      RECT 0.515000  1.710000 0.895000 1.955000 ;
      RECT 0.515000  1.955000 0.750000 1.980000 ;
      RECT 0.855000  0.465000 1.075000 1.190000 ;
      RECT 0.895000  1.360000 1.075000 1.370000 ;
      RECT 0.895000  1.370000 2.270000 1.540000 ;
      RECT 1.160000  1.540000 2.270000 1.590000 ;
      RECT 1.160000  1.590000 2.165000 1.885000 ;
      RECT 1.910000  2.090000 2.165000 2.635000 ;
      RECT 1.930000  0.085000 2.100000 0.625000 ;
      RECT 2.040000  0.990000 2.270000 1.370000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3_1


MACRO sky130_fd_sc_hdll__a211o_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.290000 1.045000 2.695000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.045000 1.960000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 1.045000 3.195000 1.275000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.045000 3.735000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.504500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.255000 0.835000 2.335000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.085000 0.385000 0.905000 ;
      RECT 0.090000  1.490000 0.385000 2.635000 ;
      RECT 1.005000  0.085000 1.770000 0.445000 ;
      RECT 1.100000  0.695000 3.935000 0.875000 ;
      RECT 1.100000  0.875000 1.355000 1.490000 ;
      RECT 1.100000  1.490000 3.935000 1.660000 ;
      RECT 1.100000  1.830000 1.355000 2.635000 ;
      RECT 1.555000  1.840000 3.045000 2.020000 ;
      RECT 1.555000  2.020000 1.935000 2.465000 ;
      RECT 2.155000  2.190000 2.430000 2.635000 ;
      RECT 2.475000  0.275000 2.855000 0.695000 ;
      RECT 2.715000  2.020000 3.045000 2.465000 ;
      RECT 3.110000  0.085000 3.385000 0.525000 ;
      RECT 3.555000  0.275000 3.935000 0.695000 ;
      RECT 3.555000  1.660000 3.935000 2.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211o_2


MACRO sky130_fd_sc_hdll__a211o_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.865000 0.995000 2.390000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 0.995000 1.695000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.590000 0.995000 3.075000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.305000 0.995000 3.585000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.447300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.265000 0.425000 1.685000 ;
        RECT 0.090000 1.685000 0.355000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.525000  1.915000 0.905000 2.635000 ;
      RECT 0.605000  0.625000 3.535000 0.815000 ;
      RECT 0.605000  0.815000 0.845000 1.505000 ;
      RECT 0.605000  1.505000 3.545000 1.685000 ;
      RECT 0.655000  0.085000 1.400000 0.455000 ;
      RECT 1.095000  1.865000 2.565000 2.095000 ;
      RECT 1.095000  2.095000 1.355000 2.455000 ;
      RECT 1.525000  2.265000 2.085000 2.635000 ;
      RECT 2.195000  0.265000 2.520000 0.625000 ;
      RECT 2.305000  2.095000 2.565000 2.455000 ;
      RECT 2.700000  0.085000 3.080000 0.455000 ;
      RECT 3.205000  1.685000 3.545000 2.455000 ;
      RECT 3.310000  0.265000 3.535000 0.625000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211o_1


MACRO sky130_fd_sc_hdll__a211o_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.360000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.535000 1.020000 5.930000 1.330000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.945000 1.020000 5.325000 1.510000 ;
        RECT 4.945000 1.510000 6.445000 1.700000 ;
        RECT 6.125000 1.020000 6.875000 1.320000 ;
        RECT 6.125000 1.320000 6.445000 1.510000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 0.985000 3.105000 1.325000 ;
        RECT 2.875000 1.325000 3.105000 1.445000 ;
        RECT 2.875000 1.445000 4.625000 1.700000 ;
        RECT 4.245000 0.985000 4.625000 1.445000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.275000 0.985000 4.045000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.071300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.635000 2.225000 0.875000 ;
        RECT 0.085000 0.875000 0.340000 1.495000 ;
        RECT 0.085000 1.495000 1.790000 1.705000 ;
        RECT 0.645000 1.705000 0.830000 2.465000 ;
        RECT 1.085000 0.255000 1.275000 0.615000 ;
        RECT 1.085000 0.615000 2.225000 0.635000 ;
        RECT 1.600000 1.705000 1.790000 2.465000 ;
        RECT 2.045000 0.255000 2.225000 0.615000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.090000  1.875000 0.425000 2.635000 ;
      RECT 0.485000  0.085000 0.865000 0.465000 ;
      RECT 0.525000  1.045000 2.620000 1.325000 ;
      RECT 1.050000  1.875000 1.380000 2.635000 ;
      RECT 1.445000  0.085000 1.825000 0.445000 ;
      RECT 2.010000  1.835000 2.260000 2.635000 ;
      RECT 2.385000  1.325000 2.620000 1.505000 ;
      RECT 2.385000  1.505000 2.705000 1.675000 ;
      RECT 2.395000  0.615000 6.040000 0.805000 ;
      RECT 2.395000  0.805000 2.620000 1.045000 ;
      RECT 2.420000  0.085000 2.805000 0.445000 ;
      RECT 2.530000  1.675000 2.705000 1.870000 ;
      RECT 2.530000  1.870000 3.860000 2.040000 ;
      RECT 2.570000  2.210000 4.900000 2.465000 ;
      RECT 3.025000  0.255000 3.270000 0.615000 ;
      RECT 3.440000  0.085000 3.820000 0.445000 ;
      RECT 4.040000  0.255000 4.420000 0.615000 ;
      RECT 4.570000  1.880000 6.995000 2.105000 ;
      RECT 4.570000  2.105000 4.900000 2.210000 ;
      RECT 4.640000  0.085000 5.010000 0.445000 ;
      RECT 5.070000  2.275000 5.450000 2.635000 ;
      RECT 5.660000  0.275000 6.040000 0.615000 ;
      RECT 5.660000  2.105000 5.970000 2.465000 ;
      RECT 6.140000  2.275000 6.520000 2.635000 ;
      RECT 6.615000  0.085000 6.995000 0.805000 ;
      RECT 6.615000  1.535000 6.995000 1.880000 ;
      RECT 6.740000  2.105000 6.995000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211o_4


MACRO sky130_fd_sc_hdll__dfstp_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.96000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.247200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.870000 1.005000 2.330000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.435000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.725000 0.265000 10.025000 0.715000 ;
        RECT  9.725000 0.715000 11.860000 0.885000 ;
        RECT  9.725000 1.470000 11.860000 1.640000 ;
        RECT  9.725000 1.640000  9.995000 2.465000 ;
        RECT 10.665000 0.265000 10.835000 0.715000 ;
        RECT 10.665000 1.640000 10.835000 2.465000 ;
        RECT 11.605000 0.265000 11.860000 0.715000 ;
        RECT 11.605000 1.640000 11.860000 2.465000 ;
        RECT 11.610000 0.885000 11.860000 1.470000 ;
    END
  END Q
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.220000 0.735000 4.510000 0.780000 ;
        RECT 4.220000 0.780000 7.735000 0.920000 ;
        RECT 4.220000 0.920000 4.510000 0.965000 ;
        RECT 7.445000 0.735000 7.735000 0.780000 ;
        RECT 7.445000 0.920000 7.735000 0.965000 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.960000 0.085000 ;
        RECT  0.515000  0.085000  0.895000 0.465000 ;
        RECT  1.555000  0.085000  1.885000 0.465000 ;
        RECT  3.910000  0.085000  4.370000 0.525000 ;
        RECT  5.140000  0.085000  5.530000 0.545000 ;
        RECT  7.320000  0.085000  8.030000 0.565000 ;
        RECT  9.190000  0.085000  9.475000 0.545000 ;
        RECT 10.195000  0.085000 10.495000 0.545000 ;
        RECT 11.055000  0.085000 11.435000 0.545000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 11.960000 2.805000 ;
        RECT  0.515000 2.135000  0.895000 2.635000 ;
        RECT  1.555000 2.135000  1.885000 2.635000 ;
        RECT  3.730000 2.255000  4.110000 2.635000 ;
        RECT  4.680000 2.255000  5.060000 2.635000 ;
        RECT  6.470000 2.255000  6.940000 2.635000 ;
        RECT  7.710000 1.945000  8.040000 2.635000 ;
        RECT  9.190000 1.835000  9.545000 2.635000 ;
        RECT 10.165000 1.810000 10.420000 2.635000 ;
        RECT 11.055000 1.810000 11.435000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.345000  0.345000 0.635000 ;
      RECT 0.175000 0.635000  0.890000 0.805000 ;
      RECT 0.175000 1.795000  0.890000 1.965000 ;
      RECT 0.175000 1.965000  0.345000 2.465000 ;
      RECT 0.660000 0.805000  0.890000 1.795000 ;
      RECT 1.115000 0.345000  1.340000 2.465000 ;
      RECT 1.530000 0.635000  2.275000 0.825000 ;
      RECT 1.530000 0.825000  1.700000 1.795000 ;
      RECT 1.530000 1.795000  2.275000 1.965000 ;
      RECT 2.105000 0.305000  2.275000 0.635000 ;
      RECT 2.105000 1.965000  2.275000 2.465000 ;
      RECT 2.500000 0.705000  2.770000 1.575000 ;
      RECT 2.500000 1.575000  3.100000 1.955000 ;
      RECT 2.510000 2.250000  3.440000 2.420000 ;
      RECT 2.625000 0.265000  3.740000 0.465000 ;
      RECT 2.950000 0.645000  3.350000 1.015000 ;
      RECT 3.270000 1.230000  3.740000 1.235000 ;
      RECT 3.270000 1.235000  4.770000 1.405000 ;
      RECT 3.270000 1.405000  3.440000 2.250000 ;
      RECT 3.520000 0.465000  3.740000 1.230000 ;
      RECT 3.610000 1.575000  3.910000 1.835000 ;
      RECT 3.610000 1.835000  5.110000 2.085000 ;
      RECT 3.910000 0.735000  4.510000 1.065000 ;
      RECT 4.340000 2.085000  4.510000 2.375000 ;
      RECT 4.470000 1.405000  4.770000 1.565000 ;
      RECT 4.790000 0.295000  4.960000 0.725000 ;
      RECT 4.790000 0.725000  5.110000 1.065000 ;
      RECT 4.940000 1.065000  5.110000 1.835000 ;
      RECT 5.330000 0.725000  6.750000 0.895000 ;
      RECT 5.330000 0.895000  5.500000 1.655000 ;
      RECT 5.330000 1.655000  5.900000 1.965000 ;
      RECT 5.560000 2.165000  6.290000 2.415000 ;
      RECT 5.720000 1.065000  5.900000 1.475000 ;
      RECT 6.070000 1.235000  8.170000 1.405000 ;
      RECT 6.070000 1.405000  6.290000 1.915000 ;
      RECT 6.070000 1.915000  7.380000 2.085000 ;
      RECT 6.070000 2.085000  6.290000 2.165000 ;
      RECT 6.190000 0.305000  7.090000 0.475000 ;
      RECT 6.370000 0.895000  6.750000 1.015000 ;
      RECT 6.460000 1.575000  8.550000 1.745000 ;
      RECT 6.920000 0.475000  7.090000 1.235000 ;
      RECT 7.140000 2.085000  7.380000 2.375000 ;
      RECT 7.260000 0.735000  7.780000 1.005000 ;
      RECT 7.260000 1.005000  7.640000 1.065000 ;
      RECT 7.790000 1.175000  8.170000 1.235000 ;
      RECT 8.210000 0.350000  8.550000 0.680000 ;
      RECT 8.210000 1.745000  8.550000 1.765000 ;
      RECT 8.210000 1.765000  8.380000 2.375000 ;
      RECT 8.340000 0.680000  8.550000 1.575000 ;
      RECT 8.650000 1.915000  8.980000 2.425000 ;
      RECT 8.730000 0.345000  8.980000 1.055000 ;
      RECT 8.730000 1.055000 11.440000 1.275000 ;
      RECT 8.730000 1.275000  8.980000 1.915000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.665000  1.740000  0.835000 1.910000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.165000  0.720000  1.335000 0.890000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.645000  1.740000  2.815000 1.910000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.155000  0.720000  3.325000 0.890000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.280000  0.765000  4.450000 0.935000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.705000  1.740000  5.875000 1.910000 ;
      RECT  5.725000  1.110000  5.895000 1.280000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  0.765000  7.675000 0.935000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.605000 1.710000 0.895000 1.800000 ;
      RECT 0.605000 1.800000 5.935000 1.940000 ;
      RECT 1.105000 0.690000 1.395000 0.780000 ;
      RECT 1.105000 0.780000 3.385000 0.920000 ;
      RECT 2.585000 1.710000 2.875000 1.800000 ;
      RECT 3.095000 0.690000 3.385000 0.780000 ;
      RECT 3.170000 0.920000 3.385000 1.120000 ;
      RECT 3.170000 1.120000 5.955000 1.260000 ;
      RECT 5.645000 1.710000 5.935000 1.800000 ;
      RECT 5.665000 1.080000 5.955000 1.120000 ;
      RECT 5.665000 1.260000 5.955000 1.310000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfstp_4


MACRO sky130_fd_sc_hdll__dfstp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.58000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.247200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.870000 1.005000 2.330000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.540000 1.495000 10.485000 1.615000 ;
        RECT 9.540000 1.615000 10.015000 2.460000 ;
        RECT 9.685000 0.265000 10.015000 0.745000 ;
        RECT 9.685000 0.745000 10.485000 0.825000 ;
        RECT 9.750000 0.825000 10.485000 1.495000 ;
    END
  END Q
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.220000 0.735000 4.510000 0.780000 ;
        RECT 4.220000 0.780000 7.735000 0.920000 ;
        RECT 4.220000 0.920000 4.510000 0.965000 ;
        RECT 7.445000 0.735000 7.735000 0.780000 ;
        RECT 7.445000 0.920000 7.735000 0.965000 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 10.580000 0.085000 ;
        RECT  0.515000  0.085000  0.895000 0.465000 ;
        RECT  1.555000  0.085000  1.885000 0.465000 ;
        RECT  3.910000  0.085000  4.370000 0.525000 ;
        RECT  5.140000  0.085000  5.530000 0.545000 ;
        RECT  7.320000  0.085000  8.030000 0.565000 ;
        RECT  9.070000  0.085000  9.450000 0.825000 ;
        RECT 10.185000  0.085000 10.450000 0.575000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 10.580000 2.805000 ;
        RECT  0.515000 2.135000  0.895000 2.635000 ;
        RECT  1.555000 2.135000  1.885000 2.635000 ;
        RECT  3.730000 2.255000  4.110000 2.635000 ;
        RECT  4.680000 2.255000  5.060000 2.635000 ;
        RECT  6.470000 2.255000  6.940000 2.635000 ;
        RECT  7.710000 1.945000  8.040000 2.635000 ;
        RECT  9.200000 1.495000  9.370000 2.635000 ;
        RECT 10.185000 1.785000 10.450000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.345000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 0.890000 0.805000 ;
      RECT 0.175000 1.795000 0.890000 1.965000 ;
      RECT 0.175000 1.965000 0.345000 2.465000 ;
      RECT 0.660000 0.805000 0.890000 1.795000 ;
      RECT 1.115000 0.345000 1.340000 2.465000 ;
      RECT 1.530000 0.635000 2.275000 0.825000 ;
      RECT 1.530000 0.825000 1.700000 1.795000 ;
      RECT 1.530000 1.795000 2.275000 1.965000 ;
      RECT 2.105000 0.305000 2.275000 0.635000 ;
      RECT 2.105000 1.965000 2.275000 2.465000 ;
      RECT 2.500000 0.705000 2.770000 1.575000 ;
      RECT 2.500000 1.575000 3.100000 1.955000 ;
      RECT 2.510000 2.250000 3.440000 2.420000 ;
      RECT 2.625000 0.265000 3.740000 0.465000 ;
      RECT 2.950000 0.645000 3.350000 1.015000 ;
      RECT 3.270000 1.230000 3.740000 1.235000 ;
      RECT 3.270000 1.235000 4.770000 1.405000 ;
      RECT 3.270000 1.405000 3.440000 2.250000 ;
      RECT 3.520000 0.465000 3.740000 1.230000 ;
      RECT 3.610000 1.575000 3.910000 1.835000 ;
      RECT 3.610000 1.835000 5.110000 2.085000 ;
      RECT 3.910000 0.735000 4.510000 1.065000 ;
      RECT 4.340000 2.085000 4.510000 2.375000 ;
      RECT 4.470000 1.405000 4.770000 1.565000 ;
      RECT 4.790000 0.295000 4.960000 0.725000 ;
      RECT 4.790000 0.725000 5.110000 1.065000 ;
      RECT 4.940000 1.065000 5.110000 1.835000 ;
      RECT 5.330000 0.725000 6.750000 0.895000 ;
      RECT 5.330000 0.895000 5.500000 1.655000 ;
      RECT 5.330000 1.655000 5.900000 1.965000 ;
      RECT 5.560000 2.165000 6.290000 2.415000 ;
      RECT 5.720000 1.065000 5.900000 1.475000 ;
      RECT 6.070000 1.235000 8.170000 1.405000 ;
      RECT 6.070000 1.405000 6.290000 1.915000 ;
      RECT 6.070000 1.915000 7.380000 2.085000 ;
      RECT 6.070000 2.085000 6.290000 2.165000 ;
      RECT 6.190000 0.305000 7.090000 0.475000 ;
      RECT 6.370000 0.895000 6.750000 1.015000 ;
      RECT 6.460000 1.575000 8.550000 1.745000 ;
      RECT 6.920000 0.475000 7.090000 1.235000 ;
      RECT 7.140000 2.085000 7.380000 2.375000 ;
      RECT 7.260000 0.735000 7.780000 1.005000 ;
      RECT 7.260000 1.005000 7.640000 1.065000 ;
      RECT 7.790000 1.175000 8.170000 1.235000 ;
      RECT 8.210000 0.350000 8.550000 0.680000 ;
      RECT 8.210000 1.745000 8.550000 1.765000 ;
      RECT 8.210000 1.765000 8.380000 2.375000 ;
      RECT 8.340000 0.680000 8.550000 1.575000 ;
      RECT 8.650000 1.915000 8.980000 2.425000 ;
      RECT 8.730000 0.345000 8.900000 0.995000 ;
      RECT 8.730000 0.995000 9.580000 1.325000 ;
      RECT 8.730000 1.325000 8.980000 1.915000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.665000  1.740000  0.835000 1.910000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.165000  0.720000  1.335000 0.890000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.645000  1.740000  2.815000 1.910000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.155000  0.720000  3.325000 0.890000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.280000  0.765000  4.450000 0.935000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.705000  1.740000  5.875000 1.910000 ;
      RECT  5.725000  1.110000  5.895000 1.280000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  0.765000  7.675000 0.935000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 0.605000 1.710000 0.895000 1.800000 ;
      RECT 0.605000 1.800000 5.935000 1.940000 ;
      RECT 1.105000 0.690000 1.395000 0.780000 ;
      RECT 1.105000 0.780000 3.385000 0.920000 ;
      RECT 2.585000 1.710000 2.875000 1.800000 ;
      RECT 3.095000 0.690000 3.385000 0.780000 ;
      RECT 3.170000 0.920000 3.385000 1.120000 ;
      RECT 3.170000 1.120000 5.955000 1.260000 ;
      RECT 5.645000 1.710000 5.935000 1.800000 ;
      RECT 5.665000 1.080000 5.955000 1.120000 ;
      RECT 5.665000 1.260000 5.955000 1.310000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfstp_2


MACRO sky130_fd_sc_hdll__dfstp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.12000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.247200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.870000 1.005000 2.330000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.518200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.740000 1.655000 10.025000 2.325000 ;
        RECT 9.755000 0.265000 10.025000 0.795000 ;
        RECT 9.800000 0.795000 10.025000 1.655000 ;
    END
  END Q
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.220000 0.735000 4.510000 0.780000 ;
        RECT 4.220000 0.780000 7.735000 0.920000 ;
        RECT 4.220000 0.920000 4.510000 0.965000 ;
        RECT 7.445000 0.735000 7.735000 0.780000 ;
        RECT 7.445000 0.920000 7.735000 0.965000 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 0.515000  0.085000  0.895000 0.465000 ;
        RECT 1.555000  0.085000  1.885000 0.465000 ;
        RECT 3.910000  0.085000  4.370000 0.525000 ;
        RECT 5.140000  0.085000  5.530000 0.545000 ;
        RECT 7.320000  0.085000  8.030000 0.565000 ;
        RECT 9.150000  0.085000  9.585000 0.545000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 0.515000 2.135000  0.895000 2.635000 ;
        RECT 1.555000 2.135000  1.885000 2.635000 ;
        RECT 3.730000 2.255000  4.110000 2.635000 ;
        RECT 4.680000 2.255000  5.060000 2.635000 ;
        RECT 6.470000 2.255000  6.940000 2.635000 ;
        RECT 7.710000 1.945000  8.040000 2.635000 ;
        RECT 9.150000 1.835000  9.570000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.345000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 0.890000 0.805000 ;
      RECT 0.175000 1.795000 0.890000 1.965000 ;
      RECT 0.175000 1.965000 0.345000 2.465000 ;
      RECT 0.660000 0.805000 0.890000 1.795000 ;
      RECT 1.115000 0.345000 1.340000 2.465000 ;
      RECT 1.530000 0.635000 2.275000 0.825000 ;
      RECT 1.530000 0.825000 1.700000 1.795000 ;
      RECT 1.530000 1.795000 2.275000 1.965000 ;
      RECT 2.105000 0.305000 2.275000 0.635000 ;
      RECT 2.105000 1.965000 2.275000 2.465000 ;
      RECT 2.500000 0.705000 2.770000 1.575000 ;
      RECT 2.500000 1.575000 3.100000 1.955000 ;
      RECT 2.510000 2.250000 3.440000 2.420000 ;
      RECT 2.625000 0.265000 3.740000 0.465000 ;
      RECT 2.950000 0.645000 3.350000 1.015000 ;
      RECT 3.270000 1.230000 3.740000 1.235000 ;
      RECT 3.270000 1.235000 4.770000 1.405000 ;
      RECT 3.270000 1.405000 3.440000 2.250000 ;
      RECT 3.520000 0.465000 3.740000 1.230000 ;
      RECT 3.610000 1.575000 3.910000 1.835000 ;
      RECT 3.610000 1.835000 5.110000 2.085000 ;
      RECT 3.910000 0.735000 4.510000 1.065000 ;
      RECT 4.340000 2.085000 4.510000 2.375000 ;
      RECT 4.470000 1.405000 4.770000 1.565000 ;
      RECT 4.790000 0.295000 4.960000 0.725000 ;
      RECT 4.790000 0.725000 5.110000 1.065000 ;
      RECT 4.940000 1.065000 5.110000 1.835000 ;
      RECT 5.330000 0.725000 6.750000 0.895000 ;
      RECT 5.330000 0.895000 5.500000 1.655000 ;
      RECT 5.330000 1.655000 5.900000 1.965000 ;
      RECT 5.560000 2.165000 6.290000 2.415000 ;
      RECT 5.720000 1.065000 5.900000 1.475000 ;
      RECT 6.070000 1.235000 8.170000 1.405000 ;
      RECT 6.070000 1.405000 6.290000 1.915000 ;
      RECT 6.070000 1.915000 7.380000 2.085000 ;
      RECT 6.070000 2.085000 6.290000 2.165000 ;
      RECT 6.190000 0.305000 7.090000 0.475000 ;
      RECT 6.370000 0.895000 6.750000 1.015000 ;
      RECT 6.460000 1.575000 8.550000 1.745000 ;
      RECT 6.920000 0.475000 7.090000 1.235000 ;
      RECT 7.140000 2.085000 7.380000 2.375000 ;
      RECT 7.260000 0.735000 7.780000 1.005000 ;
      RECT 7.260000 1.005000 7.640000 1.065000 ;
      RECT 7.790000 1.175000 8.170000 1.235000 ;
      RECT 8.210000 0.350000 8.550000 0.680000 ;
      RECT 8.210000 1.745000 8.550000 1.765000 ;
      RECT 8.210000 1.765000 8.380000 2.375000 ;
      RECT 8.340000 0.680000 8.550000 1.575000 ;
      RECT 8.650000 1.915000 8.980000 2.425000 ;
      RECT 8.730000 0.345000 8.980000 0.995000 ;
      RECT 8.730000 0.995000 9.580000 1.325000 ;
      RECT 8.730000 1.325000 8.980000 1.915000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.665000  1.740000 0.835000 1.910000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.165000  0.720000 1.335000 0.890000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.645000  1.740000 2.815000 1.910000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.155000  0.720000 3.325000 0.890000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.280000  0.765000 4.450000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.705000  1.740000 5.875000 1.910000 ;
      RECT 5.725000  1.110000 5.895000 1.280000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  0.765000 7.675000 0.935000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 0.605000 1.710000 0.895000 1.800000 ;
      RECT 0.605000 1.800000 5.935000 1.940000 ;
      RECT 1.105000 0.690000 1.395000 0.780000 ;
      RECT 1.105000 0.780000 3.385000 0.920000 ;
      RECT 2.585000 1.710000 2.875000 1.800000 ;
      RECT 3.095000 0.690000 3.385000 0.780000 ;
      RECT 3.170000 0.920000 3.385000 1.120000 ;
      RECT 3.170000 1.120000 5.955000 1.260000 ;
      RECT 5.645000 1.710000 5.935000 1.800000 ;
      RECT 5.665000 1.080000 5.955000 1.120000 ;
      RECT 5.665000 1.260000 5.955000 1.310000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfstp_1


MACRO sky130_fd_sc_hdll__tapvgnd_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE WELLTAP ;
  SYMMETRY X Y R90 ;
  SIZE  0.460000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
  END VPWR
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__tapvgnd_1


MACRO sky130_fd_sc_hdll__tapvgnd2_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE WELLTAP ;
  SYMMETRY X Y R90 ;
  SIZE  0.460000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
  END VPWR
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__tapvgnd2_1


MACRO sky130_fd_sc_hdll__diode_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  1.840000 BY  2.720000 ;
  SITE unithd ;
  PIN DIODE
    ANTENNADIFFAREA  1.055700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 1.755000 2.465000 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
  END VPWR
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__diode_4


MACRO sky130_fd_sc_hdll__diode_6
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN DIODE
    ANTENNADIFFAREA  1.718100 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 2.675000 2.465000 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
  END VPWR
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__diode_6


MACRO sky130_fd_sc_hdll__diode_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  0.920000 BY  2.720000 ;
  SITE unithd ;
  PIN DIODE
    ANTENNADIFFAREA  0.434700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.835000 2.465000 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
  END VPWR
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__diode_2


MACRO sky130_fd_sc_hdll__diode_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN DIODE
    ANTENNADIFFAREA  2.352900 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 3.595000 2.465000 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
  END VPWR
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__diode_8


MACRO sky130_fd_sc_hdll__o22a_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.900000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.710000 1.075000 5.130000 1.445000 ;
        RECT 4.710000 1.445000 6.285000 1.615000 ;
        RECT 6.075000 1.075000 6.815000 1.275000 ;
        RECT 6.075000 1.275000 6.285000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.350000 1.075000 5.905000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.620000 1.075000 3.180000 1.445000 ;
        RECT 2.620000 1.445000 4.540000 1.615000 ;
        RECT 4.200000 1.075000 4.540000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 1.075000 4.030000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.725000 1.920000 0.905000 ;
        RECT 0.085000 0.905000 0.370000 1.445000 ;
        RECT 0.085000 1.445000 1.880000 1.615000 ;
        RECT 0.600000 0.265000 0.980000 0.725000 ;
        RECT 0.690000 1.615000 0.940000 2.465000 ;
        RECT 1.540000 0.255000 1.920000 0.725000 ;
        RECT 1.630000 1.615000 1.880000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.220000  1.825000 0.470000 2.635000 ;
      RECT 0.260000  0.085000 0.430000 0.555000 ;
      RECT 0.540000  1.075000 2.430000 1.275000 ;
      RECT 1.160000  1.795000 1.410000 2.635000 ;
      RECT 1.200000  0.085000 1.370000 0.555000 ;
      RECT 2.100000  1.275000 2.430000 1.785000 ;
      RECT 2.100000  1.785000 5.770000 1.955000 ;
      RECT 2.100000  2.125000 2.870000 2.635000 ;
      RECT 2.140000  0.085000 2.310000 0.555000 ;
      RECT 2.140000  0.735000 4.320000 0.905000 ;
      RECT 2.140000  0.905000 2.430000 1.075000 ;
      RECT 2.580000  0.255000 4.870000 0.475000 ;
      RECT 2.615000  0.645000 4.320000 0.735000 ;
      RECT 3.090000  2.125000 3.340000 2.295000 ;
      RECT 3.090000  2.295000 4.280000 2.465000 ;
      RECT 3.560000  1.955000 3.810000 2.125000 ;
      RECT 4.030000  2.125000 4.280000 2.295000 ;
      RECT 4.500000  2.125000 4.830000 2.635000 ;
      RECT 4.540000  0.475000 4.870000 0.735000 ;
      RECT 4.540000  0.735000 6.750000 0.905000 ;
      RECT 5.050000  2.125000 5.300000 2.295000 ;
      RECT 5.050000  2.295000 6.240000 2.465000 ;
      RECT 5.090000  0.085000 5.260000 0.555000 ;
      RECT 5.430000  0.255000 5.810000 0.725000 ;
      RECT 5.430000  0.725000 6.750000 0.735000 ;
      RECT 5.520000  1.955000 5.770000 2.125000 ;
      RECT 5.990000  1.785000 6.240000 2.295000 ;
      RECT 6.030000  0.085000 6.200000 0.555000 ;
      RECT 6.370000  0.255000 6.750000 0.725000 ;
      RECT 6.505000  1.455000 6.710000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22a_4


MACRO sky130_fd_sc_hdll__o22a_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.835000 1.075000 3.310000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335000 1.075000 2.665000 1.325000 ;
        RECT 2.445000 1.325000 2.665000 2.405000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.535000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.730000 1.075000 2.155000 1.325000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.472000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.365000 0.365000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.535000  0.715000 1.805000 0.895000 ;
      RECT 0.535000  0.895000 0.860000 1.495000 ;
      RECT 0.535000  1.495000 2.275000 1.705000 ;
      RECT 0.605000  1.875000 1.360000 2.635000 ;
      RECT 0.615000  0.085000 0.785000 0.545000 ;
      RECT 1.055000  0.295000 2.395000 0.475000 ;
      RECT 1.440000  0.645000 1.805000 0.715000 ;
      RECT 1.805000  1.705000 2.275000 2.465000 ;
      RECT 2.065000  0.475000 2.395000 0.695000 ;
      RECT 2.065000  0.695000 3.355000 0.865000 ;
      RECT 2.625000  0.085000 2.795000 0.525000 ;
      RECT 2.965000  0.280000 3.355000 0.695000 ;
      RECT 2.985000  1.455000 3.540000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22a_1


MACRO sky130_fd_sc_hdll__o22a_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.345000 1.075000 3.705000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.795000 1.075000 3.175000 1.275000 ;
        RECT 2.905000 1.275000 3.175000 2.405000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.075000 1.890000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 1.075000 2.625000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.491500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.365000 0.855000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.115000  1.445000 0.365000 2.635000 ;
      RECT 0.185000  0.085000 0.355000 0.885000 ;
      RECT 1.075000  0.715000 2.365000 0.895000 ;
      RECT 1.075000  0.895000 1.355000 1.455000 ;
      RECT 1.075000  1.455000 2.695000 1.705000 ;
      RECT 1.095000  1.875000 1.895000 2.635000 ;
      RECT 1.125000  0.085000 1.305000 0.545000 ;
      RECT 1.565000  0.295000 2.930000 0.475000 ;
      RECT 1.950000  0.645000 2.365000 0.715000 ;
      RECT 2.340000  1.705000 2.695000 2.465000 ;
      RECT 2.590000  0.475000 2.930000 0.695000 ;
      RECT 2.590000  0.695000 3.890000 0.865000 ;
      RECT 3.195000  0.085000 3.365000 0.525000 ;
      RECT 3.555000  0.280000 3.890000 0.695000 ;
      RECT 3.570000  1.795000 3.890000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22a_2


MACRO sky130_fd_sc_hdll__dfrtp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.12000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.615000 1.905000 1.665000 ;
        RECT 1.455000 1.665000 1.770000 2.005000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.150000 0.255000  9.530000 0.735000 ;
        RECT 9.150000 0.735000 10.010000 0.905000 ;
        RECT 9.240000 1.455000 10.010000 1.625000 ;
        RECT 9.240000 1.625000  9.530000 2.465000 ;
        RECT 9.625000 0.905000 10.010000 1.455000 ;
    END
  END Q
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.995000 0.735000 4.745000 0.780000 ;
        RECT 3.995000 0.780000 7.865000 0.920000 ;
        RECT 3.995000 0.920000 4.745000 0.965000 ;
        RECT 7.575000 0.735000 7.865000 0.780000 ;
        RECT 7.575000 0.920000 7.865000 0.965000 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.090000  0.345000  0.345000 0.635000 ;
      RECT 0.090000  0.635000  0.890000 0.805000 ;
      RECT 0.090000  1.795000  0.890000 1.965000 ;
      RECT 0.090000  1.965000  0.345000 2.465000 ;
      RECT 0.515000  0.085000  0.895000 0.465000 ;
      RECT 0.515000  2.135000  0.895000 2.635000 ;
      RECT 0.660000  0.805000  0.890000 1.795000 ;
      RECT 1.115000  0.345000  1.285000 2.465000 ;
      RECT 1.575000  0.085000  1.905000 0.445000 ;
      RECT 1.770000  2.175000  1.940000 2.635000 ;
      RECT 2.075000  0.305000  2.495000 0.475000 ;
      RECT 2.075000  0.475000  2.245000 1.835000 ;
      RECT 2.075000  1.835000  2.340000 2.005000 ;
      RECT 2.170000  2.005000  2.340000 2.135000 ;
      RECT 2.170000  2.135000  2.420000 2.465000 ;
      RECT 2.425000  0.765000  2.685000 1.385000 ;
      RECT 2.510000  1.575000  3.025000 1.965000 ;
      RECT 2.685000  2.135000  3.365000 2.465000 ;
      RECT 2.695000  0.305000  3.600000 0.475000 ;
      RECT 2.855000  0.765000  3.210000 0.985000 ;
      RECT 2.855000  0.985000  3.025000 1.575000 ;
      RECT 3.195000  1.185000  4.985000 1.355000 ;
      RECT 3.195000  1.355000  3.365000 2.135000 ;
      RECT 3.430000  0.475000  3.600000 1.185000 ;
      RECT 3.535000  1.865000  4.710000 2.035000 ;
      RECT 3.535000  2.035000  3.705000 2.375000 ;
      RECT 3.725000  1.525000  5.325000 1.695000 ;
      RECT 3.805000  0.765000  4.645000 1.015000 ;
      RECT 3.990000  2.205000  4.320000 2.635000 ;
      RECT 4.525000  0.085000  4.855000 0.545000 ;
      RECT 4.540000  2.035000  4.710000 2.375000 ;
      RECT 4.815000  1.005000  4.985000 1.185000 ;
      RECT 5.005000  2.175000  5.425000 2.635000 ;
      RECT 5.065000  0.275000  5.465000 0.445000 ;
      RECT 5.065000  0.445000  5.325000 0.835000 ;
      RECT 5.155000  0.835000  5.325000 1.525000 ;
      RECT 5.155000  1.695000  5.325000 1.835000 ;
      RECT 5.155000  1.835000  5.815000 2.005000 ;
      RECT 5.605000  0.705000  5.775000 1.495000 ;
      RECT 5.605000  1.495000  6.315000 1.655000 ;
      RECT 5.605000  1.655000  6.660000 1.665000 ;
      RECT 5.645000  2.005000  5.815000 2.465000 ;
      RECT 5.735000  0.255000  6.655000 0.535000 ;
      RECT 5.945000  0.705000  6.315000 1.325000 ;
      RECT 6.050000  2.125000  7.005000 2.465000 ;
      RECT 6.145000  1.665000  6.660000 1.955000 ;
      RECT 6.485000  0.535000  6.655000 1.315000 ;
      RECT 6.485000  1.315000  7.055000 1.485000 ;
      RECT 6.825000  0.085000  6.995000 0.525000 ;
      RECT 6.835000  1.485000  7.055000 1.575000 ;
      RECT 6.835000  1.575000  8.270000 1.745000 ;
      RECT 6.835000  1.745000  7.005000 2.125000 ;
      RECT 6.955000  0.695000  7.335000 0.865000 ;
      RECT 6.955000  0.865000  7.225000 1.145000 ;
      RECT 7.165000  0.295000  8.635000 0.465000 ;
      RECT 7.165000  0.465000  7.335000 0.695000 ;
      RECT 7.340000  2.175000  7.590000 2.635000 ;
      RECT 7.505000  0.635000  7.905000 1.405000 ;
      RECT 7.810000  1.915000  8.610000 2.085000 ;
      RECT 7.810000  2.085000  7.980000 2.375000 ;
      RECT 8.160000  2.255000  8.540000 2.635000 ;
      RECT 8.290000  0.465000  8.635000 1.075000 ;
      RECT 8.290000  1.075000  9.335000 1.285000 ;
      RECT 8.290000  1.285000  8.610000 1.295000 ;
      RECT 8.440000  1.295000  8.610000 1.915000 ;
      RECT 8.810000  0.085000  8.980000 0.895000 ;
      RECT 8.810000  1.575000  8.980000 2.635000 ;
      RECT 9.750000  0.085000  9.920000 0.555000 ;
      RECT 9.750000  1.795000  9.920000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.660000  1.105000 0.830000 1.275000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.115000  1.785000 1.285000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.480000  1.105000 2.650000 1.275000 ;
      RECT 2.725000  1.785000 2.895000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.105000  0.765000 4.275000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.465000  0.765000 4.635000 0.935000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.020000  1.105000 6.190000 1.275000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.470000  1.785000 6.640000 1.955000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.635000  0.765000 7.805000 0.935000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 0.600000 1.075000 0.890000 1.120000 ;
      RECT 0.600000 1.120000 6.250000 1.260000 ;
      RECT 0.600000 1.260000 0.890000 1.305000 ;
      RECT 1.005000 1.755000 1.345000 1.800000 ;
      RECT 1.005000 1.800000 6.700000 1.940000 ;
      RECT 1.005000 1.940000 1.345000 1.985000 ;
      RECT 2.420000 1.075000 2.710000 1.120000 ;
      RECT 2.420000 1.260000 2.710000 1.305000 ;
      RECT 2.665000 1.755000 2.955000 1.800000 ;
      RECT 2.665000 1.940000 2.955000 1.985000 ;
      RECT 5.960000 1.075000 6.250000 1.120000 ;
      RECT 5.960000 1.260000 6.250000 1.305000 ;
      RECT 6.410000 1.755000 6.700000 1.800000 ;
      RECT 6.410000 1.940000 6.700000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfrtp_2


MACRO sky130_fd_sc_hdll__dfrtp_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.50000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.615000 1.975000 1.665000 ;
        RECT 1.455000 1.665000 1.780000 2.450000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.475000 0.255000  9.855000 0.735000 ;
        RECT  9.475000 0.735000 11.405000 0.905000 ;
        RECT  9.565000 1.455000 11.405000 1.625000 ;
        RECT  9.565000 1.625000  9.855000 2.465000 ;
        RECT 10.415000 0.255000 10.795000 0.735000 ;
        RECT 10.505000 1.625000 10.755000 2.465000 ;
        RECT 10.995000 0.905000 11.405000 1.455000 ;
    END
  END Q
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.175000 0.735000 4.925000 0.780000 ;
        RECT 4.175000 0.780000 8.395000 0.920000 ;
        RECT 4.175000 0.920000 4.925000 0.965000 ;
        RECT 7.810000 0.920000 8.395000 1.280000 ;
        RECT 8.105000 0.735000 8.395000 0.780000 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.500000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.500000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.500000 0.085000 ;
      RECT  0.000000  2.635000 11.500000 2.805000 ;
      RECT  0.090000  0.345000  0.345000 0.635000 ;
      RECT  0.090000  0.635000  0.890000 0.805000 ;
      RECT  0.090000  1.795000  0.890000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.515000  2.135000  0.895000 2.635000 ;
      RECT  0.660000  0.805000  0.890000 1.795000 ;
      RECT  1.115000  0.345000  1.285000 2.465000 ;
      RECT  1.645000  0.085000  1.975000 0.445000 ;
      RECT  1.950000  2.175000  2.200000 2.635000 ;
      RECT  2.145000  0.305000  2.690000 0.475000 ;
      RECT  2.145000  0.475000  2.315000 1.835000 ;
      RECT  2.145000  1.835000  2.590000 2.005000 ;
      RECT  2.420000  2.005000  2.590000 2.135000 ;
      RECT  2.420000  2.135000  2.670000 2.465000 ;
      RECT  2.535000  0.765000  2.935000 1.385000 ;
      RECT  2.760000  1.575000  3.275000 1.965000 ;
      RECT  2.935000  2.135000  3.665000 2.465000 ;
      RECT  2.945000  0.305000  3.850000 0.475000 ;
      RECT  3.105000  0.765000  3.510000 0.985000 ;
      RECT  3.105000  0.985000  3.275000 1.575000 ;
      RECT  3.495000  1.185000  5.285000 1.355000 ;
      RECT  3.495000  1.355000  3.665000 2.135000 ;
      RECT  3.680000  0.475000  3.850000 1.185000 ;
      RECT  3.835000  1.865000  5.010000 2.035000 ;
      RECT  3.835000  2.035000  4.005000 2.375000 ;
      RECT  4.025000  1.525000  5.675000 1.695000 ;
      RECT  4.175000  0.765000  4.945000 1.015000 ;
      RECT  4.290000  2.205000  4.620000 2.635000 ;
      RECT  4.825000  0.085000  5.155000 0.545000 ;
      RECT  4.840000  2.035000  5.010000 2.375000 ;
      RECT  5.115000  1.005000  5.285000 1.185000 ;
      RECT  5.305000  2.175000  5.725000 2.635000 ;
      RECT  5.365000  0.275000  5.765000 0.445000 ;
      RECT  5.365000  0.445000  5.675000 0.835000 ;
      RECT  5.505000  0.835000  5.675000 1.525000 ;
      RECT  5.505000  1.695000  5.675000 1.835000 ;
      RECT  5.505000  1.835000  6.115000 2.005000 ;
      RECT  5.915000  0.705000  6.125000 1.495000 ;
      RECT  5.915000  1.495000  6.690000 1.655000 ;
      RECT  5.915000  1.655000  7.030000 1.665000 ;
      RECT  5.945000  2.005000  6.115000 2.465000 ;
      RECT  6.035000  0.255000  7.135000 0.535000 ;
      RECT  6.295000  0.705000  6.745000 1.325000 ;
      RECT  6.350000  2.125000  7.470000 2.465000 ;
      RECT  6.470000  1.665000  7.030000 1.955000 ;
      RECT  6.965000  0.535000  7.135000 1.315000 ;
      RECT  6.965000  1.315000  7.470000 1.485000 ;
      RECT  7.250000  1.485000  7.470000 1.575000 ;
      RECT  7.250000  1.575000  8.620000 1.745000 ;
      RECT  7.250000  1.745000  7.470000 2.125000 ;
      RECT  7.355000  0.085000  7.595000 0.525000 ;
      RECT  7.355000  0.695000  7.935000 0.865000 ;
      RECT  7.355000  0.865000  7.625000 1.145000 ;
      RECT  7.640000  2.175000  7.890000 2.635000 ;
      RECT  7.765000  0.295000  8.935000 0.465000 ;
      RECT  7.765000  0.465000  7.935000 0.695000 ;
      RECT  7.805000  1.035000  8.395000 1.405000 ;
      RECT  8.110000  1.915000  8.960000 2.085000 ;
      RECT  8.110000  2.085000  8.280000 2.375000 ;
      RECT  8.155000  0.635000  8.395000 1.035000 ;
      RECT  8.460000  2.255000  8.840000 2.635000 ;
      RECT  8.615000  0.465000  8.935000 0.820000 ;
      RECT  8.615000  0.820000  8.940000 1.075000 ;
      RECT  8.615000  1.075000 10.795000 1.285000 ;
      RECT  8.615000  1.285000  8.960000 1.295000 ;
      RECT  8.790000  1.295000  8.960000 1.915000 ;
      RECT  9.135000  0.085000  9.305000 0.895000 ;
      RECT  9.135000  1.575000  9.305000 2.635000 ;
      RECT 10.075000  0.085000 10.245000 0.555000 ;
      RECT 10.075000  1.795000 10.245000 2.635000 ;
      RECT 11.015000  0.085000 11.185000 0.555000 ;
      RECT 11.015000  1.795000 11.185000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.660000  1.105000  0.830000 1.275000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.115000  1.785000  1.285000 1.955000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.595000  1.105000  2.765000 1.275000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.105000  1.785000  3.275000 1.955000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  0.765000  4.455000 0.935000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.645000  0.765000  4.815000 0.935000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.525000  1.105000  6.695000 1.275000 ;
      RECT  6.525000  1.785000  6.695000 1.955000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.870000  1.080000  8.040000 1.250000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.165000  0.765000  8.335000 0.935000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
    LAYER met1 ;
      RECT 0.600000 1.075000 0.890000 1.120000 ;
      RECT 0.600000 1.120000 6.805000 1.260000 ;
      RECT 0.600000 1.260000 0.890000 1.305000 ;
      RECT 1.005000 1.755000 1.345000 1.800000 ;
      RECT 1.005000 1.800000 6.805000 1.940000 ;
      RECT 1.005000 1.940000 1.345000 1.985000 ;
      RECT 2.535000 1.075000 2.825000 1.120000 ;
      RECT 2.535000 1.260000 2.825000 1.305000 ;
      RECT 3.045000 1.755000 3.335000 1.800000 ;
      RECT 3.045000 1.940000 3.335000 1.985000 ;
      RECT 6.465000 1.075000 6.805000 1.120000 ;
      RECT 6.465000 1.260000 6.805000 1.305000 ;
      RECT 6.465000 1.755000 6.805000 1.800000 ;
      RECT 6.465000 1.940000 6.805000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfrtp_4


MACRO sky130_fd_sc_hdll__dfrtp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.660000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.615000 1.905000 1.665000 ;
        RECT 1.455000 1.665000 1.770000 2.005000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.472000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.240000 0.255000 9.575000 2.465000 ;
    END
  END Q
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.995000 0.735000 4.745000 0.780000 ;
        RECT 3.995000 0.780000 7.865000 0.920000 ;
        RECT 3.995000 0.920000 4.745000 0.965000 ;
        RECT 7.575000 0.735000 7.865000 0.780000 ;
        RECT 7.575000 0.920000 7.865000 0.965000 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.090000  0.345000 0.345000 0.635000 ;
      RECT 0.090000  0.635000 0.890000 0.805000 ;
      RECT 0.090000  1.795000 0.890000 1.965000 ;
      RECT 0.090000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.895000 0.465000 ;
      RECT 0.515000  2.135000 0.895000 2.635000 ;
      RECT 0.660000  0.805000 0.890000 1.795000 ;
      RECT 1.115000  0.345000 1.285000 2.465000 ;
      RECT 1.575000  0.085000 1.905000 0.445000 ;
      RECT 1.770000  2.175000 1.940000 2.635000 ;
      RECT 2.075000  0.305000 2.495000 0.475000 ;
      RECT 2.075000  0.475000 2.245000 1.835000 ;
      RECT 2.075000  1.835000 2.340000 2.005000 ;
      RECT 2.170000  2.005000 2.340000 2.135000 ;
      RECT 2.170000  2.135000 2.420000 2.465000 ;
      RECT 2.425000  0.765000 2.685000 1.385000 ;
      RECT 2.510000  1.575000 3.025000 1.965000 ;
      RECT 2.685000  2.135000 3.365000 2.465000 ;
      RECT 2.695000  0.305000 3.600000 0.475000 ;
      RECT 2.855000  0.765000 3.210000 0.985000 ;
      RECT 2.855000  0.985000 3.025000 1.575000 ;
      RECT 3.195000  1.185000 4.985000 1.355000 ;
      RECT 3.195000  1.355000 3.365000 2.135000 ;
      RECT 3.430000  0.475000 3.600000 1.185000 ;
      RECT 3.535000  1.865000 4.710000 2.035000 ;
      RECT 3.535000  2.035000 3.705000 2.375000 ;
      RECT 3.725000  1.525000 5.325000 1.695000 ;
      RECT 3.805000  0.765000 4.645000 1.015000 ;
      RECT 3.990000  2.205000 4.320000 2.635000 ;
      RECT 4.525000  0.085000 4.855000 0.545000 ;
      RECT 4.540000  2.035000 4.710000 2.375000 ;
      RECT 4.815000  1.005000 4.985000 1.185000 ;
      RECT 5.005000  2.175000 5.425000 2.635000 ;
      RECT 5.065000  0.275000 5.465000 0.445000 ;
      RECT 5.065000  0.445000 5.325000 0.835000 ;
      RECT 5.155000  0.835000 5.325000 1.525000 ;
      RECT 5.155000  1.695000 5.325000 1.835000 ;
      RECT 5.155000  1.835000 5.815000 2.005000 ;
      RECT 5.605000  0.705000 5.775000 1.495000 ;
      RECT 5.605000  1.495000 6.315000 1.655000 ;
      RECT 5.605000  1.655000 6.660000 1.665000 ;
      RECT 5.645000  2.005000 5.815000 2.465000 ;
      RECT 5.735000  0.255000 6.655000 0.535000 ;
      RECT 5.945000  0.705000 6.315000 1.325000 ;
      RECT 6.050000  2.125000 7.005000 2.465000 ;
      RECT 6.145000  1.665000 6.660000 1.955000 ;
      RECT 6.485000  0.535000 6.655000 1.315000 ;
      RECT 6.485000  1.315000 7.055000 1.485000 ;
      RECT 6.825000  0.085000 6.995000 0.525000 ;
      RECT 6.835000  1.485000 7.055000 1.575000 ;
      RECT 6.835000  1.575000 8.270000 1.745000 ;
      RECT 6.835000  1.745000 7.005000 2.125000 ;
      RECT 6.955000  0.695000 7.335000 0.865000 ;
      RECT 6.955000  0.865000 7.225000 1.145000 ;
      RECT 7.165000  0.295000 8.635000 0.465000 ;
      RECT 7.165000  0.465000 7.335000 0.695000 ;
      RECT 7.340000  2.175000 7.590000 2.635000 ;
      RECT 7.505000  0.635000 7.905000 1.405000 ;
      RECT 7.810000  1.915000 8.610000 2.085000 ;
      RECT 7.810000  2.085000 7.980000 2.375000 ;
      RECT 8.160000  2.255000 8.540000 2.635000 ;
      RECT 8.290000  0.465000 8.635000 1.075000 ;
      RECT 8.290000  1.075000 9.070000 1.285000 ;
      RECT 8.290000  1.285000 8.610000 1.295000 ;
      RECT 8.440000  1.295000 8.610000 1.915000 ;
      RECT 8.810000  0.085000 8.980000 0.895000 ;
      RECT 8.810000  1.575000 8.980000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.660000  1.105000 0.830000 1.275000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.115000  1.785000 1.285000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.480000  1.105000 2.650000 1.275000 ;
      RECT 2.725000  1.785000 2.895000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.105000  0.765000 4.275000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.465000  0.765000 4.635000 0.935000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.020000  1.105000 6.190000 1.275000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.470000  1.785000 6.640000 1.955000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.635000  0.765000 7.805000 0.935000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.600000 1.075000 0.890000 1.120000 ;
      RECT 0.600000 1.120000 6.250000 1.260000 ;
      RECT 0.600000 1.260000 0.890000 1.305000 ;
      RECT 1.005000 1.755000 1.345000 1.800000 ;
      RECT 1.005000 1.800000 6.700000 1.940000 ;
      RECT 1.005000 1.940000 1.345000 1.985000 ;
      RECT 2.420000 1.075000 2.710000 1.120000 ;
      RECT 2.420000 1.260000 2.710000 1.305000 ;
      RECT 2.665000 1.755000 2.955000 1.800000 ;
      RECT 2.665000 1.940000 2.955000 1.985000 ;
      RECT 5.960000 1.075000 6.250000 1.120000 ;
      RECT 5.960000 1.260000 6.250000 1.305000 ;
      RECT 6.410000 1.755000 6.700000 1.800000 ;
      RECT 6.410000 1.940000 6.700000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfrtp_1


MACRO sky130_fd_sc_hdll__sdfrtp_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  14.26000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.160200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.120000 1.355000 3.655000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.171500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.425000 0.265000 12.755000 0.995000 ;
        RECT 12.425000 0.995000 13.695000 1.325000 ;
        RECT 12.425000 1.325000 12.755000 2.325000 ;
        RECT 13.445000 0.265000 13.695000 0.995000 ;
        RECT 13.445000 1.325000 13.695000 2.325000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.145000 0.735000  7.900000 0.780000 ;
        RECT  7.145000 0.780000 11.405000 0.920000 ;
        RECT  7.145000 0.920000  7.900000 0.965000 ;
        RECT 10.775000 0.920000 11.405000 0.965000 ;
        RECT 10.775000 0.965000 11.065000 1.310000 ;
        RECT 11.115000 0.735000 11.405000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.172800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.610000 0.710000 4.955000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.467400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.070000 1.990000 1.335000 ;
        RECT 1.585000 1.335000 2.220000 1.745000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.090000  1.795000  0.915000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.885000 0.805000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.530000  2.135000  0.910000 2.635000 ;
      RECT  0.710000  0.805000  0.885000 0.995000 ;
      RECT  0.710000  0.995000  1.025000 1.325000 ;
      RECT  0.710000  1.325000  0.915000 1.795000 ;
      RECT  1.115000  0.345000  1.365000 0.675000 ;
      RECT  1.135000  1.730000  1.365000 2.465000 ;
      RECT  1.195000  0.675000  1.365000 1.730000 ;
      RECT  1.695000  0.395000  1.865000 0.730000 ;
      RECT  1.695000  0.730000  2.435000 0.900000 ;
      RECT  2.035000  0.085000  2.415000 0.560000 ;
      RECT  2.110000  1.915000  2.730000 2.085000 ;
      RECT  2.110000  2.085000  2.380000 2.400000 ;
      RECT  2.265000  0.900000  2.435000 0.995000 ;
      RECT  2.265000  0.995000  3.445000 1.165000 ;
      RECT  2.475000  1.165000  3.445000 1.185000 ;
      RECT  2.475000  1.185000  2.730000 1.915000 ;
      RECT  2.600000  2.255000  2.930000 2.635000 ;
      RECT  2.655000  0.085000  3.035000 0.825000 ;
      RECT  3.275000  0.255000  4.435000 0.425000 ;
      RECT  3.275000  0.425000  3.445000 0.995000 ;
      RECT  3.665000  0.675000  4.045000 1.075000 ;
      RECT  3.870000  1.075000  4.045000 1.935000 ;
      RECT  3.870000  1.935000  5.650000 2.105000 ;
      RECT  3.870000  2.105000  4.040000 2.465000 ;
      RECT  4.265000  0.425000  4.435000 1.685000 ;
      RECT  4.855000  2.275000  5.205000 2.635000 ;
      RECT  5.005000  0.085000  5.350000 0.540000 ;
      RECT  5.140000  0.715000  5.720000 0.895000 ;
      RECT  5.140000  0.895000  5.310000 1.935000 ;
      RECT  5.480000  1.065000  5.650000 1.395000 ;
      RECT  5.480000  2.105000  5.650000 2.185000 ;
      RECT  5.480000  2.185000  5.850000 2.435000 ;
      RECT  5.550000  0.335000  5.890000 0.505000 ;
      RECT  5.550000  0.505000  5.720000 0.715000 ;
      RECT  5.820000  1.575000  6.120000 1.955000 ;
      RECT  5.900000  0.705000  6.650000 1.035000 ;
      RECT  5.900000  1.035000  6.120000 1.575000 ;
      RECT  6.095000  2.135000  6.460000 2.465000 ;
      RECT  6.110000  0.305000  7.010000 0.475000 ;
      RECT  6.290000  1.215000  8.150000 1.385000 ;
      RECT  6.290000  1.385000  6.460000 2.135000 ;
      RECT  6.680000  1.935000  7.940000 2.105000 ;
      RECT  6.680000  2.105000  6.850000 2.375000 ;
      RECT  6.840000  0.475000  7.010000 1.215000 ;
      RECT  6.960000  1.595000  8.540000 1.765000 ;
      RECT  7.135000  2.355000  7.465000 2.635000 ;
      RECT  7.230000  0.765000  7.810000 1.045000 ;
      RECT  7.690000  0.085000  8.020000 0.545000 ;
      RECT  7.770000  2.105000  7.940000 2.375000 ;
      RECT  7.980000  1.005000  8.150000 1.215000 ;
      RECT  8.150000  2.175000  8.570000 2.635000 ;
      RECT  8.230000  0.275000  8.610000 0.445000 ;
      RECT  8.230000  0.445000  8.540000 0.835000 ;
      RECT  8.230000  1.765000  8.540000 1.835000 ;
      RECT  8.230000  1.835000  8.985000 2.005000 ;
      RECT  8.370000  0.835000  8.540000 1.595000 ;
      RECT  8.710000  0.705000  8.970000 1.495000 ;
      RECT  8.710000  1.495000  9.445000 1.660000 ;
      RECT  8.710000  1.660000  9.845000 1.665000 ;
      RECT  8.780000  0.255000  9.890000 0.535000 ;
      RECT  8.815000  2.005000  8.985000 2.465000 ;
      RECT  9.185000  1.665000  9.845000 1.955000 ;
      RECT  9.195000  2.125000 10.215000 2.465000 ;
      RECT  9.235000  0.920000  9.405000 1.325000 ;
      RECT  9.670000  0.535000  9.890000 1.315000 ;
      RECT  9.670000  1.315000 10.285000 1.485000 ;
      RECT 10.040000  1.485000 10.285000 1.575000 ;
      RECT 10.040000  1.575000 11.370000 1.745000 ;
      RECT 10.040000  1.745000 10.215000 2.125000 ;
      RECT 10.110000  0.085000 10.330000 0.525000 ;
      RECT 10.150000  0.695000 10.730000 0.865000 ;
      RECT 10.150000  0.865000 10.370000 1.145000 ;
      RECT 10.415000  2.195000 10.665000 2.635000 ;
      RECT 10.560000  0.295000 11.735000 0.465000 ;
      RECT 10.560000  0.465000 10.730000 0.695000 ;
      RECT 10.600000  1.065000 11.370000 1.275000 ;
      RECT 10.910000  1.915000 11.730000 2.085000 ;
      RECT 10.910000  2.085000 11.080000 2.375000 ;
      RECT 11.065000  0.635000 11.370000 1.065000 ;
      RECT 11.255000  2.255000 11.635000 2.635000 ;
      RECT 11.560000  0.465000 11.735000 0.995000 ;
      RECT 11.560000  0.995000 12.205000 1.325000 ;
      RECT 11.560000  1.325000 11.730000 1.915000 ;
      RECT 11.905000  0.085000 12.075000 0.545000 ;
      RECT 11.905000  1.495000 12.155000 2.635000 ;
      RECT 12.975000  0.085000 13.145000 0.545000 ;
      RECT 12.975000  1.495000 13.225000 2.635000 ;
      RECT 13.915000  0.085000 14.085000 0.545000 ;
      RECT 13.915000  1.495000 14.165000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.855000  1.105000  1.025000 1.275000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.135000  1.785000  1.305000 1.955000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.480000  1.105000  5.650000 1.275000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.950000  1.785000  6.120000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.255000  0.765000  7.425000 0.935000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.615000  0.765000  7.785000 0.935000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.235000  1.105000  9.405000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.565000  1.785000  9.735000 1.955000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.835000  1.085000 11.005000 1.255000 ;
      RECT 11.175000  0.765000 11.345000 0.935000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT 0.795000 1.075000 1.085000 1.120000 ;
      RECT 0.795000 1.120000 9.465000 1.260000 ;
      RECT 0.795000 1.260000 1.085000 1.305000 ;
      RECT 1.070000 1.755000 1.370000 1.800000 ;
      RECT 1.070000 1.800000 9.795000 1.940000 ;
      RECT 1.070000 1.940000 1.370000 1.985000 ;
      RECT 5.420000 1.075000 5.710000 1.120000 ;
      RECT 5.420000 1.260000 5.710000 1.305000 ;
      RECT 5.890000 1.755000 6.180000 1.800000 ;
      RECT 5.890000 1.940000 6.180000 1.985000 ;
      RECT 9.155000 1.075000 9.465000 1.120000 ;
      RECT 9.155000 1.260000 9.465000 1.305000 ;
      RECT 9.500000 1.755000 9.795000 1.800000 ;
      RECT 9.500000 1.940000 9.795000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrtp_4


MACRO sky130_fd_sc_hdll__sdfrtp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  13.34000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.160200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.120000 1.355000 3.655000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.500000 0.265000 12.785000 2.325000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.145000 0.735000  7.900000 0.780000 ;
        RECT  7.145000 0.780000 11.370000 0.920000 ;
        RECT  7.145000 0.920000  7.900000 0.965000 ;
        RECT 11.080000 0.735000 11.370000 0.780000 ;
        RECT 11.080000 0.920000 11.370000 0.965000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.172800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.610000 0.710000 4.955000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.467400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.070000 1.990000 1.335000 ;
        RECT 1.585000 1.335000 2.220000 1.745000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.340000 0.085000 ;
      RECT  0.000000  2.635000 13.340000 2.805000 ;
      RECT  0.090000  1.795000  0.915000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.885000 0.805000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.530000  2.135000  0.910000 2.635000 ;
      RECT  0.710000  0.805000  0.885000 0.995000 ;
      RECT  0.710000  0.995000  1.025000 1.325000 ;
      RECT  0.710000  1.325000  0.915000 1.795000 ;
      RECT  1.115000  0.345000  1.365000 0.675000 ;
      RECT  1.135000  1.730000  1.365000 2.465000 ;
      RECT  1.195000  0.675000  1.365000 1.730000 ;
      RECT  1.695000  0.395000  1.865000 0.730000 ;
      RECT  1.695000  0.730000  2.435000 0.900000 ;
      RECT  2.035000  0.085000  2.415000 0.560000 ;
      RECT  2.110000  1.915000  2.730000 2.085000 ;
      RECT  2.110000  2.085000  2.380000 2.400000 ;
      RECT  2.265000  0.900000  2.435000 0.995000 ;
      RECT  2.265000  0.995000  3.445000 1.165000 ;
      RECT  2.475000  1.165000  3.445000 1.185000 ;
      RECT  2.475000  1.185000  2.730000 1.915000 ;
      RECT  2.600000  2.255000  2.930000 2.635000 ;
      RECT  2.655000  0.085000  3.035000 0.825000 ;
      RECT  3.275000  0.255000  4.435000 0.425000 ;
      RECT  3.275000  0.425000  3.445000 0.995000 ;
      RECT  3.665000  0.675000  4.045000 1.075000 ;
      RECT  3.870000  1.075000  4.045000 1.935000 ;
      RECT  3.870000  1.935000  5.650000 2.105000 ;
      RECT  3.870000  2.105000  4.040000 2.465000 ;
      RECT  4.265000  0.425000  4.435000 1.685000 ;
      RECT  4.855000  2.275000  5.205000 2.635000 ;
      RECT  5.005000  0.085000  5.350000 0.540000 ;
      RECT  5.140000  0.715000  5.720000 0.895000 ;
      RECT  5.140000  0.895000  5.310000 1.935000 ;
      RECT  5.480000  1.065000  5.650000 1.395000 ;
      RECT  5.480000  2.105000  5.650000 2.185000 ;
      RECT  5.480000  2.185000  5.850000 2.435000 ;
      RECT  5.550000  0.335000  5.890000 0.505000 ;
      RECT  5.550000  0.505000  5.720000 0.715000 ;
      RECT  5.820000  1.575000  6.120000 1.955000 ;
      RECT  5.900000  0.705000  6.650000 1.035000 ;
      RECT  5.900000  1.035000  6.120000 1.575000 ;
      RECT  6.095000  2.135000  6.460000 2.465000 ;
      RECT  6.110000  0.305000  7.010000 0.475000 ;
      RECT  6.290000  1.215000  8.150000 1.385000 ;
      RECT  6.290000  1.385000  6.460000 2.135000 ;
      RECT  6.680000  1.935000  7.940000 2.105000 ;
      RECT  6.680000  2.105000  6.850000 2.375000 ;
      RECT  6.840000  0.475000  7.010000 1.215000 ;
      RECT  6.960000  1.595000  8.540000 1.765000 ;
      RECT  7.135000  2.355000  7.465000 2.635000 ;
      RECT  7.230000  0.765000  7.810000 1.045000 ;
      RECT  7.690000  0.085000  8.020000 0.545000 ;
      RECT  7.770000  2.105000  7.940000 2.375000 ;
      RECT  7.980000  1.005000  8.150000 1.215000 ;
      RECT  8.150000  2.175000  8.570000 2.635000 ;
      RECT  8.230000  0.275000  8.610000 0.445000 ;
      RECT  8.230000  0.445000  8.540000 0.835000 ;
      RECT  8.230000  1.765000  8.540000 1.835000 ;
      RECT  8.230000  1.835000  8.985000 2.005000 ;
      RECT  8.370000  0.835000  8.540000 1.595000 ;
      RECT  8.710000  0.705000  8.970000 1.495000 ;
      RECT  8.710000  1.495000  9.445000 1.660000 ;
      RECT  8.710000  1.660000  9.845000 1.665000 ;
      RECT  8.780000  0.255000  9.890000 0.535000 ;
      RECT  8.815000  2.005000  8.985000 2.465000 ;
      RECT  9.185000  1.665000  9.845000 1.955000 ;
      RECT  9.195000  2.125000 10.215000 2.465000 ;
      RECT  9.235000  0.920000  9.405000 1.325000 ;
      RECT  9.670000  0.535000  9.890000 1.315000 ;
      RECT  9.670000  1.315000 10.285000 1.485000 ;
      RECT 10.040000  1.485000 10.285000 1.575000 ;
      RECT 10.040000  1.575000 11.370000 1.745000 ;
      RECT 10.040000  1.745000 10.215000 2.125000 ;
      RECT 10.110000  0.085000 10.330000 0.525000 ;
      RECT 10.150000  0.695000 10.730000 0.865000 ;
      RECT 10.150000  0.865000 10.370000 1.145000 ;
      RECT 10.415000  2.195000 10.665000 2.635000 ;
      RECT 10.560000  0.295000 11.735000 0.465000 ;
      RECT 10.560000  0.465000 10.730000 0.695000 ;
      RECT 10.600000  1.065000 11.370000 1.275000 ;
      RECT 10.910000  1.915000 11.730000 2.085000 ;
      RECT 10.910000  2.085000 11.080000 2.375000 ;
      RECT 11.065000  0.635000 11.370000 1.065000 ;
      RECT 11.255000  2.255000 11.635000 2.635000 ;
      RECT 11.560000  0.465000 11.735000 0.995000 ;
      RECT 11.560000  0.995000 12.235000 1.325000 ;
      RECT 11.560000  1.325000 11.730000 1.915000 ;
      RECT 11.905000  0.085000 12.325000 0.670000 ;
      RECT 11.905000  1.495000 12.330000 2.635000 ;
      RECT 12.995000  0.085000 13.165000 0.545000 ;
      RECT 12.995000  1.495000 13.245000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.855000  1.105000  1.025000 1.275000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.135000  1.785000  1.305000 1.955000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.480000  1.105000  5.650000 1.275000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.950000  1.785000  6.120000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.255000  0.765000  7.425000 0.935000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.615000  0.765000  7.785000 0.935000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.235000  1.105000  9.405000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.565000  1.785000  9.735000 1.955000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.140000  0.765000 11.310000 0.935000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
    LAYER met1 ;
      RECT 0.795000 1.075000 1.085000 1.120000 ;
      RECT 0.795000 1.120000 9.465000 1.260000 ;
      RECT 0.795000 1.260000 1.085000 1.305000 ;
      RECT 1.070000 1.755000 1.370000 1.800000 ;
      RECT 1.070000 1.800000 9.795000 1.940000 ;
      RECT 1.070000 1.940000 1.370000 1.985000 ;
      RECT 5.420000 1.075000 5.710000 1.120000 ;
      RECT 5.420000 1.260000 5.710000 1.305000 ;
      RECT 5.890000 1.755000 6.180000 1.800000 ;
      RECT 5.890000 1.940000 6.180000 1.985000 ;
      RECT 9.155000 1.075000 9.465000 1.120000 ;
      RECT 9.155000 1.260000 9.465000 1.305000 ;
      RECT 9.500000 1.755000 9.795000 1.800000 ;
      RECT 9.500000 1.940000 9.795000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrtp_2


MACRO sky130_fd_sc_hdll__sdfrtp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  12.88000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.160200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.120000 1.355000 3.655000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.513200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.420000 0.265000 12.785000 2.325000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.145000 0.735000  7.900000 0.780000 ;
        RECT  7.145000 0.780000 11.405000 0.920000 ;
        RECT  7.145000 0.920000  7.900000 0.965000 ;
        RECT 11.115000 0.735000 11.405000 0.780000 ;
        RECT 11.115000 0.920000 11.405000 0.965000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.172800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.610000 0.710000 4.955000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.467400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.070000 1.990000 1.335000 ;
        RECT 1.585000 1.335000 2.220000 1.745000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.880000 0.085000 ;
      RECT  0.000000  2.635000 12.880000 2.805000 ;
      RECT  0.090000  1.795000  0.915000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.885000 0.805000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.530000  2.135000  0.910000 2.635000 ;
      RECT  0.710000  0.805000  0.885000 0.995000 ;
      RECT  0.710000  0.995000  1.025000 1.325000 ;
      RECT  0.710000  1.325000  0.915000 1.795000 ;
      RECT  1.115000  0.345000  1.365000 0.675000 ;
      RECT  1.135000  1.730000  1.365000 2.465000 ;
      RECT  1.195000  0.675000  1.365000 1.730000 ;
      RECT  1.695000  0.395000  1.865000 0.730000 ;
      RECT  1.695000  0.730000  2.435000 0.900000 ;
      RECT  2.035000  0.085000  2.415000 0.560000 ;
      RECT  2.110000  1.915000  2.730000 2.085000 ;
      RECT  2.110000  2.085000  2.380000 2.400000 ;
      RECT  2.265000  0.900000  2.435000 0.995000 ;
      RECT  2.265000  0.995000  3.445000 1.165000 ;
      RECT  2.475000  1.165000  3.445000 1.185000 ;
      RECT  2.475000  1.185000  2.730000 1.915000 ;
      RECT  2.600000  2.255000  2.930000 2.635000 ;
      RECT  2.655000  0.085000  3.035000 0.825000 ;
      RECT  3.275000  0.255000  4.435000 0.425000 ;
      RECT  3.275000  0.425000  3.445000 0.995000 ;
      RECT  3.665000  0.675000  4.045000 1.075000 ;
      RECT  3.870000  1.075000  4.045000 1.935000 ;
      RECT  3.870000  1.935000  5.650000 2.105000 ;
      RECT  3.870000  2.105000  4.040000 2.465000 ;
      RECT  4.265000  0.425000  4.435000 1.685000 ;
      RECT  4.855000  2.275000  5.205000 2.635000 ;
      RECT  5.005000  0.085000  5.350000 0.540000 ;
      RECT  5.140000  0.715000  5.720000 0.895000 ;
      RECT  5.140000  0.895000  5.310000 1.935000 ;
      RECT  5.480000  1.065000  5.650000 1.395000 ;
      RECT  5.480000  2.105000  5.650000 2.185000 ;
      RECT  5.480000  2.185000  5.850000 2.435000 ;
      RECT  5.550000  0.335000  5.890000 0.505000 ;
      RECT  5.550000  0.505000  5.720000 0.715000 ;
      RECT  5.820000  1.575000  6.120000 1.955000 ;
      RECT  5.900000  0.705000  6.650000 1.035000 ;
      RECT  5.900000  1.035000  6.120000 1.575000 ;
      RECT  6.095000  2.135000  6.460000 2.465000 ;
      RECT  6.110000  0.305000  7.010000 0.475000 ;
      RECT  6.290000  1.215000  8.150000 1.385000 ;
      RECT  6.290000  1.385000  6.460000 2.135000 ;
      RECT  6.680000  1.935000  7.940000 2.105000 ;
      RECT  6.680000  2.105000  6.850000 2.375000 ;
      RECT  6.840000  0.475000  7.010000 1.215000 ;
      RECT  6.960000  1.595000  8.540000 1.765000 ;
      RECT  7.135000  2.355000  7.465000 2.635000 ;
      RECT  7.230000  0.765000  7.810000 1.045000 ;
      RECT  7.690000  0.085000  8.020000 0.545000 ;
      RECT  7.770000  2.105000  7.940000 2.375000 ;
      RECT  7.980000  1.005000  8.150000 1.215000 ;
      RECT  8.150000  2.175000  8.570000 2.635000 ;
      RECT  8.230000  0.275000  8.610000 0.445000 ;
      RECT  8.230000  0.445000  8.540000 0.835000 ;
      RECT  8.230000  1.765000  8.540000 1.835000 ;
      RECT  8.230000  1.835000  8.985000 2.005000 ;
      RECT  8.370000  0.835000  8.540000 1.595000 ;
      RECT  8.710000  0.705000  8.970000 1.495000 ;
      RECT  8.710000  1.495000  9.445000 1.660000 ;
      RECT  8.710000  1.660000  9.845000 1.665000 ;
      RECT  8.780000  0.255000  9.890000 0.535000 ;
      RECT  8.815000  2.005000  8.985000 2.465000 ;
      RECT  9.185000  1.665000  9.845000 1.955000 ;
      RECT  9.195000  2.125000 10.215000 2.465000 ;
      RECT  9.235000  0.920000  9.405000 1.325000 ;
      RECT  9.670000  0.535000  9.890000 1.315000 ;
      RECT  9.670000  1.315000 10.285000 1.485000 ;
      RECT 10.040000  1.485000 10.285000 1.575000 ;
      RECT 10.040000  1.575000 11.370000 1.745000 ;
      RECT 10.040000  1.745000 10.215000 2.125000 ;
      RECT 10.110000  0.085000 10.330000 0.525000 ;
      RECT 10.150000  0.695000 10.730000 0.865000 ;
      RECT 10.150000  0.865000 10.370000 1.145000 ;
      RECT 10.415000  2.195000 10.665000 2.635000 ;
      RECT 10.560000  0.295000 11.735000 0.465000 ;
      RECT 10.560000  0.465000 10.730000 0.695000 ;
      RECT 10.600000  1.065000 11.370000 1.275000 ;
      RECT 10.910000  1.915000 11.730000 2.085000 ;
      RECT 10.910000  2.085000 11.080000 2.375000 ;
      RECT 11.065000  0.635000 11.370000 1.065000 ;
      RECT 11.255000  2.255000 11.635000 2.635000 ;
      RECT 11.560000  0.465000 11.735000 0.995000 ;
      RECT 11.560000  0.995000 12.205000 1.325000 ;
      RECT 11.560000  1.325000 11.730000 1.915000 ;
      RECT 11.905000  0.085000 12.190000 0.710000 ;
      RECT 11.905000  1.495000 12.190000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.855000  1.105000  1.025000 1.275000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.135000  1.785000  1.305000 1.955000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.480000  1.105000  5.650000 1.275000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.950000  1.785000  6.120000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.255000  0.765000  7.425000 0.935000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.615000  0.765000  7.785000 0.935000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.235000  1.105000  9.405000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.565000  1.785000  9.735000 1.955000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.175000  0.765000 11.345000 0.935000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
    LAYER met1 ;
      RECT 0.795000 1.075000 1.085000 1.120000 ;
      RECT 0.795000 1.120000 9.465000 1.260000 ;
      RECT 0.795000 1.260000 1.085000 1.305000 ;
      RECT 1.070000 1.755000 1.370000 1.800000 ;
      RECT 1.070000 1.800000 9.795000 1.940000 ;
      RECT 1.070000 1.940000 1.370000 1.985000 ;
      RECT 5.420000 1.075000 5.710000 1.120000 ;
      RECT 5.420000 1.260000 5.710000 1.305000 ;
      RECT 5.890000 1.755000 6.180000 1.800000 ;
      RECT 5.890000 1.940000 6.180000 1.985000 ;
      RECT 9.155000 1.075000 9.465000 1.120000 ;
      RECT 9.155000 1.260000 9.465000 1.305000 ;
      RECT 9.500000 1.755000 9.795000 1.800000 ;
      RECT 9.500000 1.940000 9.795000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrtp_1


MACRO sky130_fd_sc_hdll__a22oi_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.645000 1.075000 3.535000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.770000 1.075000 4.620000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 1.075000 1.745000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 1.075000 0.830000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.278500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.485000 2.360000 1.655000 ;
        RECT 0.095000 1.655000 0.345000 2.465000 ;
        RECT 0.985000 1.655000 1.365000 2.125000 ;
        RECT 1.455000 0.675000 3.295000 0.845000 ;
        RECT 1.925000 1.655000 2.360000 2.125000 ;
        RECT 1.930000 0.845000 2.360000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.060000 0.085000 ;
        RECT 0.515000  0.085000 0.895000 0.510000 ;
        RECT 3.980000  0.085000 4.360000 0.510000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.060000 2.805000 ;
        RECT 3.045000 1.825000 3.215000 2.635000 ;
        RECT 4.085000 1.825000 4.255000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.255000 0.345000 0.680000 ;
      RECT 0.095000 0.680000 1.285000 0.850000 ;
      RECT 0.515000 1.825000 0.815000 2.295000 ;
      RECT 0.515000 2.295000 2.825000 2.465000 ;
      RECT 1.115000 0.255000 2.305000 0.505000 ;
      RECT 1.115000 0.505000 1.285000 0.680000 ;
      RECT 1.585000 1.825000 1.755000 2.295000 ;
      RECT 2.495000 0.255000 3.785000 0.505000 ;
      RECT 2.575000 1.485000 4.805000 1.655000 ;
      RECT 2.575000 1.655000 2.825000 2.295000 ;
      RECT 3.385000 1.655000 3.865000 2.465000 ;
      RECT 3.615000 0.505000 3.785000 0.680000 ;
      RECT 3.615000 0.680000 4.875000 0.850000 ;
      RECT 4.425000 1.655000 4.805000 2.465000 ;
      RECT 4.555000 0.255000 4.875000 0.680000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22oi_2


MACRO sky130_fd_sc_hdll__a22oi_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.675000 1.735000 1.055000 ;
        RECT 1.525000 1.055000 2.085000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265000 0.995000 2.625000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.815000 1.075000 1.315000 1.275000 ;
        RECT 1.065000 0.675000 1.315000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.765000 0.625000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.917000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.445000 3.135000 1.615000 ;
        RECT 0.095000 1.615000 0.425000 2.295000 ;
        RECT 0.095000 2.295000 1.375000 2.465000 ;
        RECT 0.870000 0.255000 2.275000 0.505000 ;
        RECT 1.035000 2.195000 1.375000 2.295000 ;
        RECT 2.095000 0.505000 2.275000 0.655000 ;
        RECT 2.095000 0.655000 3.135000 0.825000 ;
        RECT 2.795000 0.825000 3.135000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.095000  0.085000 0.595000 0.595000 ;
      RECT 0.645000  1.785000 2.275000 1.980000 ;
      RECT 0.645000  1.980000 0.815000 2.115000 ;
      RECT 1.555000  2.255000 1.910000 2.635000 ;
      RECT 2.105000  1.980000 2.275000 2.165000 ;
      RECT 2.505000  0.085000 2.835000 0.485000 ;
      RECT 2.560000  1.855000 2.825000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22oi_1


MACRO sky130_fd_sc_hdll__a22oi_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.740000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675000 1.075000 6.285000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.510000 1.075000 8.535000 1.285000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 1.075000 4.440000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 2.095000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.645000 1.445000 3.675000 1.625000 ;
        RECT 0.645000 1.625000 0.855000 2.125000 ;
        RECT 1.545000 1.625000 1.795000 2.125000 ;
        RECT 2.395000 0.645000 6.115000 0.885000 ;
        RECT 2.395000 0.885000 2.695000 1.445000 ;
        RECT 2.485000 1.625000 2.735000 2.125000 ;
        RECT 3.425000 1.625000 3.675000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.090000  1.455000 0.425000 2.295000 ;
      RECT 0.090000  2.295000 4.665000 2.465000 ;
      RECT 0.095000  0.255000 0.425000 0.725000 ;
      RECT 0.095000  0.725000 2.225000 0.905000 ;
      RECT 0.645000  0.085000 0.815000 0.555000 ;
      RECT 0.985000  0.255000 1.365000 0.725000 ;
      RECT 1.075000  1.795000 1.325000 2.295000 ;
      RECT 1.585000  0.085000 1.755000 0.555000 ;
      RECT 1.925000  0.255000 4.185000 0.475000 ;
      RECT 1.925000  0.475000 2.225000 0.725000 ;
      RECT 2.015000  1.795000 2.265000 2.295000 ;
      RECT 2.955000  1.795000 3.205000 2.295000 ;
      RECT 3.895000  1.455000 8.425000 1.625000 ;
      RECT 3.895000  1.625000 4.665000 2.295000 ;
      RECT 4.375000  0.255000 6.585000 0.475000 ;
      RECT 4.885000  1.795000 5.135000 2.635000 ;
      RECT 5.355000  1.625000 5.605000 2.465000 ;
      RECT 5.825000  1.795000 6.075000 2.635000 ;
      RECT 6.295000  1.625000 6.545000 2.465000 ;
      RECT 6.335000  0.475000 6.585000 0.725000 ;
      RECT 6.335000  0.725000 8.465000 0.905000 ;
      RECT 6.765000  1.795000 7.015000 2.635000 ;
      RECT 6.805000  0.085000 6.975000 0.555000 ;
      RECT 7.145000  0.255000 7.525000 0.725000 ;
      RECT 7.235000  1.625000 7.485000 2.465000 ;
      RECT 7.705000  1.795000 7.955000 2.635000 ;
      RECT 7.745000  0.085000 7.915000 0.555000 ;
      RECT 8.085000  0.255000 8.465000 0.725000 ;
      RECT 8.175000  1.625000 8.425000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22oi_4


MACRO sky130_fd_sc_hdll__muxb16to1_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  25.76000 BY  5.440000 ;
  SITE unithd ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.055000 0.915000 1.325000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.525000 1.055000 6.345000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 1.055000 7.355000 1.325000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.965000 1.055000 12.785000 1.325000 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.975000 1.055000 13.795000 1.325000 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.405000 1.055000 19.225000 1.325000 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.415000 1.055000 20.235000 1.325000 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.845000 1.055000 25.665000 1.325000 ;
    END
  END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 4.115000 0.915000 4.385000 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.525000 4.115000 6.345000 4.385000 ;
    END
  END D[9]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 4.115000 7.355000 4.385000 ;
    END
  END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.965000 4.115000 12.785000 4.385000 ;
    END
  END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.975000 4.115000 13.795000 4.385000 ;
    END
  END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.405000 4.115000 19.225000 4.385000 ;
    END
  END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.415000 4.115000 20.235000 4.385000 ;
    END
  END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.845000 4.115000 25.665000 4.385000 ;
    END
  END D[15]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 1.025000 3.125000 1.295000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.025000 3.650000 1.295000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.230000 1.025000 9.565000 1.295000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.755000 1.025000 10.090000 1.295000 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.670000 1.025000 16.005000 1.295000 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.195000 1.025000 16.530000 1.295000 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.110000 1.025000 22.445000 1.295000 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.635000 1.025000 22.970000 1.295000 ;
    END
  END S[7]
  PIN S[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 4.145000 3.125000 4.415000 ;
    END
  END S[8]
  PIN S[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 4.145000 3.650000 4.415000 ;
    END
  END S[9]
  PIN S[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.230000 4.145000 9.565000 4.415000 ;
    END
  END S[10]
  PIN S[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.755000 4.145000 10.090000 4.415000 ;
    END
  END S[11]
  PIN S[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.670000 4.145000 16.005000 4.415000 ;
    END
  END S[12]
  PIN S[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.195000 4.145000 16.530000 4.415000 ;
    END
  END S[13]
  PIN S[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.110000 4.145000 22.445000 4.415000 ;
    END
  END S[14]
  PIN S[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.635000 4.145000 22.970000 4.415000 ;
    END
  END S[15]
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  1.465000 1.755000  1.755000 1.800000 ;
        RECT  1.465000 1.800000 24.295000 1.940000 ;
        RECT  1.465000 1.940000  1.755000 1.985000 ;
        RECT  1.465000 3.455000  1.755000 3.500000 ;
        RECT  1.465000 3.500000 24.295000 3.640000 ;
        RECT  1.465000 3.640000  1.755000 3.685000 ;
        RECT  4.685000 1.755000  4.975000 1.800000 ;
        RECT  4.685000 1.940000  4.975000 1.985000 ;
        RECT  4.685000 3.455000  4.975000 3.500000 ;
        RECT  4.685000 3.640000  4.975000 3.685000 ;
        RECT  7.905000 1.755000  8.195000 1.800000 ;
        RECT  7.905000 1.940000  8.195000 1.985000 ;
        RECT  7.905000 3.455000  8.195000 3.500000 ;
        RECT  7.905000 3.640000  8.195000 3.685000 ;
        RECT 11.125000 1.755000 11.415000 1.800000 ;
        RECT 11.125000 1.940000 11.415000 1.985000 ;
        RECT 11.125000 3.455000 11.415000 3.500000 ;
        RECT 11.125000 3.640000 11.415000 3.685000 ;
        RECT 14.345000 1.755000 14.635000 1.800000 ;
        RECT 14.345000 1.940000 14.635000 1.985000 ;
        RECT 14.345000 3.455000 14.635000 3.500000 ;
        RECT 14.345000 3.640000 14.635000 3.685000 ;
        RECT 17.565000 1.755000 17.855000 1.800000 ;
        RECT 17.565000 1.940000 17.855000 1.985000 ;
        RECT 17.565000 3.455000 17.855000 3.500000 ;
        RECT 17.565000 3.640000 17.855000 3.685000 ;
        RECT 20.785000 1.755000 21.075000 1.800000 ;
        RECT 20.785000 1.940000 21.075000 1.985000 ;
        RECT 20.785000 3.455000 21.075000 3.500000 ;
        RECT 20.785000 3.640000 21.075000 3.685000 ;
        RECT 24.005000 1.755000 24.295000 1.800000 ;
        RECT 24.005000 1.940000 24.295000 1.985000 ;
        RECT 24.005000 3.455000 24.295000 3.500000 ;
        RECT 24.005000 3.640000 24.295000 3.685000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 25.760000 0.240000 ;
        RECT 0.000000  5.200000 25.760000 5.680000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 25.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 25.760000 0.085000 ;
      RECT  0.000000  2.635000  1.415000 2.805000 ;
      RECT  0.000000  5.355000 25.760000 5.525000 ;
      RECT  0.095000  1.495000  1.285000 1.665000 ;
      RECT  0.095000  1.665000  0.395000 2.210000 ;
      RECT  0.095000  2.210000  0.425000 2.465000 ;
      RECT  0.095000  2.975000  0.425000 3.230000 ;
      RECT  0.095000  3.230000  0.395000 3.775000 ;
      RECT  0.095000  3.775000  1.285000 3.945000 ;
      RECT  0.145000  0.255000  0.475000 0.715000 ;
      RECT  0.145000  0.715000  1.335000 0.885000 ;
      RECT  0.145000  4.555000  1.335000 4.725000 ;
      RECT  0.145000  4.725000  0.475000 5.185000 ;
      RECT  0.565000  1.835000  0.895000 2.105000 ;
      RECT  0.565000  3.335000  0.895000 3.605000 ;
      RECT  0.595000  2.105000  0.895000 2.635000 ;
      RECT  0.595000  2.805000  0.895000 3.335000 ;
      RECT  0.645000  0.085000  0.860000 0.545000 ;
      RECT  0.645000  4.895000  0.860000 5.355000 ;
      RECT  1.030000  0.255000  2.175000 0.425000 ;
      RECT  1.030000  0.425000  1.335000 0.715000 ;
      RECT  1.030000  0.885000  1.335000 0.925000 ;
      RECT  1.030000  4.515000  1.335000 4.555000 ;
      RECT  1.030000  4.725000  1.335000 5.015000 ;
      RECT  1.030000  5.015000  2.175000 5.185000 ;
      RECT  1.115000  1.665000  1.285000 2.295000 ;
      RECT  1.115000  2.295000  1.415000 2.465000 ;
      RECT  1.115000  2.975000  1.415000 3.145000 ;
      RECT  1.115000  3.145000  1.285000 3.775000 ;
      RECT  1.465000  1.755000  1.895000 2.125000 ;
      RECT  1.465000  3.315000  1.895000 3.685000 ;
      RECT  1.505000  0.595000  1.835000 0.885000 ;
      RECT  1.505000  4.555000  1.835000 4.845000 ;
      RECT  1.585000  0.885000  1.755000 1.755000 ;
      RECT  1.585000  2.125000  1.755000 3.315000 ;
      RECT  1.585000  3.685000  1.755000 4.555000 ;
      RECT  1.925000  2.295000  2.280000 2.465000 ;
      RECT  1.925000  2.635000  4.515000 2.805000 ;
      RECT  1.925000  2.975000  2.280000 3.145000 ;
      RECT  2.005000  0.425000  2.175000 0.770000 ;
      RECT  2.005000  4.670000  2.175000 5.015000 ;
      RECT  2.100000  1.205000  2.515000 1.305000 ;
      RECT  2.100000  1.305000  2.620000 1.465000 ;
      RECT  2.100000  1.465000  2.880000 1.475000 ;
      RECT  2.100000  3.965000  2.880000 3.975000 ;
      RECT  2.100000  3.975000  2.620000 4.135000 ;
      RECT  2.100000  4.135000  2.515000 4.235000 ;
      RECT  2.110000  1.645000  2.280000 2.295000 ;
      RECT  2.110000  3.145000  2.280000 3.795000 ;
      RECT  2.345000  0.585000  2.925000 0.755000 ;
      RECT  2.345000  0.755000  2.515000 1.205000 ;
      RECT  2.345000  4.235000  2.515000 4.685000 ;
      RECT  2.345000  4.685000  2.925000 4.855000 ;
      RECT  2.450000  1.475000  2.880000 1.635000 ;
      RECT  2.450000  3.805000  2.880000 3.965000 ;
      RECT  2.550000  1.635000  2.880000 2.465000 ;
      RECT  2.550000  2.975000  2.880000 3.805000 ;
      RECT  2.675000  0.330000  2.925000 0.585000 ;
      RECT  2.675000  4.855000  2.925000 5.110000 ;
      RECT  3.055000  1.465000  3.385000 2.635000 ;
      RECT  3.055000  2.805000  3.385000 3.975000 ;
      RECT  3.095000  0.085000  3.345000 0.660000 ;
      RECT  3.095000  4.780000  3.345000 5.355000 ;
      RECT  3.515000  0.330000  3.765000 0.585000 ;
      RECT  3.515000  0.585000  4.095000 0.755000 ;
      RECT  3.515000  4.685000  4.095000 4.855000 ;
      RECT  3.515000  4.855000  3.765000 5.110000 ;
      RECT  3.560000  1.465000  4.340000 1.475000 ;
      RECT  3.560000  1.475000  3.990000 1.635000 ;
      RECT  3.560000  1.635000  3.890000 2.465000 ;
      RECT  3.560000  2.975000  3.890000 3.805000 ;
      RECT  3.560000  3.805000  3.990000 3.965000 ;
      RECT  3.560000  3.965000  4.340000 3.975000 ;
      RECT  3.820000  1.305000  4.340000 1.465000 ;
      RECT  3.820000  3.975000  4.340000 4.135000 ;
      RECT  3.925000  0.755000  4.095000 1.205000 ;
      RECT  3.925000  1.205000  4.340000 1.305000 ;
      RECT  3.925000  4.135000  4.340000 4.235000 ;
      RECT  3.925000  4.235000  4.095000 4.685000 ;
      RECT  4.160000  1.645000  4.330000 2.295000 ;
      RECT  4.160000  2.295000  4.515000 2.465000 ;
      RECT  4.160000  2.975000  4.515000 3.145000 ;
      RECT  4.160000  3.145000  4.330000 3.795000 ;
      RECT  4.265000  0.255000  5.410000 0.425000 ;
      RECT  4.265000  0.425000  4.435000 0.770000 ;
      RECT  4.265000  4.670000  4.435000 5.015000 ;
      RECT  4.265000  5.015000  5.410000 5.185000 ;
      RECT  4.545000  1.755000  4.975000 2.125000 ;
      RECT  4.545000  3.315000  4.975000 3.685000 ;
      RECT  4.605000  0.595000  4.935000 0.885000 ;
      RECT  4.605000  4.555000  4.935000 4.845000 ;
      RECT  4.685000  0.885000  4.855000 1.755000 ;
      RECT  4.685000  2.125000  4.855000 3.315000 ;
      RECT  4.685000  3.685000  4.855000 4.555000 ;
      RECT  5.025000  2.295000  5.325000 2.465000 ;
      RECT  5.025000  2.635000  7.855000 2.805000 ;
      RECT  5.025000  2.975000  5.325000 3.145000 ;
      RECT  5.105000  0.425000  5.410000 0.715000 ;
      RECT  5.105000  0.715000  6.295000 0.885000 ;
      RECT  5.105000  0.885000  5.410000 0.925000 ;
      RECT  5.105000  4.515000  5.410000 4.555000 ;
      RECT  5.105000  4.555000  6.295000 4.725000 ;
      RECT  5.105000  4.725000  5.410000 5.015000 ;
      RECT  5.155000  1.495000  6.345000 1.665000 ;
      RECT  5.155000  1.665000  5.325000 2.295000 ;
      RECT  5.155000  3.145000  5.325000 3.775000 ;
      RECT  5.155000  3.775000  6.345000 3.945000 ;
      RECT  5.545000  1.835000  5.875000 2.105000 ;
      RECT  5.545000  2.105000  5.845000 2.635000 ;
      RECT  5.545000  2.805000  5.845000 3.335000 ;
      RECT  5.545000  3.335000  5.875000 3.605000 ;
      RECT  5.580000  0.085000  5.795000 0.545000 ;
      RECT  5.580000  4.895000  5.795000 5.355000 ;
      RECT  5.965000  0.255000  6.295000 0.715000 ;
      RECT  5.965000  4.725000  6.295000 5.185000 ;
      RECT  6.015000  2.210000  6.345000 2.465000 ;
      RECT  6.015000  2.975000  6.345000 3.230000 ;
      RECT  6.045000  1.665000  6.345000 2.210000 ;
      RECT  6.045000  3.230000  6.345000 3.775000 ;
      RECT  6.535000  1.495000  7.725000 1.665000 ;
      RECT  6.535000  1.665000  6.835000 2.210000 ;
      RECT  6.535000  2.210000  6.865000 2.465000 ;
      RECT  6.535000  2.975000  6.865000 3.230000 ;
      RECT  6.535000  3.230000  6.835000 3.775000 ;
      RECT  6.535000  3.775000  7.725000 3.945000 ;
      RECT  6.585000  0.255000  6.915000 0.715000 ;
      RECT  6.585000  0.715000  7.775000 0.885000 ;
      RECT  6.585000  4.555000  7.775000 4.725000 ;
      RECT  6.585000  4.725000  6.915000 5.185000 ;
      RECT  7.005000  1.835000  7.335000 2.105000 ;
      RECT  7.005000  3.335000  7.335000 3.605000 ;
      RECT  7.035000  2.105000  7.335000 2.635000 ;
      RECT  7.035000  2.805000  7.335000 3.335000 ;
      RECT  7.085000  0.085000  7.300000 0.545000 ;
      RECT  7.085000  4.895000  7.300000 5.355000 ;
      RECT  7.470000  0.255000  8.615000 0.425000 ;
      RECT  7.470000  0.425000  7.775000 0.715000 ;
      RECT  7.470000  0.885000  7.775000 0.925000 ;
      RECT  7.470000  4.515000  7.775000 4.555000 ;
      RECT  7.470000  4.725000  7.775000 5.015000 ;
      RECT  7.470000  5.015000  8.615000 5.185000 ;
      RECT  7.555000  1.665000  7.725000 2.295000 ;
      RECT  7.555000  2.295000  7.855000 2.465000 ;
      RECT  7.555000  2.975000  7.855000 3.145000 ;
      RECT  7.555000  3.145000  7.725000 3.775000 ;
      RECT  7.905000  1.755000  8.335000 2.125000 ;
      RECT  7.905000  3.315000  8.335000 3.685000 ;
      RECT  7.945000  0.595000  8.275000 0.885000 ;
      RECT  7.945000  4.555000  8.275000 4.845000 ;
      RECT  8.025000  0.885000  8.195000 1.755000 ;
      RECT  8.025000  2.125000  8.195000 3.315000 ;
      RECT  8.025000  3.685000  8.195000 4.555000 ;
      RECT  8.365000  2.295000  8.720000 2.465000 ;
      RECT  8.365000  2.635000 10.955000 2.805000 ;
      RECT  8.365000  2.975000  8.720000 3.145000 ;
      RECT  8.445000  0.425000  8.615000 0.770000 ;
      RECT  8.445000  4.670000  8.615000 5.015000 ;
      RECT  8.540000  1.205000  8.955000 1.305000 ;
      RECT  8.540000  1.305000  9.060000 1.465000 ;
      RECT  8.540000  1.465000  9.320000 1.475000 ;
      RECT  8.540000  3.965000  9.320000 3.975000 ;
      RECT  8.540000  3.975000  9.060000 4.135000 ;
      RECT  8.540000  4.135000  8.955000 4.235000 ;
      RECT  8.550000  1.645000  8.720000 2.295000 ;
      RECT  8.550000  3.145000  8.720000 3.795000 ;
      RECT  8.785000  0.585000  9.365000 0.755000 ;
      RECT  8.785000  0.755000  8.955000 1.205000 ;
      RECT  8.785000  4.235000  8.955000 4.685000 ;
      RECT  8.785000  4.685000  9.365000 4.855000 ;
      RECT  8.890000  1.475000  9.320000 1.635000 ;
      RECT  8.890000  3.805000  9.320000 3.965000 ;
      RECT  8.990000  1.635000  9.320000 2.465000 ;
      RECT  8.990000  2.975000  9.320000 3.805000 ;
      RECT  9.115000  0.330000  9.365000 0.585000 ;
      RECT  9.115000  4.855000  9.365000 5.110000 ;
      RECT  9.495000  1.465000  9.825000 2.635000 ;
      RECT  9.495000  2.805000  9.825000 3.975000 ;
      RECT  9.535000  0.085000  9.785000 0.660000 ;
      RECT  9.535000  4.780000  9.785000 5.355000 ;
      RECT  9.955000  0.330000 10.205000 0.585000 ;
      RECT  9.955000  0.585000 10.535000 0.755000 ;
      RECT  9.955000  4.685000 10.535000 4.855000 ;
      RECT  9.955000  4.855000 10.205000 5.110000 ;
      RECT 10.000000  1.465000 10.780000 1.475000 ;
      RECT 10.000000  1.475000 10.430000 1.635000 ;
      RECT 10.000000  1.635000 10.330000 2.465000 ;
      RECT 10.000000  2.975000 10.330000 3.805000 ;
      RECT 10.000000  3.805000 10.430000 3.965000 ;
      RECT 10.000000  3.965000 10.780000 3.975000 ;
      RECT 10.260000  1.305000 10.780000 1.465000 ;
      RECT 10.260000  3.975000 10.780000 4.135000 ;
      RECT 10.365000  0.755000 10.535000 1.205000 ;
      RECT 10.365000  1.205000 10.780000 1.305000 ;
      RECT 10.365000  4.135000 10.780000 4.235000 ;
      RECT 10.365000  4.235000 10.535000 4.685000 ;
      RECT 10.600000  1.645000 10.770000 2.295000 ;
      RECT 10.600000  2.295000 10.955000 2.465000 ;
      RECT 10.600000  2.975000 10.955000 3.145000 ;
      RECT 10.600000  3.145000 10.770000 3.795000 ;
      RECT 10.705000  0.255000 11.850000 0.425000 ;
      RECT 10.705000  0.425000 10.875000 0.770000 ;
      RECT 10.705000  4.670000 10.875000 5.015000 ;
      RECT 10.705000  5.015000 11.850000 5.185000 ;
      RECT 10.985000  1.755000 11.415000 2.125000 ;
      RECT 10.985000  3.315000 11.415000 3.685000 ;
      RECT 11.045000  0.595000 11.375000 0.885000 ;
      RECT 11.045000  4.555000 11.375000 4.845000 ;
      RECT 11.125000  0.885000 11.295000 1.755000 ;
      RECT 11.125000  2.125000 11.295000 3.315000 ;
      RECT 11.125000  3.685000 11.295000 4.555000 ;
      RECT 11.465000  2.295000 11.765000 2.465000 ;
      RECT 11.465000  2.635000 14.295000 2.805000 ;
      RECT 11.465000  2.975000 11.765000 3.145000 ;
      RECT 11.545000  0.425000 11.850000 0.715000 ;
      RECT 11.545000  0.715000 12.735000 0.885000 ;
      RECT 11.545000  0.885000 11.850000 0.925000 ;
      RECT 11.545000  4.515000 11.850000 4.555000 ;
      RECT 11.545000  4.555000 12.735000 4.725000 ;
      RECT 11.545000  4.725000 11.850000 5.015000 ;
      RECT 11.595000  1.495000 12.785000 1.665000 ;
      RECT 11.595000  1.665000 11.765000 2.295000 ;
      RECT 11.595000  3.145000 11.765000 3.775000 ;
      RECT 11.595000  3.775000 12.785000 3.945000 ;
      RECT 11.985000  1.835000 12.315000 2.105000 ;
      RECT 11.985000  2.105000 12.285000 2.635000 ;
      RECT 11.985000  2.805000 12.285000 3.335000 ;
      RECT 11.985000  3.335000 12.315000 3.605000 ;
      RECT 12.020000  0.085000 12.235000 0.545000 ;
      RECT 12.020000  4.895000 12.235000 5.355000 ;
      RECT 12.405000  0.255000 12.735000 0.715000 ;
      RECT 12.405000  4.725000 12.735000 5.185000 ;
      RECT 12.455000  2.210000 12.785000 2.465000 ;
      RECT 12.455000  2.975000 12.785000 3.230000 ;
      RECT 12.485000  1.665000 12.785000 2.210000 ;
      RECT 12.485000  3.230000 12.785000 3.775000 ;
      RECT 12.975000  1.495000 14.165000 1.665000 ;
      RECT 12.975000  1.665000 13.275000 2.210000 ;
      RECT 12.975000  2.210000 13.305000 2.465000 ;
      RECT 12.975000  2.975000 13.305000 3.230000 ;
      RECT 12.975000  3.230000 13.275000 3.775000 ;
      RECT 12.975000  3.775000 14.165000 3.945000 ;
      RECT 13.025000  0.255000 13.355000 0.715000 ;
      RECT 13.025000  0.715000 14.215000 0.885000 ;
      RECT 13.025000  4.555000 14.215000 4.725000 ;
      RECT 13.025000  4.725000 13.355000 5.185000 ;
      RECT 13.445000  1.835000 13.775000 2.105000 ;
      RECT 13.445000  3.335000 13.775000 3.605000 ;
      RECT 13.475000  2.105000 13.775000 2.635000 ;
      RECT 13.475000  2.805000 13.775000 3.335000 ;
      RECT 13.525000  0.085000 13.740000 0.545000 ;
      RECT 13.525000  4.895000 13.740000 5.355000 ;
      RECT 13.910000  0.255000 15.055000 0.425000 ;
      RECT 13.910000  0.425000 14.215000 0.715000 ;
      RECT 13.910000  0.885000 14.215000 0.925000 ;
      RECT 13.910000  4.515000 14.215000 4.555000 ;
      RECT 13.910000  4.725000 14.215000 5.015000 ;
      RECT 13.910000  5.015000 15.055000 5.185000 ;
      RECT 13.995000  1.665000 14.165000 2.295000 ;
      RECT 13.995000  2.295000 14.295000 2.465000 ;
      RECT 13.995000  2.975000 14.295000 3.145000 ;
      RECT 13.995000  3.145000 14.165000 3.775000 ;
      RECT 14.345000  1.755000 14.775000 2.125000 ;
      RECT 14.345000  3.315000 14.775000 3.685000 ;
      RECT 14.385000  0.595000 14.715000 0.885000 ;
      RECT 14.385000  4.555000 14.715000 4.845000 ;
      RECT 14.465000  0.885000 14.635000 1.755000 ;
      RECT 14.465000  2.125000 14.635000 3.315000 ;
      RECT 14.465000  3.685000 14.635000 4.555000 ;
      RECT 14.805000  2.295000 15.160000 2.465000 ;
      RECT 14.805000  2.635000 17.395000 2.805000 ;
      RECT 14.805000  2.975000 15.160000 3.145000 ;
      RECT 14.885000  0.425000 15.055000 0.770000 ;
      RECT 14.885000  4.670000 15.055000 5.015000 ;
      RECT 14.980000  1.205000 15.395000 1.305000 ;
      RECT 14.980000  1.305000 15.500000 1.465000 ;
      RECT 14.980000  1.465000 15.760000 1.475000 ;
      RECT 14.980000  3.965000 15.760000 3.975000 ;
      RECT 14.980000  3.975000 15.500000 4.135000 ;
      RECT 14.980000  4.135000 15.395000 4.235000 ;
      RECT 14.990000  1.645000 15.160000 2.295000 ;
      RECT 14.990000  3.145000 15.160000 3.795000 ;
      RECT 15.225000  0.585000 15.805000 0.755000 ;
      RECT 15.225000  0.755000 15.395000 1.205000 ;
      RECT 15.225000  4.235000 15.395000 4.685000 ;
      RECT 15.225000  4.685000 15.805000 4.855000 ;
      RECT 15.330000  1.475000 15.760000 1.635000 ;
      RECT 15.330000  3.805000 15.760000 3.965000 ;
      RECT 15.430000  1.635000 15.760000 2.465000 ;
      RECT 15.430000  2.975000 15.760000 3.805000 ;
      RECT 15.555000  0.330000 15.805000 0.585000 ;
      RECT 15.555000  4.855000 15.805000 5.110000 ;
      RECT 15.935000  1.465000 16.265000 2.635000 ;
      RECT 15.935000  2.805000 16.265000 3.975000 ;
      RECT 15.975000  0.085000 16.225000 0.660000 ;
      RECT 15.975000  4.780000 16.225000 5.355000 ;
      RECT 16.395000  0.330000 16.645000 0.585000 ;
      RECT 16.395000  0.585000 16.975000 0.755000 ;
      RECT 16.395000  4.685000 16.975000 4.855000 ;
      RECT 16.395000  4.855000 16.645000 5.110000 ;
      RECT 16.440000  1.465000 17.220000 1.475000 ;
      RECT 16.440000  1.475000 16.870000 1.635000 ;
      RECT 16.440000  1.635000 16.770000 2.465000 ;
      RECT 16.440000  2.975000 16.770000 3.805000 ;
      RECT 16.440000  3.805000 16.870000 3.965000 ;
      RECT 16.440000  3.965000 17.220000 3.975000 ;
      RECT 16.700000  1.305000 17.220000 1.465000 ;
      RECT 16.700000  3.975000 17.220000 4.135000 ;
      RECT 16.805000  0.755000 16.975000 1.205000 ;
      RECT 16.805000  1.205000 17.220000 1.305000 ;
      RECT 16.805000  4.135000 17.220000 4.235000 ;
      RECT 16.805000  4.235000 16.975000 4.685000 ;
      RECT 17.040000  1.645000 17.210000 2.295000 ;
      RECT 17.040000  2.295000 17.395000 2.465000 ;
      RECT 17.040000  2.975000 17.395000 3.145000 ;
      RECT 17.040000  3.145000 17.210000 3.795000 ;
      RECT 17.145000  0.255000 18.290000 0.425000 ;
      RECT 17.145000  0.425000 17.315000 0.770000 ;
      RECT 17.145000  4.670000 17.315000 5.015000 ;
      RECT 17.145000  5.015000 18.290000 5.185000 ;
      RECT 17.425000  1.755000 17.855000 2.125000 ;
      RECT 17.425000  3.315000 17.855000 3.685000 ;
      RECT 17.485000  0.595000 17.815000 0.885000 ;
      RECT 17.485000  4.555000 17.815000 4.845000 ;
      RECT 17.565000  0.885000 17.735000 1.755000 ;
      RECT 17.565000  2.125000 17.735000 3.315000 ;
      RECT 17.565000  3.685000 17.735000 4.555000 ;
      RECT 17.905000  2.295000 18.205000 2.465000 ;
      RECT 17.905000  2.635000 20.735000 2.805000 ;
      RECT 17.905000  2.975000 18.205000 3.145000 ;
      RECT 17.985000  0.425000 18.290000 0.715000 ;
      RECT 17.985000  0.715000 19.175000 0.885000 ;
      RECT 17.985000  0.885000 18.290000 0.925000 ;
      RECT 17.985000  4.515000 18.290000 4.555000 ;
      RECT 17.985000  4.555000 19.175000 4.725000 ;
      RECT 17.985000  4.725000 18.290000 5.015000 ;
      RECT 18.035000  1.495000 19.225000 1.665000 ;
      RECT 18.035000  1.665000 18.205000 2.295000 ;
      RECT 18.035000  3.145000 18.205000 3.775000 ;
      RECT 18.035000  3.775000 19.225000 3.945000 ;
      RECT 18.425000  1.835000 18.755000 2.105000 ;
      RECT 18.425000  2.105000 18.725000 2.635000 ;
      RECT 18.425000  2.805000 18.725000 3.335000 ;
      RECT 18.425000  3.335000 18.755000 3.605000 ;
      RECT 18.460000  0.085000 18.675000 0.545000 ;
      RECT 18.460000  4.895000 18.675000 5.355000 ;
      RECT 18.845000  0.255000 19.175000 0.715000 ;
      RECT 18.845000  4.725000 19.175000 5.185000 ;
      RECT 18.895000  2.210000 19.225000 2.465000 ;
      RECT 18.895000  2.975000 19.225000 3.230000 ;
      RECT 18.925000  1.665000 19.225000 2.210000 ;
      RECT 18.925000  3.230000 19.225000 3.775000 ;
      RECT 19.415000  1.495000 20.605000 1.665000 ;
      RECT 19.415000  1.665000 19.715000 2.210000 ;
      RECT 19.415000  2.210000 19.745000 2.465000 ;
      RECT 19.415000  2.975000 19.745000 3.230000 ;
      RECT 19.415000  3.230000 19.715000 3.775000 ;
      RECT 19.415000  3.775000 20.605000 3.945000 ;
      RECT 19.465000  0.255000 19.795000 0.715000 ;
      RECT 19.465000  0.715000 20.655000 0.885000 ;
      RECT 19.465000  4.555000 20.655000 4.725000 ;
      RECT 19.465000  4.725000 19.795000 5.185000 ;
      RECT 19.885000  1.835000 20.215000 2.105000 ;
      RECT 19.885000  3.335000 20.215000 3.605000 ;
      RECT 19.915000  2.105000 20.215000 2.635000 ;
      RECT 19.915000  2.805000 20.215000 3.335000 ;
      RECT 19.965000  0.085000 20.180000 0.545000 ;
      RECT 19.965000  4.895000 20.180000 5.355000 ;
      RECT 20.350000  0.255000 21.495000 0.425000 ;
      RECT 20.350000  0.425000 20.655000 0.715000 ;
      RECT 20.350000  0.885000 20.655000 0.925000 ;
      RECT 20.350000  4.515000 20.655000 4.555000 ;
      RECT 20.350000  4.725000 20.655000 5.015000 ;
      RECT 20.350000  5.015000 21.495000 5.185000 ;
      RECT 20.435000  1.665000 20.605000 2.295000 ;
      RECT 20.435000  2.295000 20.735000 2.465000 ;
      RECT 20.435000  2.975000 20.735000 3.145000 ;
      RECT 20.435000  3.145000 20.605000 3.775000 ;
      RECT 20.785000  1.755000 21.215000 2.125000 ;
      RECT 20.785000  3.315000 21.215000 3.685000 ;
      RECT 20.825000  0.595000 21.155000 0.885000 ;
      RECT 20.825000  4.555000 21.155000 4.845000 ;
      RECT 20.905000  0.885000 21.075000 1.755000 ;
      RECT 20.905000  2.125000 21.075000 3.315000 ;
      RECT 20.905000  3.685000 21.075000 4.555000 ;
      RECT 21.245000  2.295000 21.600000 2.465000 ;
      RECT 21.245000  2.635000 23.835000 2.805000 ;
      RECT 21.245000  2.975000 21.600000 3.145000 ;
      RECT 21.325000  0.425000 21.495000 0.770000 ;
      RECT 21.325000  4.670000 21.495000 5.015000 ;
      RECT 21.420000  1.205000 21.835000 1.305000 ;
      RECT 21.420000  1.305000 21.940000 1.465000 ;
      RECT 21.420000  1.465000 22.200000 1.475000 ;
      RECT 21.420000  3.965000 22.200000 3.975000 ;
      RECT 21.420000  3.975000 21.940000 4.135000 ;
      RECT 21.420000  4.135000 21.835000 4.235000 ;
      RECT 21.430000  1.645000 21.600000 2.295000 ;
      RECT 21.430000  3.145000 21.600000 3.795000 ;
      RECT 21.665000  0.585000 22.245000 0.755000 ;
      RECT 21.665000  0.755000 21.835000 1.205000 ;
      RECT 21.665000  4.235000 21.835000 4.685000 ;
      RECT 21.665000  4.685000 22.245000 4.855000 ;
      RECT 21.770000  1.475000 22.200000 1.635000 ;
      RECT 21.770000  3.805000 22.200000 3.965000 ;
      RECT 21.870000  1.635000 22.200000 2.465000 ;
      RECT 21.870000  2.975000 22.200000 3.805000 ;
      RECT 21.995000  0.330000 22.245000 0.585000 ;
      RECT 21.995000  4.855000 22.245000 5.110000 ;
      RECT 22.375000  1.465000 22.705000 2.635000 ;
      RECT 22.375000  2.805000 22.705000 3.975000 ;
      RECT 22.415000  0.085000 22.665000 0.660000 ;
      RECT 22.415000  4.780000 22.665000 5.355000 ;
      RECT 22.835000  0.330000 23.085000 0.585000 ;
      RECT 22.835000  0.585000 23.415000 0.755000 ;
      RECT 22.835000  4.685000 23.415000 4.855000 ;
      RECT 22.835000  4.855000 23.085000 5.110000 ;
      RECT 22.880000  1.465000 23.660000 1.475000 ;
      RECT 22.880000  1.475000 23.310000 1.635000 ;
      RECT 22.880000  1.635000 23.210000 2.465000 ;
      RECT 22.880000  2.975000 23.210000 3.805000 ;
      RECT 22.880000  3.805000 23.310000 3.965000 ;
      RECT 22.880000  3.965000 23.660000 3.975000 ;
      RECT 23.140000  1.305000 23.660000 1.465000 ;
      RECT 23.140000  3.975000 23.660000 4.135000 ;
      RECT 23.245000  0.755000 23.415000 1.205000 ;
      RECT 23.245000  1.205000 23.660000 1.305000 ;
      RECT 23.245000  4.135000 23.660000 4.235000 ;
      RECT 23.245000  4.235000 23.415000 4.685000 ;
      RECT 23.480000  1.645000 23.650000 2.295000 ;
      RECT 23.480000  2.295000 23.835000 2.465000 ;
      RECT 23.480000  2.975000 23.835000 3.145000 ;
      RECT 23.480000  3.145000 23.650000 3.795000 ;
      RECT 23.585000  0.255000 24.730000 0.425000 ;
      RECT 23.585000  0.425000 23.755000 0.770000 ;
      RECT 23.585000  4.670000 23.755000 5.015000 ;
      RECT 23.585000  5.015000 24.730000 5.185000 ;
      RECT 23.865000  1.755000 24.295000 2.125000 ;
      RECT 23.865000  3.315000 24.295000 3.685000 ;
      RECT 23.925000  0.595000 24.255000 0.885000 ;
      RECT 23.925000  4.555000 24.255000 4.845000 ;
      RECT 24.005000  0.885000 24.175000 1.755000 ;
      RECT 24.005000  2.125000 24.175000 3.315000 ;
      RECT 24.005000  3.685000 24.175000 4.555000 ;
      RECT 24.345000  2.295000 24.645000 2.465000 ;
      RECT 24.345000  2.635000 25.760000 2.805000 ;
      RECT 24.345000  2.975000 24.645000 3.145000 ;
      RECT 24.425000  0.425000 24.730000 0.715000 ;
      RECT 24.425000  0.715000 25.615000 0.885000 ;
      RECT 24.425000  0.885000 24.730000 0.925000 ;
      RECT 24.425000  4.515000 24.730000 4.555000 ;
      RECT 24.425000  4.555000 25.615000 4.725000 ;
      RECT 24.425000  4.725000 24.730000 5.015000 ;
      RECT 24.475000  1.495000 25.665000 1.665000 ;
      RECT 24.475000  1.665000 24.645000 2.295000 ;
      RECT 24.475000  3.145000 24.645000 3.775000 ;
      RECT 24.475000  3.775000 25.665000 3.945000 ;
      RECT 24.865000  1.835000 25.195000 2.105000 ;
      RECT 24.865000  2.105000 25.165000 2.635000 ;
      RECT 24.865000  2.805000 25.165000 3.335000 ;
      RECT 24.865000  3.335000 25.195000 3.605000 ;
      RECT 24.900000  0.085000 25.115000 0.545000 ;
      RECT 24.900000  4.895000 25.115000 5.355000 ;
      RECT 25.285000  0.255000 25.615000 0.715000 ;
      RECT 25.285000  4.725000 25.615000 5.185000 ;
      RECT 25.335000  2.210000 25.665000 2.465000 ;
      RECT 25.335000  2.975000 25.665000 3.230000 ;
      RECT 25.365000  1.665000 25.665000 2.210000 ;
      RECT 25.365000  3.230000 25.665000 3.775000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.145000  5.355000  0.315000 5.525000 ;
      RECT  0.175000  2.140000  0.345000 2.310000 ;
      RECT  0.175000  3.130000  0.345000 3.300000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.605000  5.355000  0.775000 5.525000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.065000  5.355000  1.235000 5.525000 ;
      RECT  1.115000  2.140000  1.285000 2.310000 ;
      RECT  1.115000  3.130000  1.285000 3.300000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.785000  1.695000 1.955000 ;
      RECT  1.525000  3.485000  1.695000 3.655000 ;
      RECT  1.525000  5.355000  1.695000 5.525000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  1.985000  5.355000  2.155000 5.525000 ;
      RECT  2.110000  2.140000  2.280000 2.310000 ;
      RECT  2.110000  3.130000  2.280000 3.300000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.445000  5.355000  2.615000 5.525000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  2.905000  5.355000  3.075000 5.525000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.365000  5.355000  3.535000 5.525000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  3.825000  5.355000  3.995000 5.525000 ;
      RECT  4.160000  2.140000  4.330000 2.310000 ;
      RECT  4.160000  3.130000  4.330000 3.300000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.285000  5.355000  4.455000 5.525000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.785000  4.915000 1.955000 ;
      RECT  4.745000  3.485000  4.915000 3.655000 ;
      RECT  4.745000  5.355000  4.915000 5.525000 ;
      RECT  5.155000  2.140000  5.325000 2.310000 ;
      RECT  5.155000  3.130000  5.325000 3.300000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.205000  5.355000  5.375000 5.525000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.665000  5.355000  5.835000 5.525000 ;
      RECT  6.095000  2.140000  6.265000 2.310000 ;
      RECT  6.095000  3.130000  6.265000 3.300000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.125000  5.355000  6.295000 5.525000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.585000  5.355000  6.755000 5.525000 ;
      RECT  6.615000  2.140000  6.785000 2.310000 ;
      RECT  6.615000  3.130000  6.785000 3.300000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.045000  5.355000  7.215000 5.525000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.505000  5.355000  7.675000 5.525000 ;
      RECT  7.555000  2.140000  7.725000 2.310000 ;
      RECT  7.555000  3.130000  7.725000 3.300000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  1.785000  8.135000 1.955000 ;
      RECT  7.965000  3.485000  8.135000 3.655000 ;
      RECT  7.965000  5.355000  8.135000 5.525000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.425000  5.355000  8.595000 5.525000 ;
      RECT  8.550000  2.140000  8.720000 2.310000 ;
      RECT  8.550000  3.130000  8.720000 3.300000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.885000  5.355000  9.055000 5.525000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.345000  5.355000  9.515000 5.525000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT  9.805000  5.355000  9.975000 5.525000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.265000  5.355000 10.435000 5.525000 ;
      RECT 10.600000  2.140000 10.770000 2.310000 ;
      RECT 10.600000  3.130000 10.770000 3.300000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.725000  5.355000 10.895000 5.525000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  1.785000 11.355000 1.955000 ;
      RECT 11.185000  3.485000 11.355000 3.655000 ;
      RECT 11.185000  5.355000 11.355000 5.525000 ;
      RECT 11.595000  2.140000 11.765000 2.310000 ;
      RECT 11.595000  3.130000 11.765000 3.300000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 11.645000  5.355000 11.815000 5.525000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.105000  5.355000 12.275000 5.525000 ;
      RECT 12.535000  2.140000 12.705000 2.310000 ;
      RECT 12.535000  3.130000 12.705000 3.300000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 12.565000  5.355000 12.735000 5.525000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.025000  5.355000 13.195000 5.525000 ;
      RECT 13.055000  2.140000 13.225000 2.310000 ;
      RECT 13.055000  3.130000 13.225000 3.300000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.485000  5.355000 13.655000 5.525000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 13.945000  5.355000 14.115000 5.525000 ;
      RECT 13.995000  2.140000 14.165000 2.310000 ;
      RECT 13.995000  3.130000 14.165000 3.300000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  1.785000 14.575000 1.955000 ;
      RECT 14.405000  3.485000 14.575000 3.655000 ;
      RECT 14.405000  5.355000 14.575000 5.525000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 14.865000  5.355000 15.035000 5.525000 ;
      RECT 14.990000  2.140000 15.160000 2.310000 ;
      RECT 14.990000  3.130000 15.160000 3.300000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.325000  5.355000 15.495000 5.525000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 15.785000  5.355000 15.955000 5.525000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.245000  5.355000 16.415000 5.525000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
      RECT 16.705000  5.355000 16.875000 5.525000 ;
      RECT 17.040000  2.140000 17.210000 2.310000 ;
      RECT 17.040000  3.130000 17.210000 3.300000 ;
      RECT 17.165000 -0.085000 17.335000 0.085000 ;
      RECT 17.165000  2.635000 17.335000 2.805000 ;
      RECT 17.165000  5.355000 17.335000 5.525000 ;
      RECT 17.625000 -0.085000 17.795000 0.085000 ;
      RECT 17.625000  1.785000 17.795000 1.955000 ;
      RECT 17.625000  3.485000 17.795000 3.655000 ;
      RECT 17.625000  5.355000 17.795000 5.525000 ;
      RECT 18.035000  2.140000 18.205000 2.310000 ;
      RECT 18.035000  3.130000 18.205000 3.300000 ;
      RECT 18.085000 -0.085000 18.255000 0.085000 ;
      RECT 18.085000  2.635000 18.255000 2.805000 ;
      RECT 18.085000  5.355000 18.255000 5.525000 ;
      RECT 18.545000 -0.085000 18.715000 0.085000 ;
      RECT 18.545000  2.635000 18.715000 2.805000 ;
      RECT 18.545000  5.355000 18.715000 5.525000 ;
      RECT 18.975000  2.140000 19.145000 2.310000 ;
      RECT 18.975000  3.130000 19.145000 3.300000 ;
      RECT 19.005000 -0.085000 19.175000 0.085000 ;
      RECT 19.005000  2.635000 19.175000 2.805000 ;
      RECT 19.005000  5.355000 19.175000 5.525000 ;
      RECT 19.465000 -0.085000 19.635000 0.085000 ;
      RECT 19.465000  2.635000 19.635000 2.805000 ;
      RECT 19.465000  5.355000 19.635000 5.525000 ;
      RECT 19.495000  2.140000 19.665000 2.310000 ;
      RECT 19.495000  3.130000 19.665000 3.300000 ;
      RECT 19.925000 -0.085000 20.095000 0.085000 ;
      RECT 19.925000  2.635000 20.095000 2.805000 ;
      RECT 19.925000  5.355000 20.095000 5.525000 ;
      RECT 20.385000 -0.085000 20.555000 0.085000 ;
      RECT 20.385000  2.635000 20.555000 2.805000 ;
      RECT 20.385000  5.355000 20.555000 5.525000 ;
      RECT 20.435000  2.140000 20.605000 2.310000 ;
      RECT 20.435000  3.130000 20.605000 3.300000 ;
      RECT 20.845000 -0.085000 21.015000 0.085000 ;
      RECT 20.845000  1.785000 21.015000 1.955000 ;
      RECT 20.845000  3.485000 21.015000 3.655000 ;
      RECT 20.845000  5.355000 21.015000 5.525000 ;
      RECT 21.305000 -0.085000 21.475000 0.085000 ;
      RECT 21.305000  2.635000 21.475000 2.805000 ;
      RECT 21.305000  5.355000 21.475000 5.525000 ;
      RECT 21.430000  2.140000 21.600000 2.310000 ;
      RECT 21.430000  3.130000 21.600000 3.300000 ;
      RECT 21.765000 -0.085000 21.935000 0.085000 ;
      RECT 21.765000  2.635000 21.935000 2.805000 ;
      RECT 21.765000  5.355000 21.935000 5.525000 ;
      RECT 22.225000 -0.085000 22.395000 0.085000 ;
      RECT 22.225000  2.635000 22.395000 2.805000 ;
      RECT 22.225000  5.355000 22.395000 5.525000 ;
      RECT 22.685000 -0.085000 22.855000 0.085000 ;
      RECT 22.685000  2.635000 22.855000 2.805000 ;
      RECT 22.685000  5.355000 22.855000 5.525000 ;
      RECT 23.145000 -0.085000 23.315000 0.085000 ;
      RECT 23.145000  2.635000 23.315000 2.805000 ;
      RECT 23.145000  5.355000 23.315000 5.525000 ;
      RECT 23.480000  2.140000 23.650000 2.310000 ;
      RECT 23.480000  3.130000 23.650000 3.300000 ;
      RECT 23.605000 -0.085000 23.775000 0.085000 ;
      RECT 23.605000  2.635000 23.775000 2.805000 ;
      RECT 23.605000  5.355000 23.775000 5.525000 ;
      RECT 24.065000 -0.085000 24.235000 0.085000 ;
      RECT 24.065000  1.785000 24.235000 1.955000 ;
      RECT 24.065000  3.485000 24.235000 3.655000 ;
      RECT 24.065000  5.355000 24.235000 5.525000 ;
      RECT 24.475000  2.140000 24.645000 2.310000 ;
      RECT 24.475000  3.130000 24.645000 3.300000 ;
      RECT 24.525000 -0.085000 24.695000 0.085000 ;
      RECT 24.525000  2.635000 24.695000 2.805000 ;
      RECT 24.525000  5.355000 24.695000 5.525000 ;
      RECT 24.985000 -0.085000 25.155000 0.085000 ;
      RECT 24.985000  2.635000 25.155000 2.805000 ;
      RECT 24.985000  5.355000 25.155000 5.525000 ;
      RECT 25.415000  2.140000 25.585000 2.310000 ;
      RECT 25.415000  3.130000 25.585000 3.300000 ;
      RECT 25.445000 -0.085000 25.615000 0.085000 ;
      RECT 25.445000  2.635000 25.615000 2.805000 ;
      RECT 25.445000  5.355000 25.615000 5.525000 ;
    LAYER met1 ;
      RECT  0.115000 2.110000  0.405000 2.155000 ;
      RECT  0.115000 2.155000  2.340000 2.295000 ;
      RECT  0.115000 2.295000  0.405000 2.340000 ;
      RECT  0.115000 3.100000  0.405000 3.145000 ;
      RECT  0.115000 3.145000  2.340000 3.285000 ;
      RECT  0.115000 3.285000  0.405000 3.330000 ;
      RECT  1.055000 2.110000  1.345000 2.155000 ;
      RECT  1.055000 2.295000  1.345000 2.340000 ;
      RECT  1.055000 3.100000  1.345000 3.145000 ;
      RECT  1.055000 3.285000  1.345000 3.330000 ;
      RECT  2.050000 2.110000  2.340000 2.155000 ;
      RECT  2.050000 2.295000  2.340000 2.340000 ;
      RECT  2.050000 3.100000  2.340000 3.145000 ;
      RECT  2.050000 3.285000  2.340000 3.330000 ;
      RECT  4.100000 2.110000  4.390000 2.155000 ;
      RECT  4.100000 2.155000  6.325000 2.295000 ;
      RECT  4.100000 2.295000  4.390000 2.340000 ;
      RECT  4.100000 3.100000  4.390000 3.145000 ;
      RECT  4.100000 3.145000  6.325000 3.285000 ;
      RECT  4.100000 3.285000  4.390000 3.330000 ;
      RECT  5.095000 2.110000  5.385000 2.155000 ;
      RECT  5.095000 2.295000  5.385000 2.340000 ;
      RECT  5.095000 3.100000  5.385000 3.145000 ;
      RECT  5.095000 3.285000  5.385000 3.330000 ;
      RECT  6.035000 2.110000  6.325000 2.155000 ;
      RECT  6.035000 2.295000  6.325000 2.340000 ;
      RECT  6.035000 3.100000  6.325000 3.145000 ;
      RECT  6.035000 3.285000  6.325000 3.330000 ;
      RECT  6.555000 2.110000  6.845000 2.155000 ;
      RECT  6.555000 2.155000  8.780000 2.295000 ;
      RECT  6.555000 2.295000  6.845000 2.340000 ;
      RECT  6.555000 3.100000  6.845000 3.145000 ;
      RECT  6.555000 3.145000  8.780000 3.285000 ;
      RECT  6.555000 3.285000  6.845000 3.330000 ;
      RECT  7.495000 2.110000  7.785000 2.155000 ;
      RECT  7.495000 2.295000  7.785000 2.340000 ;
      RECT  7.495000 3.100000  7.785000 3.145000 ;
      RECT  7.495000 3.285000  7.785000 3.330000 ;
      RECT  8.490000 2.110000  8.780000 2.155000 ;
      RECT  8.490000 2.295000  8.780000 2.340000 ;
      RECT  8.490000 3.100000  8.780000 3.145000 ;
      RECT  8.490000 3.285000  8.780000 3.330000 ;
      RECT 10.540000 2.110000 10.830000 2.155000 ;
      RECT 10.540000 2.155000 12.765000 2.295000 ;
      RECT 10.540000 2.295000 10.830000 2.340000 ;
      RECT 10.540000 3.100000 10.830000 3.145000 ;
      RECT 10.540000 3.145000 12.765000 3.285000 ;
      RECT 10.540000 3.285000 10.830000 3.330000 ;
      RECT 11.535000 2.110000 11.825000 2.155000 ;
      RECT 11.535000 2.295000 11.825000 2.340000 ;
      RECT 11.535000 3.100000 11.825000 3.145000 ;
      RECT 11.535000 3.285000 11.825000 3.330000 ;
      RECT 12.475000 2.110000 12.765000 2.155000 ;
      RECT 12.475000 2.295000 12.765000 2.340000 ;
      RECT 12.475000 3.100000 12.765000 3.145000 ;
      RECT 12.475000 3.285000 12.765000 3.330000 ;
      RECT 12.995000 2.110000 13.285000 2.155000 ;
      RECT 12.995000 2.155000 15.220000 2.295000 ;
      RECT 12.995000 2.295000 13.285000 2.340000 ;
      RECT 12.995000 3.100000 13.285000 3.145000 ;
      RECT 12.995000 3.145000 15.220000 3.285000 ;
      RECT 12.995000 3.285000 13.285000 3.330000 ;
      RECT 13.935000 2.110000 14.225000 2.155000 ;
      RECT 13.935000 2.295000 14.225000 2.340000 ;
      RECT 13.935000 3.100000 14.225000 3.145000 ;
      RECT 13.935000 3.285000 14.225000 3.330000 ;
      RECT 14.930000 2.110000 15.220000 2.155000 ;
      RECT 14.930000 2.295000 15.220000 2.340000 ;
      RECT 14.930000 3.100000 15.220000 3.145000 ;
      RECT 14.930000 3.285000 15.220000 3.330000 ;
      RECT 16.980000 2.110000 17.270000 2.155000 ;
      RECT 16.980000 2.155000 19.205000 2.295000 ;
      RECT 16.980000 2.295000 17.270000 2.340000 ;
      RECT 16.980000 3.100000 17.270000 3.145000 ;
      RECT 16.980000 3.145000 19.205000 3.285000 ;
      RECT 16.980000 3.285000 17.270000 3.330000 ;
      RECT 17.975000 2.110000 18.265000 2.155000 ;
      RECT 17.975000 2.295000 18.265000 2.340000 ;
      RECT 17.975000 3.100000 18.265000 3.145000 ;
      RECT 17.975000 3.285000 18.265000 3.330000 ;
      RECT 18.915000 2.110000 19.205000 2.155000 ;
      RECT 18.915000 2.295000 19.205000 2.340000 ;
      RECT 18.915000 3.100000 19.205000 3.145000 ;
      RECT 18.915000 3.285000 19.205000 3.330000 ;
      RECT 19.435000 2.110000 19.725000 2.155000 ;
      RECT 19.435000 2.155000 21.660000 2.295000 ;
      RECT 19.435000 2.295000 19.725000 2.340000 ;
      RECT 19.435000 3.100000 19.725000 3.145000 ;
      RECT 19.435000 3.145000 21.660000 3.285000 ;
      RECT 19.435000 3.285000 19.725000 3.330000 ;
      RECT 20.375000 2.110000 20.665000 2.155000 ;
      RECT 20.375000 2.295000 20.665000 2.340000 ;
      RECT 20.375000 3.100000 20.665000 3.145000 ;
      RECT 20.375000 3.285000 20.665000 3.330000 ;
      RECT 21.370000 2.110000 21.660000 2.155000 ;
      RECT 21.370000 2.295000 21.660000 2.340000 ;
      RECT 21.370000 3.100000 21.660000 3.145000 ;
      RECT 21.370000 3.285000 21.660000 3.330000 ;
      RECT 23.420000 2.110000 23.710000 2.155000 ;
      RECT 23.420000 2.155000 25.645000 2.295000 ;
      RECT 23.420000 2.295000 23.710000 2.340000 ;
      RECT 23.420000 3.100000 23.710000 3.145000 ;
      RECT 23.420000 3.145000 25.645000 3.285000 ;
      RECT 23.420000 3.285000 23.710000 3.330000 ;
      RECT 24.415000 2.110000 24.705000 2.155000 ;
      RECT 24.415000 2.295000 24.705000 2.340000 ;
      RECT 24.415000 3.100000 24.705000 3.145000 ;
      RECT 24.415000 3.285000 24.705000 3.330000 ;
      RECT 25.355000 2.110000 25.645000 2.155000 ;
      RECT 25.355000 2.295000 25.645000 2.340000 ;
      RECT 25.355000 3.100000 25.645000 3.145000 ;
      RECT 25.355000 3.285000 25.645000 3.330000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb16to1_2


MACRO sky130_fd_sc_hdll__muxb16to1_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  51.98000 BY  5.440000 ;
  SITE unithd ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 1.055000 1.785000 1.325000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.095000 1.055000 12.485000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.275000 1.055000 14.665000 1.325000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 23.975000 1.055000 25.365000 1.325000 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 26.615000 1.055000 28.005000 1.325000 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 37.315000 1.055000 38.705000 1.325000 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 39.495000 1.055000 40.885000 1.325000 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 50.195000 1.055000 51.585000 1.325000 ;
    END
  END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 4.115000 1.785000 4.385000 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.095000 4.115000 12.485000 4.385000 ;
    END
  END D[9]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.275000 4.115000 14.665000 4.385000 ;
    END
  END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 23.975000 4.115000 25.365000 4.385000 ;
    END
  END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 26.615000 4.115000 28.005000 4.385000 ;
    END
  END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 37.315000 4.115000 38.705000 4.385000 ;
    END
  END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 39.495000 4.115000 40.885000 4.385000 ;
    END
  END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 50.195000 4.115000 51.585000 4.385000 ;
    END
  END D[15]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 0.995000 6.355000 1.325000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.525000 0.995000 7.120000 1.325000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.640000 0.995000 19.235000 1.325000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.405000 0.995000 20.000000 1.325000 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.980000 0.995000 32.575000 1.325000 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 32.745000 0.995000 33.340000 1.325000 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 44.860000 0.995000 45.455000 1.325000 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 45.625000 0.995000 46.220000 1.325000 ;
    END
  END S[7]
  PIN S[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 4.115000 6.355000 4.445000 ;
    END
  END S[8]
  PIN S[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.525000 4.115000 7.120000 4.445000 ;
    END
  END S[9]
  PIN S[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.640000 4.115000 19.235000 4.445000 ;
    END
  END S[10]
  PIN S[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.405000 4.115000 20.000000 4.445000 ;
    END
  END S[11]
  PIN S[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.980000 4.115000 32.575000 4.445000 ;
    END
  END S[12]
  PIN S[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 32.745000 4.115000 33.340000 4.445000 ;
    END
  END S[13]
  PIN S[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 44.860000 4.115000 45.455000 4.445000 ;
    END
  END S[14]
  PIN S[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 45.625000 4.115000 46.220000 4.445000 ;
    END
  END S[15]
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  2.985000 1.755000  3.275000 1.800000 ;
        RECT  2.985000 1.800000 48.995000 1.940000 ;
        RECT  2.985000 1.940000  3.275000 1.985000 ;
        RECT  2.985000 3.455000  3.275000 3.500000 ;
        RECT  2.985000 3.500000 48.995000 3.640000 ;
        RECT  2.985000 3.640000  3.275000 3.685000 ;
        RECT  3.925000 1.755000  4.215000 1.800000 ;
        RECT  3.925000 1.940000  4.215000 1.985000 ;
        RECT  3.925000 3.455000  4.215000 3.500000 ;
        RECT  3.925000 3.640000  4.215000 3.685000 ;
        RECT  8.665000 1.755000  8.955000 1.800000 ;
        RECT  8.665000 1.940000  8.955000 1.985000 ;
        RECT  8.665000 3.455000  8.955000 3.500000 ;
        RECT  8.665000 3.640000  8.955000 3.685000 ;
        RECT  9.605000 1.755000  9.895000 1.800000 ;
        RECT  9.605000 1.940000  9.895000 1.985000 ;
        RECT  9.605000 3.455000  9.895000 3.500000 ;
        RECT  9.605000 3.640000  9.895000 3.685000 ;
        RECT 15.865000 1.755000 16.155000 1.800000 ;
        RECT 15.865000 1.940000 16.155000 1.985000 ;
        RECT 15.865000 3.455000 16.155000 3.500000 ;
        RECT 15.865000 3.640000 16.155000 3.685000 ;
        RECT 16.805000 1.755000 17.095000 1.800000 ;
        RECT 16.805000 1.940000 17.095000 1.985000 ;
        RECT 16.805000 3.455000 17.095000 3.500000 ;
        RECT 16.805000 3.640000 17.095000 3.685000 ;
        RECT 21.545000 1.755000 21.835000 1.800000 ;
        RECT 21.545000 1.940000 21.835000 1.985000 ;
        RECT 21.545000 3.455000 21.835000 3.500000 ;
        RECT 21.545000 3.640000 21.835000 3.685000 ;
        RECT 22.485000 1.755000 22.775000 1.800000 ;
        RECT 22.485000 1.940000 22.775000 1.985000 ;
        RECT 22.485000 3.455000 22.775000 3.500000 ;
        RECT 22.485000 3.640000 22.775000 3.685000 ;
        RECT 29.205000 1.755000 29.495000 1.800000 ;
        RECT 29.205000 1.940000 29.495000 1.985000 ;
        RECT 29.205000 3.455000 29.495000 3.500000 ;
        RECT 29.205000 3.640000 29.495000 3.685000 ;
        RECT 30.145000 1.755000 30.435000 1.800000 ;
        RECT 30.145000 1.940000 30.435000 1.985000 ;
        RECT 30.145000 3.455000 30.435000 3.500000 ;
        RECT 30.145000 3.640000 30.435000 3.685000 ;
        RECT 34.885000 1.755000 35.175000 1.800000 ;
        RECT 34.885000 1.940000 35.175000 1.985000 ;
        RECT 34.885000 3.455000 35.175000 3.500000 ;
        RECT 34.885000 3.640000 35.175000 3.685000 ;
        RECT 35.825000 1.755000 36.115000 1.800000 ;
        RECT 35.825000 1.940000 36.115000 1.985000 ;
        RECT 35.825000 3.455000 36.115000 3.500000 ;
        RECT 35.825000 3.640000 36.115000 3.685000 ;
        RECT 42.085000 1.755000 42.375000 1.800000 ;
        RECT 42.085000 1.940000 42.375000 1.985000 ;
        RECT 42.085000 3.455000 42.375000 3.500000 ;
        RECT 42.085000 3.640000 42.375000 3.685000 ;
        RECT 43.025000 1.755000 43.315000 1.800000 ;
        RECT 43.025000 1.940000 43.315000 1.985000 ;
        RECT 43.025000 3.455000 43.315000 3.500000 ;
        RECT 43.025000 3.640000 43.315000 3.685000 ;
        RECT 47.765000 1.755000 48.055000 1.800000 ;
        RECT 47.765000 1.940000 48.055000 1.985000 ;
        RECT 47.765000 3.455000 48.055000 3.500000 ;
        RECT 47.765000 3.640000 48.055000 3.685000 ;
        RECT 48.705000 1.755000 48.995000 1.800000 ;
        RECT 48.705000 1.940000 48.995000 1.985000 ;
        RECT 48.705000 3.455000 48.995000 3.500000 ;
        RECT 48.705000 3.640000 48.995000 3.685000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 51.980000 0.240000 ;
        RECT 0.000000  5.200000 51.980000 5.680000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 51.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 51.980000 0.085000 ;
      RECT  0.000000  2.635000  2.795000 2.805000 ;
      RECT  0.000000  5.355000 51.980000 5.525000 ;
      RECT  0.125000  1.495000  0.395000 2.635000 ;
      RECT  0.125000  2.805000  0.395000 3.945000 ;
      RECT  0.145000  0.085000  0.395000 0.885000 ;
      RECT  0.145000  4.555000  0.395000 5.355000 ;
      RECT  0.565000  0.255000  0.895000 0.715000 ;
      RECT  0.565000  0.715000  2.695000 0.885000 ;
      RECT  0.565000  1.495000  2.795000 1.665000 ;
      RECT  0.565000  1.665000  0.895000 2.465000 ;
      RECT  0.565000  2.975000  0.895000 3.775000 ;
      RECT  0.565000  3.775000  2.795000 3.945000 ;
      RECT  0.565000  4.555000  2.695000 4.725000 ;
      RECT  0.565000  4.725000  0.895000 5.185000 ;
      RECT  1.065000  0.085000  1.335000 0.545000 ;
      RECT  1.065000  1.835000  1.335000 2.635000 ;
      RECT  1.065000  2.805000  1.335000 3.605000 ;
      RECT  1.065000  4.895000  1.335000 5.355000 ;
      RECT  1.505000  0.255000  1.835000 0.715000 ;
      RECT  1.505000  1.665000  1.835000 2.465000 ;
      RECT  1.505000  2.975000  1.835000 3.775000 ;
      RECT  1.505000  4.725000  1.835000 5.185000 ;
      RECT  2.005000  0.085000  2.255000 0.545000 ;
      RECT  2.005000  1.835000  2.275000 2.635000 ;
      RECT  2.005000  2.805000  2.275000 3.605000 ;
      RECT  2.005000  4.895000  2.255000 5.355000 ;
      RECT  2.425000  0.255000  4.455000 0.425000 ;
      RECT  2.425000  0.425000  2.695000 0.715000 ;
      RECT  2.425000  4.725000  2.695000 5.015000 ;
      RECT  2.425000  5.015000  4.455000 5.185000 ;
      RECT  2.495000  1.665000  2.795000 2.465000 ;
      RECT  2.495000  2.975000  2.795000 3.775000 ;
      RECT  2.865000  0.595000  3.195000 0.885000 ;
      RECT  2.865000  4.555000  3.195000 4.845000 ;
      RECT  2.965000  0.885000  3.195000 1.065000 ;
      RECT  2.965000  1.065000  4.235000 1.365000 ;
      RECT  2.965000  1.365000  3.295000 4.075000 ;
      RECT  2.965000  4.075000  4.235000 4.375000 ;
      RECT  2.965000  4.375000  3.195000 4.555000 ;
      RECT  3.365000  0.425000  3.535000 0.770000 ;
      RECT  3.365000  4.670000  3.535000 5.015000 ;
      RECT  3.465000  1.535000  3.735000 2.465000 ;
      RECT  3.465000  2.975000  3.735000 3.905000 ;
      RECT  3.705000  0.595000  4.035000 1.065000 ;
      RECT  3.705000  4.375000  4.035000 4.845000 ;
      RECT  3.905000  1.365000  4.235000 4.075000 ;
      RECT  4.205000  0.425000  4.455000 0.770000 ;
      RECT  4.205000  4.670000  4.455000 5.015000 ;
      RECT  4.405000  1.065000  5.590000 1.395000 ;
      RECT  4.405000  1.565000  4.705000 2.465000 ;
      RECT  4.405000  2.635000  8.475000 2.805000 ;
      RECT  4.405000  2.975000  4.705000 3.875000 ;
      RECT  4.405000  4.045000  5.590000 4.375000 ;
      RECT  4.950000  1.605000  5.225000 2.635000 ;
      RECT  4.950000  2.805000  5.225000 3.835000 ;
      RECT  4.960000  0.085000  5.250000 0.610000 ;
      RECT  4.960000  4.830000  5.250000 5.355000 ;
      RECT  5.420000  0.280000  5.670000 0.825000 ;
      RECT  5.420000  0.825000  5.590000 1.065000 ;
      RECT  5.420000  1.395000  5.590000 1.605000 ;
      RECT  5.420000  1.605000  5.750000 2.465000 ;
      RECT  5.420000  2.975000  5.750000 3.835000 ;
      RECT  5.420000  3.835000  5.590000 4.045000 ;
      RECT  5.420000  4.375000  5.590000 4.615000 ;
      RECT  5.420000  4.615000  5.670000 5.160000 ;
      RECT  5.880000  0.085000  6.170000 0.610000 ;
      RECT  5.880000  4.830000  6.170000 5.355000 ;
      RECT  5.920000  1.605000  6.220000 2.635000 ;
      RECT  5.920000  2.805000  6.220000 3.835000 ;
      RECT  6.660000  1.605000  6.960000 2.635000 ;
      RECT  6.660000  2.805000  6.960000 3.835000 ;
      RECT  6.710000  0.085000  7.000000 0.610000 ;
      RECT  6.710000  4.830000  7.000000 5.355000 ;
      RECT  7.130000  1.605000  7.460000 2.465000 ;
      RECT  7.130000  2.975000  7.460000 3.835000 ;
      RECT  7.210000  0.280000  7.460000 0.825000 ;
      RECT  7.210000  4.615000  7.460000 5.160000 ;
      RECT  7.290000  0.825000  7.460000 1.065000 ;
      RECT  7.290000  1.065000  8.475000 1.395000 ;
      RECT  7.290000  1.395000  7.460000 1.605000 ;
      RECT  7.290000  3.835000  7.460000 4.045000 ;
      RECT  7.290000  4.045000  8.475000 4.375000 ;
      RECT  7.290000  4.375000  7.460000 4.615000 ;
      RECT  7.630000  0.085000  7.920000 0.610000 ;
      RECT  7.630000  4.830000  7.920000 5.355000 ;
      RECT  7.655000  1.605000  7.930000 2.635000 ;
      RECT  7.655000  2.805000  7.930000 3.835000 ;
      RECT  8.175000  1.565000  8.475000 2.465000 ;
      RECT  8.175000  2.975000  8.475000 3.875000 ;
      RECT  8.425000  0.255000 10.455000 0.425000 ;
      RECT  8.425000  0.425000  8.675000 0.770000 ;
      RECT  8.425000  4.670000  8.675000 5.015000 ;
      RECT  8.425000  5.015000 10.455000 5.185000 ;
      RECT  8.645000  1.065000  9.915000 1.365000 ;
      RECT  8.645000  1.365000  8.975000 4.075000 ;
      RECT  8.645000  4.075000  9.915000 4.375000 ;
      RECT  8.845000  0.595000  9.175000 1.065000 ;
      RECT  8.845000  4.375000  9.175000 4.845000 ;
      RECT  9.145000  1.535000  9.415000 2.465000 ;
      RECT  9.145000  2.975000  9.415000 3.905000 ;
      RECT  9.345000  0.425000  9.515000 0.770000 ;
      RECT  9.345000  4.670000  9.515000 5.015000 ;
      RECT  9.585000  1.365000  9.915000 4.075000 ;
      RECT  9.685000  0.595000 10.015000 0.885000 ;
      RECT  9.685000  0.885000  9.915000 1.065000 ;
      RECT  9.685000  4.375000  9.915000 4.555000 ;
      RECT  9.685000  4.555000 10.015000 4.845000 ;
      RECT 10.085000  1.495000 12.315000 1.665000 ;
      RECT 10.085000  1.665000 10.385000 2.465000 ;
      RECT 10.085000  2.635000 15.675000 2.805000 ;
      RECT 10.085000  2.975000 10.385000 3.775000 ;
      RECT 10.085000  3.775000 12.315000 3.945000 ;
      RECT 10.185000  0.425000 10.455000 0.715000 ;
      RECT 10.185000  0.715000 12.315000 0.885000 ;
      RECT 10.185000  4.555000 12.315000 4.725000 ;
      RECT 10.185000  4.725000 10.455000 5.015000 ;
      RECT 10.605000  1.835000 10.875000 2.635000 ;
      RECT 10.605000  2.805000 10.875000 3.605000 ;
      RECT 10.625000  0.085000 10.875000 0.545000 ;
      RECT 10.625000  4.895000 10.875000 5.355000 ;
      RECT 11.045000  0.255000 11.375000 0.715000 ;
      RECT 11.045000  1.665000 11.375000 2.465000 ;
      RECT 11.045000  2.975000 11.375000 3.775000 ;
      RECT 11.045000  4.725000 11.375000 5.185000 ;
      RECT 11.545000  0.085000 11.815000 0.545000 ;
      RECT 11.545000  1.835000 11.815000 2.635000 ;
      RECT 11.545000  2.805000 11.815000 3.605000 ;
      RECT 11.545000  4.895000 11.815000 5.355000 ;
      RECT 11.985000  0.255000 12.315000 0.715000 ;
      RECT 11.985000  1.665000 12.315000 2.465000 ;
      RECT 11.985000  2.975000 12.315000 3.775000 ;
      RECT 11.985000  4.725000 12.315000 5.185000 ;
      RECT 12.485000  0.085000 12.735000 0.885000 ;
      RECT 12.485000  1.495000 12.755000 2.635000 ;
      RECT 12.485000  2.805000 12.755000 3.945000 ;
      RECT 12.485000  4.555000 12.735000 5.355000 ;
      RECT 13.005000  1.495000 13.275000 2.635000 ;
      RECT 13.005000  2.805000 13.275000 3.945000 ;
      RECT 13.025000  0.085000 13.275000 0.885000 ;
      RECT 13.025000  4.555000 13.275000 5.355000 ;
      RECT 13.445000  0.255000 13.775000 0.715000 ;
      RECT 13.445000  0.715000 15.575000 0.885000 ;
      RECT 13.445000  1.495000 15.675000 1.665000 ;
      RECT 13.445000  1.665000 13.775000 2.465000 ;
      RECT 13.445000  2.975000 13.775000 3.775000 ;
      RECT 13.445000  3.775000 15.675000 3.945000 ;
      RECT 13.445000  4.555000 15.575000 4.725000 ;
      RECT 13.445000  4.725000 13.775000 5.185000 ;
      RECT 13.945000  0.085000 14.215000 0.545000 ;
      RECT 13.945000  1.835000 14.215000 2.635000 ;
      RECT 13.945000  2.805000 14.215000 3.605000 ;
      RECT 13.945000  4.895000 14.215000 5.355000 ;
      RECT 14.385000  0.255000 14.715000 0.715000 ;
      RECT 14.385000  1.665000 14.715000 2.465000 ;
      RECT 14.385000  2.975000 14.715000 3.775000 ;
      RECT 14.385000  4.725000 14.715000 5.185000 ;
      RECT 14.885000  0.085000 15.135000 0.545000 ;
      RECT 14.885000  1.835000 15.155000 2.635000 ;
      RECT 14.885000  2.805000 15.155000 3.605000 ;
      RECT 14.885000  4.895000 15.135000 5.355000 ;
      RECT 15.305000  0.255000 17.335000 0.425000 ;
      RECT 15.305000  0.425000 15.575000 0.715000 ;
      RECT 15.305000  4.725000 15.575000 5.015000 ;
      RECT 15.305000  5.015000 17.335000 5.185000 ;
      RECT 15.375000  1.665000 15.675000 2.465000 ;
      RECT 15.375000  2.975000 15.675000 3.775000 ;
      RECT 15.745000  0.595000 16.075000 0.885000 ;
      RECT 15.745000  4.555000 16.075000 4.845000 ;
      RECT 15.845000  0.885000 16.075000 1.065000 ;
      RECT 15.845000  1.065000 17.115000 1.365000 ;
      RECT 15.845000  1.365000 16.175000 4.075000 ;
      RECT 15.845000  4.075000 17.115000 4.375000 ;
      RECT 15.845000  4.375000 16.075000 4.555000 ;
      RECT 16.245000  0.425000 16.415000 0.770000 ;
      RECT 16.245000  4.670000 16.415000 5.015000 ;
      RECT 16.345000  1.535000 16.615000 2.465000 ;
      RECT 16.345000  2.975000 16.615000 3.905000 ;
      RECT 16.585000  0.595000 16.915000 1.065000 ;
      RECT 16.585000  4.375000 16.915000 4.845000 ;
      RECT 16.785000  1.365000 17.115000 4.075000 ;
      RECT 17.085000  0.425000 17.335000 0.770000 ;
      RECT 17.085000  4.670000 17.335000 5.015000 ;
      RECT 17.285000  1.065000 18.470000 1.395000 ;
      RECT 17.285000  1.565000 17.585000 2.465000 ;
      RECT 17.285000  2.635000 21.355000 2.805000 ;
      RECT 17.285000  2.975000 17.585000 3.875000 ;
      RECT 17.285000  4.045000 18.470000 4.375000 ;
      RECT 17.830000  1.605000 18.105000 2.635000 ;
      RECT 17.830000  2.805000 18.105000 3.835000 ;
      RECT 17.840000  0.085000 18.130000 0.610000 ;
      RECT 17.840000  4.830000 18.130000 5.355000 ;
      RECT 18.300000  0.280000 18.550000 0.825000 ;
      RECT 18.300000  0.825000 18.470000 1.065000 ;
      RECT 18.300000  1.395000 18.470000 1.605000 ;
      RECT 18.300000  1.605000 18.630000 2.465000 ;
      RECT 18.300000  2.975000 18.630000 3.835000 ;
      RECT 18.300000  3.835000 18.470000 4.045000 ;
      RECT 18.300000  4.375000 18.470000 4.615000 ;
      RECT 18.300000  4.615000 18.550000 5.160000 ;
      RECT 18.760000  0.085000 19.050000 0.610000 ;
      RECT 18.760000  4.830000 19.050000 5.355000 ;
      RECT 18.800000  1.605000 19.100000 2.635000 ;
      RECT 18.800000  2.805000 19.100000 3.835000 ;
      RECT 19.540000  1.605000 19.840000 2.635000 ;
      RECT 19.540000  2.805000 19.840000 3.835000 ;
      RECT 19.590000  0.085000 19.880000 0.610000 ;
      RECT 19.590000  4.830000 19.880000 5.355000 ;
      RECT 20.010000  1.605000 20.340000 2.465000 ;
      RECT 20.010000  2.975000 20.340000 3.835000 ;
      RECT 20.090000  0.280000 20.340000 0.825000 ;
      RECT 20.090000  4.615000 20.340000 5.160000 ;
      RECT 20.170000  0.825000 20.340000 1.065000 ;
      RECT 20.170000  1.065000 21.355000 1.395000 ;
      RECT 20.170000  1.395000 20.340000 1.605000 ;
      RECT 20.170000  3.835000 20.340000 4.045000 ;
      RECT 20.170000  4.045000 21.355000 4.375000 ;
      RECT 20.170000  4.375000 20.340000 4.615000 ;
      RECT 20.510000  0.085000 20.800000 0.610000 ;
      RECT 20.510000  4.830000 20.800000 5.355000 ;
      RECT 20.535000  1.605000 20.810000 2.635000 ;
      RECT 20.535000  2.805000 20.810000 3.835000 ;
      RECT 21.055000  1.565000 21.355000 2.465000 ;
      RECT 21.055000  2.975000 21.355000 3.875000 ;
      RECT 21.305000  0.255000 23.335000 0.425000 ;
      RECT 21.305000  0.425000 21.555000 0.770000 ;
      RECT 21.305000  4.670000 21.555000 5.015000 ;
      RECT 21.305000  5.015000 23.335000 5.185000 ;
      RECT 21.525000  1.065000 22.795000 1.365000 ;
      RECT 21.525000  1.365000 21.855000 4.075000 ;
      RECT 21.525000  4.075000 22.795000 4.375000 ;
      RECT 21.725000  0.595000 22.055000 1.065000 ;
      RECT 21.725000  4.375000 22.055000 4.845000 ;
      RECT 22.025000  1.535000 22.295000 2.465000 ;
      RECT 22.025000  2.975000 22.295000 3.905000 ;
      RECT 22.225000  0.425000 22.395000 0.770000 ;
      RECT 22.225000  4.670000 22.395000 5.015000 ;
      RECT 22.465000  1.365000 22.795000 4.075000 ;
      RECT 22.565000  0.595000 22.895000 0.885000 ;
      RECT 22.565000  0.885000 22.795000 1.065000 ;
      RECT 22.565000  4.375000 22.795000 4.555000 ;
      RECT 22.565000  4.555000 22.895000 4.845000 ;
      RECT 22.965000  1.495000 25.195000 1.665000 ;
      RECT 22.965000  1.665000 23.265000 2.465000 ;
      RECT 22.965000  2.635000 29.015000 2.805000 ;
      RECT 22.965000  2.975000 23.265000 3.775000 ;
      RECT 22.965000  3.775000 25.195000 3.945000 ;
      RECT 23.065000  0.425000 23.335000 0.715000 ;
      RECT 23.065000  0.715000 25.195000 0.885000 ;
      RECT 23.065000  4.555000 25.195000 4.725000 ;
      RECT 23.065000  4.725000 23.335000 5.015000 ;
      RECT 23.485000  1.835000 23.755000 2.635000 ;
      RECT 23.485000  2.805000 23.755000 3.605000 ;
      RECT 23.505000  0.085000 23.755000 0.545000 ;
      RECT 23.505000  4.895000 23.755000 5.355000 ;
      RECT 23.925000  0.255000 24.255000 0.715000 ;
      RECT 23.925000  1.665000 24.255000 2.465000 ;
      RECT 23.925000  2.975000 24.255000 3.775000 ;
      RECT 23.925000  4.725000 24.255000 5.185000 ;
      RECT 24.425000  0.085000 24.695000 0.545000 ;
      RECT 24.425000  1.835000 24.695000 2.635000 ;
      RECT 24.425000  2.805000 24.695000 3.605000 ;
      RECT 24.425000  4.895000 24.695000 5.355000 ;
      RECT 24.865000  0.255000 25.195000 0.715000 ;
      RECT 24.865000  1.665000 25.195000 2.465000 ;
      RECT 24.865000  2.975000 25.195000 3.775000 ;
      RECT 24.865000  4.725000 25.195000 5.185000 ;
      RECT 25.365000  0.085000 25.615000 0.885000 ;
      RECT 25.365000  1.495000 25.635000 2.635000 ;
      RECT 25.365000  2.805000 25.635000 3.945000 ;
      RECT 25.365000  4.555000 25.615000 5.355000 ;
      RECT 26.345000  1.495000 26.615000 2.635000 ;
      RECT 26.345000  2.805000 26.615000 3.945000 ;
      RECT 26.365000  0.085000 26.615000 0.885000 ;
      RECT 26.365000  4.555000 26.615000 5.355000 ;
      RECT 26.785000  0.255000 27.115000 0.715000 ;
      RECT 26.785000  0.715000 28.915000 0.885000 ;
      RECT 26.785000  1.495000 29.015000 1.665000 ;
      RECT 26.785000  1.665000 27.115000 2.465000 ;
      RECT 26.785000  2.975000 27.115000 3.775000 ;
      RECT 26.785000  3.775000 29.015000 3.945000 ;
      RECT 26.785000  4.555000 28.915000 4.725000 ;
      RECT 26.785000  4.725000 27.115000 5.185000 ;
      RECT 27.285000  0.085000 27.555000 0.545000 ;
      RECT 27.285000  1.835000 27.555000 2.635000 ;
      RECT 27.285000  2.805000 27.555000 3.605000 ;
      RECT 27.285000  4.895000 27.555000 5.355000 ;
      RECT 27.725000  0.255000 28.055000 0.715000 ;
      RECT 27.725000  1.665000 28.055000 2.465000 ;
      RECT 27.725000  2.975000 28.055000 3.775000 ;
      RECT 27.725000  4.725000 28.055000 5.185000 ;
      RECT 28.225000  0.085000 28.475000 0.545000 ;
      RECT 28.225000  1.835000 28.495000 2.635000 ;
      RECT 28.225000  2.805000 28.495000 3.605000 ;
      RECT 28.225000  4.895000 28.475000 5.355000 ;
      RECT 28.645000  0.255000 30.675000 0.425000 ;
      RECT 28.645000  0.425000 28.915000 0.715000 ;
      RECT 28.645000  4.725000 28.915000 5.015000 ;
      RECT 28.645000  5.015000 30.675000 5.185000 ;
      RECT 28.715000  1.665000 29.015000 2.465000 ;
      RECT 28.715000  2.975000 29.015000 3.775000 ;
      RECT 29.085000  0.595000 29.415000 0.885000 ;
      RECT 29.085000  4.555000 29.415000 4.845000 ;
      RECT 29.185000  0.885000 29.415000 1.065000 ;
      RECT 29.185000  1.065000 30.455000 1.365000 ;
      RECT 29.185000  1.365000 29.515000 4.075000 ;
      RECT 29.185000  4.075000 30.455000 4.375000 ;
      RECT 29.185000  4.375000 29.415000 4.555000 ;
      RECT 29.585000  0.425000 29.755000 0.770000 ;
      RECT 29.585000  4.670000 29.755000 5.015000 ;
      RECT 29.685000  1.535000 29.955000 2.465000 ;
      RECT 29.685000  2.975000 29.955000 3.905000 ;
      RECT 29.925000  0.595000 30.255000 1.065000 ;
      RECT 29.925000  4.375000 30.255000 4.845000 ;
      RECT 30.125000  1.365000 30.455000 4.075000 ;
      RECT 30.425000  0.425000 30.675000 0.770000 ;
      RECT 30.425000  4.670000 30.675000 5.015000 ;
      RECT 30.625000  1.065000 31.810000 1.395000 ;
      RECT 30.625000  1.565000 30.925000 2.465000 ;
      RECT 30.625000  2.635000 34.695000 2.805000 ;
      RECT 30.625000  2.975000 30.925000 3.875000 ;
      RECT 30.625000  4.045000 31.810000 4.375000 ;
      RECT 31.170000  1.605000 31.445000 2.635000 ;
      RECT 31.170000  2.805000 31.445000 3.835000 ;
      RECT 31.180000  0.085000 31.470000 0.610000 ;
      RECT 31.180000  4.830000 31.470000 5.355000 ;
      RECT 31.640000  0.280000 31.890000 0.825000 ;
      RECT 31.640000  0.825000 31.810000 1.065000 ;
      RECT 31.640000  1.395000 31.810000 1.605000 ;
      RECT 31.640000  1.605000 31.970000 2.465000 ;
      RECT 31.640000  2.975000 31.970000 3.835000 ;
      RECT 31.640000  3.835000 31.810000 4.045000 ;
      RECT 31.640000  4.375000 31.810000 4.615000 ;
      RECT 31.640000  4.615000 31.890000 5.160000 ;
      RECT 32.100000  0.085000 32.390000 0.610000 ;
      RECT 32.100000  4.830000 32.390000 5.355000 ;
      RECT 32.140000  1.605000 32.440000 2.635000 ;
      RECT 32.140000  2.805000 32.440000 3.835000 ;
      RECT 32.880000  1.605000 33.180000 2.635000 ;
      RECT 32.880000  2.805000 33.180000 3.835000 ;
      RECT 32.930000  0.085000 33.220000 0.610000 ;
      RECT 32.930000  4.830000 33.220000 5.355000 ;
      RECT 33.350000  1.605000 33.680000 2.465000 ;
      RECT 33.350000  2.975000 33.680000 3.835000 ;
      RECT 33.430000  0.280000 33.680000 0.825000 ;
      RECT 33.430000  4.615000 33.680000 5.160000 ;
      RECT 33.510000  0.825000 33.680000 1.065000 ;
      RECT 33.510000  1.065000 34.695000 1.395000 ;
      RECT 33.510000  1.395000 33.680000 1.605000 ;
      RECT 33.510000  3.835000 33.680000 4.045000 ;
      RECT 33.510000  4.045000 34.695000 4.375000 ;
      RECT 33.510000  4.375000 33.680000 4.615000 ;
      RECT 33.850000  0.085000 34.140000 0.610000 ;
      RECT 33.850000  4.830000 34.140000 5.355000 ;
      RECT 33.875000  1.605000 34.150000 2.635000 ;
      RECT 33.875000  2.805000 34.150000 3.835000 ;
      RECT 34.395000  1.565000 34.695000 2.465000 ;
      RECT 34.395000  2.975000 34.695000 3.875000 ;
      RECT 34.645000  0.255000 36.675000 0.425000 ;
      RECT 34.645000  0.425000 34.895000 0.770000 ;
      RECT 34.645000  4.670000 34.895000 5.015000 ;
      RECT 34.645000  5.015000 36.675000 5.185000 ;
      RECT 34.865000  1.065000 36.135000 1.365000 ;
      RECT 34.865000  1.365000 35.195000 4.075000 ;
      RECT 34.865000  4.075000 36.135000 4.375000 ;
      RECT 35.065000  0.595000 35.395000 1.065000 ;
      RECT 35.065000  4.375000 35.395000 4.845000 ;
      RECT 35.365000  1.535000 35.635000 2.465000 ;
      RECT 35.365000  2.975000 35.635000 3.905000 ;
      RECT 35.565000  0.425000 35.735000 0.770000 ;
      RECT 35.565000  4.670000 35.735000 5.015000 ;
      RECT 35.805000  1.365000 36.135000 4.075000 ;
      RECT 35.905000  0.595000 36.235000 0.885000 ;
      RECT 35.905000  0.885000 36.135000 1.065000 ;
      RECT 35.905000  4.375000 36.135000 4.555000 ;
      RECT 35.905000  4.555000 36.235000 4.845000 ;
      RECT 36.305000  1.495000 38.535000 1.665000 ;
      RECT 36.305000  1.665000 36.605000 2.465000 ;
      RECT 36.305000  2.635000 41.895000 2.805000 ;
      RECT 36.305000  2.975000 36.605000 3.775000 ;
      RECT 36.305000  3.775000 38.535000 3.945000 ;
      RECT 36.405000  0.425000 36.675000 0.715000 ;
      RECT 36.405000  0.715000 38.535000 0.885000 ;
      RECT 36.405000  4.555000 38.535000 4.725000 ;
      RECT 36.405000  4.725000 36.675000 5.015000 ;
      RECT 36.825000  1.835000 37.095000 2.635000 ;
      RECT 36.825000  2.805000 37.095000 3.605000 ;
      RECT 36.845000  0.085000 37.095000 0.545000 ;
      RECT 36.845000  4.895000 37.095000 5.355000 ;
      RECT 37.265000  0.255000 37.595000 0.715000 ;
      RECT 37.265000  1.665000 37.595000 2.465000 ;
      RECT 37.265000  2.975000 37.595000 3.775000 ;
      RECT 37.265000  4.725000 37.595000 5.185000 ;
      RECT 37.765000  0.085000 38.035000 0.545000 ;
      RECT 37.765000  1.835000 38.035000 2.635000 ;
      RECT 37.765000  2.805000 38.035000 3.605000 ;
      RECT 37.765000  4.895000 38.035000 5.355000 ;
      RECT 38.205000  0.255000 38.535000 0.715000 ;
      RECT 38.205000  1.665000 38.535000 2.465000 ;
      RECT 38.205000  2.975000 38.535000 3.775000 ;
      RECT 38.205000  4.725000 38.535000 5.185000 ;
      RECT 38.705000  0.085000 38.955000 0.885000 ;
      RECT 38.705000  1.495000 38.975000 2.635000 ;
      RECT 38.705000  2.805000 38.975000 3.945000 ;
      RECT 38.705000  4.555000 38.955000 5.355000 ;
      RECT 39.225000  1.495000 39.495000 2.635000 ;
      RECT 39.225000  2.805000 39.495000 3.945000 ;
      RECT 39.245000  0.085000 39.495000 0.885000 ;
      RECT 39.245000  4.555000 39.495000 5.355000 ;
      RECT 39.665000  0.255000 39.995000 0.715000 ;
      RECT 39.665000  0.715000 41.795000 0.885000 ;
      RECT 39.665000  1.495000 41.895000 1.665000 ;
      RECT 39.665000  1.665000 39.995000 2.465000 ;
      RECT 39.665000  2.975000 39.995000 3.775000 ;
      RECT 39.665000  3.775000 41.895000 3.945000 ;
      RECT 39.665000  4.555000 41.795000 4.725000 ;
      RECT 39.665000  4.725000 39.995000 5.185000 ;
      RECT 40.165000  0.085000 40.435000 0.545000 ;
      RECT 40.165000  1.835000 40.435000 2.635000 ;
      RECT 40.165000  2.805000 40.435000 3.605000 ;
      RECT 40.165000  4.895000 40.435000 5.355000 ;
      RECT 40.605000  0.255000 40.935000 0.715000 ;
      RECT 40.605000  1.665000 40.935000 2.465000 ;
      RECT 40.605000  2.975000 40.935000 3.775000 ;
      RECT 40.605000  4.725000 40.935000 5.185000 ;
      RECT 41.105000  0.085000 41.355000 0.545000 ;
      RECT 41.105000  1.835000 41.375000 2.635000 ;
      RECT 41.105000  2.805000 41.375000 3.605000 ;
      RECT 41.105000  4.895000 41.355000 5.355000 ;
      RECT 41.525000  0.255000 43.555000 0.425000 ;
      RECT 41.525000  0.425000 41.795000 0.715000 ;
      RECT 41.525000  4.725000 41.795000 5.015000 ;
      RECT 41.525000  5.015000 43.555000 5.185000 ;
      RECT 41.595000  1.665000 41.895000 2.465000 ;
      RECT 41.595000  2.975000 41.895000 3.775000 ;
      RECT 41.965000  0.595000 42.295000 0.885000 ;
      RECT 41.965000  4.555000 42.295000 4.845000 ;
      RECT 42.065000  0.885000 42.295000 1.065000 ;
      RECT 42.065000  1.065000 43.335000 1.365000 ;
      RECT 42.065000  1.365000 42.395000 4.075000 ;
      RECT 42.065000  4.075000 43.335000 4.375000 ;
      RECT 42.065000  4.375000 42.295000 4.555000 ;
      RECT 42.465000  0.425000 42.635000 0.770000 ;
      RECT 42.465000  4.670000 42.635000 5.015000 ;
      RECT 42.565000  1.535000 42.835000 2.465000 ;
      RECT 42.565000  2.975000 42.835000 3.905000 ;
      RECT 42.805000  0.595000 43.135000 1.065000 ;
      RECT 42.805000  4.375000 43.135000 4.845000 ;
      RECT 43.005000  1.365000 43.335000 4.075000 ;
      RECT 43.305000  0.425000 43.555000 0.770000 ;
      RECT 43.305000  4.670000 43.555000 5.015000 ;
      RECT 43.505000  1.065000 44.690000 1.395000 ;
      RECT 43.505000  1.565000 43.805000 2.465000 ;
      RECT 43.505000  2.635000 47.575000 2.805000 ;
      RECT 43.505000  2.975000 43.805000 3.875000 ;
      RECT 43.505000  4.045000 44.690000 4.375000 ;
      RECT 44.050000  1.605000 44.325000 2.635000 ;
      RECT 44.050000  2.805000 44.325000 3.835000 ;
      RECT 44.060000  0.085000 44.350000 0.610000 ;
      RECT 44.060000  4.830000 44.350000 5.355000 ;
      RECT 44.520000  0.280000 44.770000 0.825000 ;
      RECT 44.520000  0.825000 44.690000 1.065000 ;
      RECT 44.520000  1.395000 44.690000 1.605000 ;
      RECT 44.520000  1.605000 44.850000 2.465000 ;
      RECT 44.520000  2.975000 44.850000 3.835000 ;
      RECT 44.520000  3.835000 44.690000 4.045000 ;
      RECT 44.520000  4.375000 44.690000 4.615000 ;
      RECT 44.520000  4.615000 44.770000 5.160000 ;
      RECT 44.980000  0.085000 45.270000 0.610000 ;
      RECT 44.980000  4.830000 45.270000 5.355000 ;
      RECT 45.020000  1.605000 45.320000 2.635000 ;
      RECT 45.020000  2.805000 45.320000 3.835000 ;
      RECT 45.760000  1.605000 46.060000 2.635000 ;
      RECT 45.760000  2.805000 46.060000 3.835000 ;
      RECT 45.810000  0.085000 46.100000 0.610000 ;
      RECT 45.810000  4.830000 46.100000 5.355000 ;
      RECT 46.230000  1.605000 46.560000 2.465000 ;
      RECT 46.230000  2.975000 46.560000 3.835000 ;
      RECT 46.310000  0.280000 46.560000 0.825000 ;
      RECT 46.310000  4.615000 46.560000 5.160000 ;
      RECT 46.390000  0.825000 46.560000 1.065000 ;
      RECT 46.390000  1.065000 47.575000 1.395000 ;
      RECT 46.390000  1.395000 46.560000 1.605000 ;
      RECT 46.390000  3.835000 46.560000 4.045000 ;
      RECT 46.390000  4.045000 47.575000 4.375000 ;
      RECT 46.390000  4.375000 46.560000 4.615000 ;
      RECT 46.730000  0.085000 47.020000 0.610000 ;
      RECT 46.730000  4.830000 47.020000 5.355000 ;
      RECT 46.755000  1.605000 47.030000 2.635000 ;
      RECT 46.755000  2.805000 47.030000 3.835000 ;
      RECT 47.275000  1.565000 47.575000 2.465000 ;
      RECT 47.275000  2.975000 47.575000 3.875000 ;
      RECT 47.525000  0.255000 49.555000 0.425000 ;
      RECT 47.525000  0.425000 47.775000 0.770000 ;
      RECT 47.525000  4.670000 47.775000 5.015000 ;
      RECT 47.525000  5.015000 49.555000 5.185000 ;
      RECT 47.745000  1.065000 49.015000 1.365000 ;
      RECT 47.745000  1.365000 48.075000 4.075000 ;
      RECT 47.745000  4.075000 49.015000 4.375000 ;
      RECT 47.945000  0.595000 48.275000 1.065000 ;
      RECT 47.945000  4.375000 48.275000 4.845000 ;
      RECT 48.245000  1.535000 48.515000 2.465000 ;
      RECT 48.245000  2.975000 48.515000 3.905000 ;
      RECT 48.445000  0.425000 48.615000 0.770000 ;
      RECT 48.445000  4.670000 48.615000 5.015000 ;
      RECT 48.685000  1.365000 49.015000 4.075000 ;
      RECT 48.785000  0.595000 49.115000 0.885000 ;
      RECT 48.785000  0.885000 49.015000 1.065000 ;
      RECT 48.785000  4.375000 49.015000 4.555000 ;
      RECT 48.785000  4.555000 49.115000 4.845000 ;
      RECT 49.185000  1.495000 51.415000 1.665000 ;
      RECT 49.185000  1.665000 49.485000 2.465000 ;
      RECT 49.185000  2.635000 51.980000 2.805000 ;
      RECT 49.185000  2.975000 49.485000 3.775000 ;
      RECT 49.185000  3.775000 51.415000 3.945000 ;
      RECT 49.285000  0.425000 49.555000 0.715000 ;
      RECT 49.285000  0.715000 51.415000 0.885000 ;
      RECT 49.285000  4.555000 51.415000 4.725000 ;
      RECT 49.285000  4.725000 49.555000 5.015000 ;
      RECT 49.705000  1.835000 49.975000 2.635000 ;
      RECT 49.705000  2.805000 49.975000 3.605000 ;
      RECT 49.725000  0.085000 49.975000 0.545000 ;
      RECT 49.725000  4.895000 49.975000 5.355000 ;
      RECT 50.145000  0.255000 50.475000 0.715000 ;
      RECT 50.145000  1.665000 50.475000 2.465000 ;
      RECT 50.145000  2.975000 50.475000 3.775000 ;
      RECT 50.145000  4.725000 50.475000 5.185000 ;
      RECT 50.645000  0.085000 50.915000 0.545000 ;
      RECT 50.645000  1.835000 50.915000 2.635000 ;
      RECT 50.645000  2.805000 50.915000 3.605000 ;
      RECT 50.645000  4.895000 50.915000 5.355000 ;
      RECT 51.085000  0.255000 51.415000 0.715000 ;
      RECT 51.085000  1.665000 51.415000 2.465000 ;
      RECT 51.085000  2.975000 51.415000 3.775000 ;
      RECT 51.085000  4.725000 51.415000 5.185000 ;
      RECT 51.585000  0.085000 51.835000 0.885000 ;
      RECT 51.585000  1.495000 51.855000 2.635000 ;
      RECT 51.585000  2.805000 51.855000 3.945000 ;
      RECT 51.585000  4.555000 51.835000 5.355000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.145000  5.355000  0.315000 5.525000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.605000  5.355000  0.775000 5.525000 ;
      RECT  0.645000  2.140000  0.815000 2.310000 ;
      RECT  0.645000  3.130000  0.815000 3.300000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.065000  5.355000  1.235000 5.525000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.525000  5.355000  1.695000 5.525000 ;
      RECT  1.585000  2.140000  1.755000 2.310000 ;
      RECT  1.585000  3.130000  1.755000 3.300000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  1.985000  5.355000  2.155000 5.525000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.445000  5.355000  2.615000 5.525000 ;
      RECT  2.565000  2.140000  2.735000 2.310000 ;
      RECT  2.565000  3.130000  2.735000 3.300000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  5.355000  3.075000 5.525000 ;
      RECT  3.045000  1.785000  3.215000 1.955000 ;
      RECT  3.045000  3.485000  3.215000 3.655000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  5.355000  3.535000 5.525000 ;
      RECT  3.515000  2.140000  3.685000 2.310000 ;
      RECT  3.515000  3.130000  3.685000 3.300000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  5.355000  3.995000 5.525000 ;
      RECT  3.985000  1.785000  4.155000 1.955000 ;
      RECT  3.985000  3.485000  4.155000 3.655000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  5.355000  4.455000 5.525000 ;
      RECT  4.465000  2.140000  4.635000 2.310000 ;
      RECT  4.465000  3.130000  4.635000 3.300000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.745000  5.355000  4.915000 5.525000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.205000  5.355000  5.375000 5.525000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.665000  5.355000  5.835000 5.525000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.125000  5.355000  6.295000 5.525000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.585000  5.355000  6.755000 5.525000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.045000  5.355000  7.215000 5.525000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.505000  5.355000  7.675000 5.525000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  7.965000  5.355000  8.135000 5.525000 ;
      RECT  8.245000  2.140000  8.415000 2.310000 ;
      RECT  8.245000  3.130000  8.415000 3.300000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  5.355000  8.595000 5.525000 ;
      RECT  8.725000  1.785000  8.895000 1.955000 ;
      RECT  8.725000  3.485000  8.895000 3.655000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  5.355000  9.055000 5.525000 ;
      RECT  9.195000  2.140000  9.365000 2.310000 ;
      RECT  9.195000  3.130000  9.365000 3.300000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  5.355000  9.515000 5.525000 ;
      RECT  9.665000  1.785000  9.835000 1.955000 ;
      RECT  9.665000  3.485000  9.835000 3.655000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  5.355000  9.975000 5.525000 ;
      RECT 10.145000  2.140000 10.315000 2.310000 ;
      RECT 10.145000  3.130000 10.315000 3.300000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.265000  5.355000 10.435000 5.525000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.725000  5.355000 10.895000 5.525000 ;
      RECT 11.125000  2.140000 11.295000 2.310000 ;
      RECT 11.125000  3.130000 11.295000 3.300000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.185000  5.355000 11.355000 5.525000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 11.645000  5.355000 11.815000 5.525000 ;
      RECT 12.065000  2.140000 12.235000 2.310000 ;
      RECT 12.065000  3.130000 12.235000 3.300000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.105000  5.355000 12.275000 5.525000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 12.565000  5.355000 12.735000 5.525000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.025000  5.355000 13.195000 5.525000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.485000  5.355000 13.655000 5.525000 ;
      RECT 13.525000  2.140000 13.695000 2.310000 ;
      RECT 13.525000  3.130000 13.695000 3.300000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 13.945000  5.355000 14.115000 5.525000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.405000  5.355000 14.575000 5.525000 ;
      RECT 14.465000  2.140000 14.635000 2.310000 ;
      RECT 14.465000  3.130000 14.635000 3.300000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 14.865000  5.355000 15.035000 5.525000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.325000  5.355000 15.495000 5.525000 ;
      RECT 15.445000  2.140000 15.615000 2.310000 ;
      RECT 15.445000  3.130000 15.615000 3.300000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  5.355000 15.955000 5.525000 ;
      RECT 15.925000  1.785000 16.095000 1.955000 ;
      RECT 15.925000  3.485000 16.095000 3.655000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  5.355000 16.415000 5.525000 ;
      RECT 16.395000  2.140000 16.565000 2.310000 ;
      RECT 16.395000  3.130000 16.565000 3.300000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  5.355000 16.875000 5.525000 ;
      RECT 16.865000  1.785000 17.035000 1.955000 ;
      RECT 16.865000  3.485000 17.035000 3.655000 ;
      RECT 17.165000 -0.085000 17.335000 0.085000 ;
      RECT 17.165000  5.355000 17.335000 5.525000 ;
      RECT 17.345000  2.140000 17.515000 2.310000 ;
      RECT 17.345000  3.130000 17.515000 3.300000 ;
      RECT 17.625000 -0.085000 17.795000 0.085000 ;
      RECT 17.625000  2.635000 17.795000 2.805000 ;
      RECT 17.625000  5.355000 17.795000 5.525000 ;
      RECT 18.085000 -0.085000 18.255000 0.085000 ;
      RECT 18.085000  2.635000 18.255000 2.805000 ;
      RECT 18.085000  5.355000 18.255000 5.525000 ;
      RECT 18.545000 -0.085000 18.715000 0.085000 ;
      RECT 18.545000  2.635000 18.715000 2.805000 ;
      RECT 18.545000  5.355000 18.715000 5.525000 ;
      RECT 19.005000 -0.085000 19.175000 0.085000 ;
      RECT 19.005000  2.635000 19.175000 2.805000 ;
      RECT 19.005000  5.355000 19.175000 5.525000 ;
      RECT 19.465000 -0.085000 19.635000 0.085000 ;
      RECT 19.465000  2.635000 19.635000 2.805000 ;
      RECT 19.465000  5.355000 19.635000 5.525000 ;
      RECT 19.925000 -0.085000 20.095000 0.085000 ;
      RECT 19.925000  2.635000 20.095000 2.805000 ;
      RECT 19.925000  5.355000 20.095000 5.525000 ;
      RECT 20.385000 -0.085000 20.555000 0.085000 ;
      RECT 20.385000  2.635000 20.555000 2.805000 ;
      RECT 20.385000  5.355000 20.555000 5.525000 ;
      RECT 20.845000 -0.085000 21.015000 0.085000 ;
      RECT 20.845000  2.635000 21.015000 2.805000 ;
      RECT 20.845000  5.355000 21.015000 5.525000 ;
      RECT 21.125000  2.140000 21.295000 2.310000 ;
      RECT 21.125000  3.130000 21.295000 3.300000 ;
      RECT 21.305000 -0.085000 21.475000 0.085000 ;
      RECT 21.305000  5.355000 21.475000 5.525000 ;
      RECT 21.605000  1.785000 21.775000 1.955000 ;
      RECT 21.605000  3.485000 21.775000 3.655000 ;
      RECT 21.765000 -0.085000 21.935000 0.085000 ;
      RECT 21.765000  5.355000 21.935000 5.525000 ;
      RECT 22.075000  2.140000 22.245000 2.310000 ;
      RECT 22.075000  3.130000 22.245000 3.300000 ;
      RECT 22.225000 -0.085000 22.395000 0.085000 ;
      RECT 22.225000  5.355000 22.395000 5.525000 ;
      RECT 22.545000  1.785000 22.715000 1.955000 ;
      RECT 22.545000  3.485000 22.715000 3.655000 ;
      RECT 22.685000 -0.085000 22.855000 0.085000 ;
      RECT 22.685000  5.355000 22.855000 5.525000 ;
      RECT 23.025000  2.140000 23.195000 2.310000 ;
      RECT 23.025000  3.130000 23.195000 3.300000 ;
      RECT 23.145000 -0.085000 23.315000 0.085000 ;
      RECT 23.145000  2.635000 23.315000 2.805000 ;
      RECT 23.145000  5.355000 23.315000 5.525000 ;
      RECT 23.605000 -0.085000 23.775000 0.085000 ;
      RECT 23.605000  2.635000 23.775000 2.805000 ;
      RECT 23.605000  5.355000 23.775000 5.525000 ;
      RECT 24.005000  2.140000 24.175000 2.310000 ;
      RECT 24.005000  3.130000 24.175000 3.300000 ;
      RECT 24.065000 -0.085000 24.235000 0.085000 ;
      RECT 24.065000  2.635000 24.235000 2.805000 ;
      RECT 24.065000  5.355000 24.235000 5.525000 ;
      RECT 24.525000 -0.085000 24.695000 0.085000 ;
      RECT 24.525000  2.635000 24.695000 2.805000 ;
      RECT 24.525000  5.355000 24.695000 5.525000 ;
      RECT 24.945000  2.140000 25.115000 2.310000 ;
      RECT 24.945000  3.130000 25.115000 3.300000 ;
      RECT 24.985000 -0.085000 25.155000 0.085000 ;
      RECT 24.985000  2.635000 25.155000 2.805000 ;
      RECT 24.985000  5.355000 25.155000 5.525000 ;
      RECT 25.445000 -0.085000 25.615000 0.085000 ;
      RECT 25.445000  2.635000 25.615000 2.805000 ;
      RECT 25.445000  5.355000 25.615000 5.525000 ;
      RECT 25.905000 -0.085000 26.075000 0.085000 ;
      RECT 25.905000  2.635000 26.075000 2.805000 ;
      RECT 25.905000  5.355000 26.075000 5.525000 ;
      RECT 26.365000 -0.085000 26.535000 0.085000 ;
      RECT 26.365000  2.635000 26.535000 2.805000 ;
      RECT 26.365000  5.355000 26.535000 5.525000 ;
      RECT 26.825000 -0.085000 26.995000 0.085000 ;
      RECT 26.825000  2.635000 26.995000 2.805000 ;
      RECT 26.825000  5.355000 26.995000 5.525000 ;
      RECT 26.865000  2.140000 27.035000 2.310000 ;
      RECT 26.865000  3.130000 27.035000 3.300000 ;
      RECT 27.285000 -0.085000 27.455000 0.085000 ;
      RECT 27.285000  2.635000 27.455000 2.805000 ;
      RECT 27.285000  5.355000 27.455000 5.525000 ;
      RECT 27.745000 -0.085000 27.915000 0.085000 ;
      RECT 27.745000  2.635000 27.915000 2.805000 ;
      RECT 27.745000  5.355000 27.915000 5.525000 ;
      RECT 27.805000  2.140000 27.975000 2.310000 ;
      RECT 27.805000  3.130000 27.975000 3.300000 ;
      RECT 28.205000 -0.085000 28.375000 0.085000 ;
      RECT 28.205000  2.635000 28.375000 2.805000 ;
      RECT 28.205000  5.355000 28.375000 5.525000 ;
      RECT 28.665000 -0.085000 28.835000 0.085000 ;
      RECT 28.665000  2.635000 28.835000 2.805000 ;
      RECT 28.665000  5.355000 28.835000 5.525000 ;
      RECT 28.785000  2.140000 28.955000 2.310000 ;
      RECT 28.785000  3.130000 28.955000 3.300000 ;
      RECT 29.125000 -0.085000 29.295000 0.085000 ;
      RECT 29.125000  5.355000 29.295000 5.525000 ;
      RECT 29.265000  1.785000 29.435000 1.955000 ;
      RECT 29.265000  3.485000 29.435000 3.655000 ;
      RECT 29.585000 -0.085000 29.755000 0.085000 ;
      RECT 29.585000  5.355000 29.755000 5.525000 ;
      RECT 29.735000  2.140000 29.905000 2.310000 ;
      RECT 29.735000  3.130000 29.905000 3.300000 ;
      RECT 30.045000 -0.085000 30.215000 0.085000 ;
      RECT 30.045000  5.355000 30.215000 5.525000 ;
      RECT 30.205000  1.785000 30.375000 1.955000 ;
      RECT 30.205000  3.485000 30.375000 3.655000 ;
      RECT 30.505000 -0.085000 30.675000 0.085000 ;
      RECT 30.505000  5.355000 30.675000 5.525000 ;
      RECT 30.685000  2.140000 30.855000 2.310000 ;
      RECT 30.685000  3.130000 30.855000 3.300000 ;
      RECT 30.965000 -0.085000 31.135000 0.085000 ;
      RECT 30.965000  2.635000 31.135000 2.805000 ;
      RECT 30.965000  5.355000 31.135000 5.525000 ;
      RECT 31.425000 -0.085000 31.595000 0.085000 ;
      RECT 31.425000  2.635000 31.595000 2.805000 ;
      RECT 31.425000  5.355000 31.595000 5.525000 ;
      RECT 31.885000 -0.085000 32.055000 0.085000 ;
      RECT 31.885000  2.635000 32.055000 2.805000 ;
      RECT 31.885000  5.355000 32.055000 5.525000 ;
      RECT 32.345000 -0.085000 32.515000 0.085000 ;
      RECT 32.345000  2.635000 32.515000 2.805000 ;
      RECT 32.345000  5.355000 32.515000 5.525000 ;
      RECT 32.805000 -0.085000 32.975000 0.085000 ;
      RECT 32.805000  2.635000 32.975000 2.805000 ;
      RECT 32.805000  5.355000 32.975000 5.525000 ;
      RECT 33.265000 -0.085000 33.435000 0.085000 ;
      RECT 33.265000  2.635000 33.435000 2.805000 ;
      RECT 33.265000  5.355000 33.435000 5.525000 ;
      RECT 33.725000 -0.085000 33.895000 0.085000 ;
      RECT 33.725000  2.635000 33.895000 2.805000 ;
      RECT 33.725000  5.355000 33.895000 5.525000 ;
      RECT 34.185000 -0.085000 34.355000 0.085000 ;
      RECT 34.185000  2.635000 34.355000 2.805000 ;
      RECT 34.185000  5.355000 34.355000 5.525000 ;
      RECT 34.465000  2.140000 34.635000 2.310000 ;
      RECT 34.465000  3.130000 34.635000 3.300000 ;
      RECT 34.645000 -0.085000 34.815000 0.085000 ;
      RECT 34.645000  5.355000 34.815000 5.525000 ;
      RECT 34.945000  1.785000 35.115000 1.955000 ;
      RECT 34.945000  3.485000 35.115000 3.655000 ;
      RECT 35.105000 -0.085000 35.275000 0.085000 ;
      RECT 35.105000  5.355000 35.275000 5.525000 ;
      RECT 35.415000  2.140000 35.585000 2.310000 ;
      RECT 35.415000  3.130000 35.585000 3.300000 ;
      RECT 35.565000 -0.085000 35.735000 0.085000 ;
      RECT 35.565000  5.355000 35.735000 5.525000 ;
      RECT 35.885000  1.785000 36.055000 1.955000 ;
      RECT 35.885000  3.485000 36.055000 3.655000 ;
      RECT 36.025000 -0.085000 36.195000 0.085000 ;
      RECT 36.025000  5.355000 36.195000 5.525000 ;
      RECT 36.365000  2.140000 36.535000 2.310000 ;
      RECT 36.365000  3.130000 36.535000 3.300000 ;
      RECT 36.485000 -0.085000 36.655000 0.085000 ;
      RECT 36.485000  2.635000 36.655000 2.805000 ;
      RECT 36.485000  5.355000 36.655000 5.525000 ;
      RECT 36.945000 -0.085000 37.115000 0.085000 ;
      RECT 36.945000  2.635000 37.115000 2.805000 ;
      RECT 36.945000  5.355000 37.115000 5.525000 ;
      RECT 37.345000  2.140000 37.515000 2.310000 ;
      RECT 37.345000  3.130000 37.515000 3.300000 ;
      RECT 37.405000 -0.085000 37.575000 0.085000 ;
      RECT 37.405000  2.635000 37.575000 2.805000 ;
      RECT 37.405000  5.355000 37.575000 5.525000 ;
      RECT 37.865000 -0.085000 38.035000 0.085000 ;
      RECT 37.865000  2.635000 38.035000 2.805000 ;
      RECT 37.865000  5.355000 38.035000 5.525000 ;
      RECT 38.285000  2.140000 38.455000 2.310000 ;
      RECT 38.285000  3.130000 38.455000 3.300000 ;
      RECT 38.325000 -0.085000 38.495000 0.085000 ;
      RECT 38.325000  2.635000 38.495000 2.805000 ;
      RECT 38.325000  5.355000 38.495000 5.525000 ;
      RECT 38.785000 -0.085000 38.955000 0.085000 ;
      RECT 38.785000  2.635000 38.955000 2.805000 ;
      RECT 38.785000  5.355000 38.955000 5.525000 ;
      RECT 39.245000 -0.085000 39.415000 0.085000 ;
      RECT 39.245000  2.635000 39.415000 2.805000 ;
      RECT 39.245000  5.355000 39.415000 5.525000 ;
      RECT 39.705000 -0.085000 39.875000 0.085000 ;
      RECT 39.705000  2.635000 39.875000 2.805000 ;
      RECT 39.705000  5.355000 39.875000 5.525000 ;
      RECT 39.745000  2.140000 39.915000 2.310000 ;
      RECT 39.745000  3.130000 39.915000 3.300000 ;
      RECT 40.165000 -0.085000 40.335000 0.085000 ;
      RECT 40.165000  2.635000 40.335000 2.805000 ;
      RECT 40.165000  5.355000 40.335000 5.525000 ;
      RECT 40.625000 -0.085000 40.795000 0.085000 ;
      RECT 40.625000  2.635000 40.795000 2.805000 ;
      RECT 40.625000  5.355000 40.795000 5.525000 ;
      RECT 40.685000  2.140000 40.855000 2.310000 ;
      RECT 40.685000  3.130000 40.855000 3.300000 ;
      RECT 41.085000 -0.085000 41.255000 0.085000 ;
      RECT 41.085000  2.635000 41.255000 2.805000 ;
      RECT 41.085000  5.355000 41.255000 5.525000 ;
      RECT 41.545000 -0.085000 41.715000 0.085000 ;
      RECT 41.545000  2.635000 41.715000 2.805000 ;
      RECT 41.545000  5.355000 41.715000 5.525000 ;
      RECT 41.665000  2.140000 41.835000 2.310000 ;
      RECT 41.665000  3.130000 41.835000 3.300000 ;
      RECT 42.005000 -0.085000 42.175000 0.085000 ;
      RECT 42.005000  5.355000 42.175000 5.525000 ;
      RECT 42.145000  1.785000 42.315000 1.955000 ;
      RECT 42.145000  3.485000 42.315000 3.655000 ;
      RECT 42.465000 -0.085000 42.635000 0.085000 ;
      RECT 42.465000  5.355000 42.635000 5.525000 ;
      RECT 42.615000  2.140000 42.785000 2.310000 ;
      RECT 42.615000  3.130000 42.785000 3.300000 ;
      RECT 42.925000 -0.085000 43.095000 0.085000 ;
      RECT 42.925000  5.355000 43.095000 5.525000 ;
      RECT 43.085000  1.785000 43.255000 1.955000 ;
      RECT 43.085000  3.485000 43.255000 3.655000 ;
      RECT 43.385000 -0.085000 43.555000 0.085000 ;
      RECT 43.385000  5.355000 43.555000 5.525000 ;
      RECT 43.565000  2.140000 43.735000 2.310000 ;
      RECT 43.565000  3.130000 43.735000 3.300000 ;
      RECT 43.845000 -0.085000 44.015000 0.085000 ;
      RECT 43.845000  2.635000 44.015000 2.805000 ;
      RECT 43.845000  5.355000 44.015000 5.525000 ;
      RECT 44.305000 -0.085000 44.475000 0.085000 ;
      RECT 44.305000  2.635000 44.475000 2.805000 ;
      RECT 44.305000  5.355000 44.475000 5.525000 ;
      RECT 44.765000 -0.085000 44.935000 0.085000 ;
      RECT 44.765000  2.635000 44.935000 2.805000 ;
      RECT 44.765000  5.355000 44.935000 5.525000 ;
      RECT 45.225000 -0.085000 45.395000 0.085000 ;
      RECT 45.225000  2.635000 45.395000 2.805000 ;
      RECT 45.225000  5.355000 45.395000 5.525000 ;
      RECT 45.685000 -0.085000 45.855000 0.085000 ;
      RECT 45.685000  2.635000 45.855000 2.805000 ;
      RECT 45.685000  5.355000 45.855000 5.525000 ;
      RECT 46.145000 -0.085000 46.315000 0.085000 ;
      RECT 46.145000  2.635000 46.315000 2.805000 ;
      RECT 46.145000  5.355000 46.315000 5.525000 ;
      RECT 46.605000 -0.085000 46.775000 0.085000 ;
      RECT 46.605000  2.635000 46.775000 2.805000 ;
      RECT 46.605000  5.355000 46.775000 5.525000 ;
      RECT 47.065000 -0.085000 47.235000 0.085000 ;
      RECT 47.065000  2.635000 47.235000 2.805000 ;
      RECT 47.065000  5.355000 47.235000 5.525000 ;
      RECT 47.345000  2.140000 47.515000 2.310000 ;
      RECT 47.345000  3.130000 47.515000 3.300000 ;
      RECT 47.525000 -0.085000 47.695000 0.085000 ;
      RECT 47.525000  5.355000 47.695000 5.525000 ;
      RECT 47.825000  1.785000 47.995000 1.955000 ;
      RECT 47.825000  3.485000 47.995000 3.655000 ;
      RECT 47.985000 -0.085000 48.155000 0.085000 ;
      RECT 47.985000  5.355000 48.155000 5.525000 ;
      RECT 48.295000  2.140000 48.465000 2.310000 ;
      RECT 48.295000  3.130000 48.465000 3.300000 ;
      RECT 48.445000 -0.085000 48.615000 0.085000 ;
      RECT 48.445000  5.355000 48.615000 5.525000 ;
      RECT 48.765000  1.785000 48.935000 1.955000 ;
      RECT 48.765000  3.485000 48.935000 3.655000 ;
      RECT 48.905000 -0.085000 49.075000 0.085000 ;
      RECT 48.905000  5.355000 49.075000 5.525000 ;
      RECT 49.245000  2.140000 49.415000 2.310000 ;
      RECT 49.245000  3.130000 49.415000 3.300000 ;
      RECT 49.365000 -0.085000 49.535000 0.085000 ;
      RECT 49.365000  2.635000 49.535000 2.805000 ;
      RECT 49.365000  5.355000 49.535000 5.525000 ;
      RECT 49.825000 -0.085000 49.995000 0.085000 ;
      RECT 49.825000  2.635000 49.995000 2.805000 ;
      RECT 49.825000  5.355000 49.995000 5.525000 ;
      RECT 50.225000  2.140000 50.395000 2.310000 ;
      RECT 50.225000  3.130000 50.395000 3.300000 ;
      RECT 50.285000 -0.085000 50.455000 0.085000 ;
      RECT 50.285000  2.635000 50.455000 2.805000 ;
      RECT 50.285000  5.355000 50.455000 5.525000 ;
      RECT 50.745000 -0.085000 50.915000 0.085000 ;
      RECT 50.745000  2.635000 50.915000 2.805000 ;
      RECT 50.745000  5.355000 50.915000 5.525000 ;
      RECT 51.165000  2.140000 51.335000 2.310000 ;
      RECT 51.165000  3.130000 51.335000 3.300000 ;
      RECT 51.205000 -0.085000 51.375000 0.085000 ;
      RECT 51.205000  2.635000 51.375000 2.805000 ;
      RECT 51.205000  5.355000 51.375000 5.525000 ;
      RECT 51.665000 -0.085000 51.835000 0.085000 ;
      RECT 51.665000  2.635000 51.835000 2.805000 ;
      RECT 51.665000  5.355000 51.835000 5.525000 ;
    LAYER met1 ;
      RECT  0.585000 2.110000  0.875000 2.155000 ;
      RECT  0.585000 2.155000  4.695000 2.295000 ;
      RECT  0.585000 2.295000  0.875000 2.340000 ;
      RECT  0.585000 3.100000  0.875000 3.145000 ;
      RECT  0.585000 3.145000  4.695000 3.285000 ;
      RECT  0.585000 3.285000  0.875000 3.330000 ;
      RECT  1.525000 2.110000  1.815000 2.155000 ;
      RECT  1.525000 2.295000  1.815000 2.340000 ;
      RECT  1.525000 3.100000  1.815000 3.145000 ;
      RECT  1.525000 3.285000  1.815000 3.330000 ;
      RECT  2.505000 2.110000  2.795000 2.155000 ;
      RECT  2.505000 2.295000  2.795000 2.340000 ;
      RECT  2.505000 3.100000  2.795000 3.145000 ;
      RECT  2.505000 3.285000  2.795000 3.330000 ;
      RECT  3.455000 2.110000  3.745000 2.155000 ;
      RECT  3.455000 2.295000  3.745000 2.340000 ;
      RECT  3.455000 3.100000  3.745000 3.145000 ;
      RECT  3.455000 3.285000  3.745000 3.330000 ;
      RECT  4.405000 2.110000  4.695000 2.155000 ;
      RECT  4.405000 2.295000  4.695000 2.340000 ;
      RECT  4.405000 3.100000  4.695000 3.145000 ;
      RECT  4.405000 3.285000  4.695000 3.330000 ;
      RECT  8.185000 2.110000  8.475000 2.155000 ;
      RECT  8.185000 2.155000 12.295000 2.295000 ;
      RECT  8.185000 2.295000  8.475000 2.340000 ;
      RECT  8.185000 3.100000  8.475000 3.145000 ;
      RECT  8.185000 3.145000 12.295000 3.285000 ;
      RECT  8.185000 3.285000  8.475000 3.330000 ;
      RECT  9.135000 2.110000  9.425000 2.155000 ;
      RECT  9.135000 2.295000  9.425000 2.340000 ;
      RECT  9.135000 3.100000  9.425000 3.145000 ;
      RECT  9.135000 3.285000  9.425000 3.330000 ;
      RECT 10.085000 2.110000 10.375000 2.155000 ;
      RECT 10.085000 2.295000 10.375000 2.340000 ;
      RECT 10.085000 3.100000 10.375000 3.145000 ;
      RECT 10.085000 3.285000 10.375000 3.330000 ;
      RECT 11.065000 2.110000 11.355000 2.155000 ;
      RECT 11.065000 2.295000 11.355000 2.340000 ;
      RECT 11.065000 3.100000 11.355000 3.145000 ;
      RECT 11.065000 3.285000 11.355000 3.330000 ;
      RECT 12.005000 2.110000 12.295000 2.155000 ;
      RECT 12.005000 2.295000 12.295000 2.340000 ;
      RECT 12.005000 3.100000 12.295000 3.145000 ;
      RECT 12.005000 3.285000 12.295000 3.330000 ;
      RECT 13.465000 2.110000 13.755000 2.155000 ;
      RECT 13.465000 2.155000 17.575000 2.295000 ;
      RECT 13.465000 2.295000 13.755000 2.340000 ;
      RECT 13.465000 3.100000 13.755000 3.145000 ;
      RECT 13.465000 3.145000 17.575000 3.285000 ;
      RECT 13.465000 3.285000 13.755000 3.330000 ;
      RECT 14.405000 2.110000 14.695000 2.155000 ;
      RECT 14.405000 2.295000 14.695000 2.340000 ;
      RECT 14.405000 3.100000 14.695000 3.145000 ;
      RECT 14.405000 3.285000 14.695000 3.330000 ;
      RECT 15.385000 2.110000 15.675000 2.155000 ;
      RECT 15.385000 2.295000 15.675000 2.340000 ;
      RECT 15.385000 3.100000 15.675000 3.145000 ;
      RECT 15.385000 3.285000 15.675000 3.330000 ;
      RECT 16.335000 2.110000 16.625000 2.155000 ;
      RECT 16.335000 2.295000 16.625000 2.340000 ;
      RECT 16.335000 3.100000 16.625000 3.145000 ;
      RECT 16.335000 3.285000 16.625000 3.330000 ;
      RECT 17.285000 2.110000 17.575000 2.155000 ;
      RECT 17.285000 2.295000 17.575000 2.340000 ;
      RECT 17.285000 3.100000 17.575000 3.145000 ;
      RECT 17.285000 3.285000 17.575000 3.330000 ;
      RECT 21.065000 2.110000 21.355000 2.155000 ;
      RECT 21.065000 2.155000 25.175000 2.295000 ;
      RECT 21.065000 2.295000 21.355000 2.340000 ;
      RECT 21.065000 3.100000 21.355000 3.145000 ;
      RECT 21.065000 3.145000 25.175000 3.285000 ;
      RECT 21.065000 3.285000 21.355000 3.330000 ;
      RECT 22.015000 2.110000 22.305000 2.155000 ;
      RECT 22.015000 2.295000 22.305000 2.340000 ;
      RECT 22.015000 3.100000 22.305000 3.145000 ;
      RECT 22.015000 3.285000 22.305000 3.330000 ;
      RECT 22.965000 2.110000 23.255000 2.155000 ;
      RECT 22.965000 2.295000 23.255000 2.340000 ;
      RECT 22.965000 3.100000 23.255000 3.145000 ;
      RECT 22.965000 3.285000 23.255000 3.330000 ;
      RECT 23.945000 2.110000 24.235000 2.155000 ;
      RECT 23.945000 2.295000 24.235000 2.340000 ;
      RECT 23.945000 3.100000 24.235000 3.145000 ;
      RECT 23.945000 3.285000 24.235000 3.330000 ;
      RECT 24.885000 2.110000 25.175000 2.155000 ;
      RECT 24.885000 2.295000 25.175000 2.340000 ;
      RECT 24.885000 3.100000 25.175000 3.145000 ;
      RECT 24.885000 3.285000 25.175000 3.330000 ;
      RECT 26.805000 2.110000 27.095000 2.155000 ;
      RECT 26.805000 2.155000 30.915000 2.295000 ;
      RECT 26.805000 2.295000 27.095000 2.340000 ;
      RECT 26.805000 3.100000 27.095000 3.145000 ;
      RECT 26.805000 3.145000 30.915000 3.285000 ;
      RECT 26.805000 3.285000 27.095000 3.330000 ;
      RECT 27.745000 2.110000 28.035000 2.155000 ;
      RECT 27.745000 2.295000 28.035000 2.340000 ;
      RECT 27.745000 3.100000 28.035000 3.145000 ;
      RECT 27.745000 3.285000 28.035000 3.330000 ;
      RECT 28.725000 2.110000 29.015000 2.155000 ;
      RECT 28.725000 2.295000 29.015000 2.340000 ;
      RECT 28.725000 3.100000 29.015000 3.145000 ;
      RECT 28.725000 3.285000 29.015000 3.330000 ;
      RECT 29.675000 2.110000 29.965000 2.155000 ;
      RECT 29.675000 2.295000 29.965000 2.340000 ;
      RECT 29.675000 3.100000 29.965000 3.145000 ;
      RECT 29.675000 3.285000 29.965000 3.330000 ;
      RECT 30.625000 2.110000 30.915000 2.155000 ;
      RECT 30.625000 2.295000 30.915000 2.340000 ;
      RECT 30.625000 3.100000 30.915000 3.145000 ;
      RECT 30.625000 3.285000 30.915000 3.330000 ;
      RECT 34.405000 2.110000 34.695000 2.155000 ;
      RECT 34.405000 2.155000 38.515000 2.295000 ;
      RECT 34.405000 2.295000 34.695000 2.340000 ;
      RECT 34.405000 3.100000 34.695000 3.145000 ;
      RECT 34.405000 3.145000 38.515000 3.285000 ;
      RECT 34.405000 3.285000 34.695000 3.330000 ;
      RECT 35.355000 2.110000 35.645000 2.155000 ;
      RECT 35.355000 2.295000 35.645000 2.340000 ;
      RECT 35.355000 3.100000 35.645000 3.145000 ;
      RECT 35.355000 3.285000 35.645000 3.330000 ;
      RECT 36.305000 2.110000 36.595000 2.155000 ;
      RECT 36.305000 2.295000 36.595000 2.340000 ;
      RECT 36.305000 3.100000 36.595000 3.145000 ;
      RECT 36.305000 3.285000 36.595000 3.330000 ;
      RECT 37.285000 2.110000 37.575000 2.155000 ;
      RECT 37.285000 2.295000 37.575000 2.340000 ;
      RECT 37.285000 3.100000 37.575000 3.145000 ;
      RECT 37.285000 3.285000 37.575000 3.330000 ;
      RECT 38.225000 2.110000 38.515000 2.155000 ;
      RECT 38.225000 2.295000 38.515000 2.340000 ;
      RECT 38.225000 3.100000 38.515000 3.145000 ;
      RECT 38.225000 3.285000 38.515000 3.330000 ;
      RECT 39.685000 2.110000 39.975000 2.155000 ;
      RECT 39.685000 2.155000 43.795000 2.295000 ;
      RECT 39.685000 2.295000 39.975000 2.340000 ;
      RECT 39.685000 3.100000 39.975000 3.145000 ;
      RECT 39.685000 3.145000 43.795000 3.285000 ;
      RECT 39.685000 3.285000 39.975000 3.330000 ;
      RECT 40.625000 2.110000 40.915000 2.155000 ;
      RECT 40.625000 2.295000 40.915000 2.340000 ;
      RECT 40.625000 3.100000 40.915000 3.145000 ;
      RECT 40.625000 3.285000 40.915000 3.330000 ;
      RECT 41.605000 2.110000 41.895000 2.155000 ;
      RECT 41.605000 2.295000 41.895000 2.340000 ;
      RECT 41.605000 3.100000 41.895000 3.145000 ;
      RECT 41.605000 3.285000 41.895000 3.330000 ;
      RECT 42.555000 2.110000 42.845000 2.155000 ;
      RECT 42.555000 2.295000 42.845000 2.340000 ;
      RECT 42.555000 3.100000 42.845000 3.145000 ;
      RECT 42.555000 3.285000 42.845000 3.330000 ;
      RECT 43.505000 2.110000 43.795000 2.155000 ;
      RECT 43.505000 2.295000 43.795000 2.340000 ;
      RECT 43.505000 3.100000 43.795000 3.145000 ;
      RECT 43.505000 3.285000 43.795000 3.330000 ;
      RECT 47.285000 2.110000 47.575000 2.155000 ;
      RECT 47.285000 2.155000 51.395000 2.295000 ;
      RECT 47.285000 2.295000 47.575000 2.340000 ;
      RECT 47.285000 3.100000 47.575000 3.145000 ;
      RECT 47.285000 3.145000 51.395000 3.285000 ;
      RECT 47.285000 3.285000 47.575000 3.330000 ;
      RECT 48.235000 2.110000 48.525000 2.155000 ;
      RECT 48.235000 2.295000 48.525000 2.340000 ;
      RECT 48.235000 3.100000 48.525000 3.145000 ;
      RECT 48.235000 3.285000 48.525000 3.330000 ;
      RECT 49.185000 2.110000 49.475000 2.155000 ;
      RECT 49.185000 2.295000 49.475000 2.340000 ;
      RECT 49.185000 3.100000 49.475000 3.145000 ;
      RECT 49.185000 3.285000 49.475000 3.330000 ;
      RECT 50.165000 2.110000 50.455000 2.155000 ;
      RECT 50.165000 2.295000 50.455000 2.340000 ;
      RECT 50.165000 3.100000 50.455000 3.145000 ;
      RECT 50.165000 3.285000 50.455000 3.330000 ;
      RECT 51.105000 2.110000 51.395000 2.155000 ;
      RECT 51.105000 2.295000 51.395000 2.340000 ;
      RECT 51.105000 3.100000 51.395000 3.145000 ;
      RECT 51.105000 3.285000 51.395000 3.330000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb16to1_4


MACRO sky130_fd_sc_hdll__muxb16to1_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  17.02000 BY  5.440000 ;
  SITE unithd ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.335000 1.055000 0.730000 1.325000 ;
        RECT 0.560000 0.395000 0.835000 0.625000 ;
        RECT 0.560000 0.625000 0.730000 1.055000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 0.395000 4.040000 0.625000 ;
        RECT 3.870000 0.625000 4.040000 1.055000 ;
        RECT 3.870000 1.055000 4.265000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 1.055000 4.870000 1.325000 ;
        RECT 4.700000 0.395000 4.975000 0.625000 ;
        RECT 4.700000 0.625000 4.870000 1.055000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.905000 0.395000 8.180000 0.625000 ;
        RECT 8.010000 0.625000 8.180000 1.055000 ;
        RECT 8.010000 1.055000 8.405000 1.325000 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.615000 1.055000 9.010000 1.325000 ;
        RECT 8.840000 0.395000 9.115000 0.625000 ;
        RECT 8.840000 0.625000 9.010000 1.055000 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.045000 0.395000 12.320000 0.625000 ;
        RECT 12.150000 0.625000 12.320000 1.055000 ;
        RECT 12.150000 1.055000 12.545000 1.325000 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755000 1.055000 13.150000 1.325000 ;
        RECT 12.980000 0.395000 13.255000 0.625000 ;
        RECT 12.980000 0.625000 13.150000 1.055000 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.185000 0.395000 16.460000 0.625000 ;
        RECT 16.290000 0.625000 16.460000 1.055000 ;
        RECT 16.290000 1.055000 16.685000 1.325000 ;
    END
  END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.335000 4.115000 0.730000 4.385000 ;
        RECT 0.560000 4.385000 0.730000 4.815000 ;
        RECT 0.560000 4.815000 0.835000 5.045000 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 4.815000 4.040000 5.045000 ;
        RECT 3.870000 4.115000 4.265000 4.385000 ;
        RECT 3.870000 4.385000 4.040000 4.815000 ;
    END
  END D[9]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 4.115000 4.870000 4.385000 ;
        RECT 4.700000 4.385000 4.870000 4.815000 ;
        RECT 4.700000 4.815000 4.975000 5.045000 ;
    END
  END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.905000 4.815000 8.180000 5.045000 ;
        RECT 8.010000 4.115000 8.405000 4.385000 ;
        RECT 8.010000 4.385000 8.180000 4.815000 ;
    END
  END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.615000 4.115000 9.010000 4.385000 ;
        RECT 8.840000 4.385000 9.010000 4.815000 ;
        RECT 8.840000 4.815000 9.115000 5.045000 ;
    END
  END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.045000 4.815000 12.320000 5.045000 ;
        RECT 12.150000 4.115000 12.545000 4.385000 ;
        RECT 12.150000 4.385000 12.320000 4.815000 ;
    END
  END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755000 4.115000 13.150000 4.385000 ;
        RECT 12.980000 4.385000 13.150000 4.815000 ;
        RECT 12.980000 4.815000 13.255000 5.045000 ;
    END
  END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.185000 4.815000 16.460000 5.045000 ;
        RECT 16.290000 4.115000 16.685000 4.385000 ;
        RECT 16.290000 4.385000 16.460000 4.815000 ;
    END
  END D[15]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 0.945000 2.205000 1.295000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.395000 0.945000 2.795000 1.295000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.945000 0.945000 6.345000 1.295000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 0.945000 6.935000 1.295000 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.085000 0.945000 10.485000 1.295000 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.675000 0.945000 11.075000 1.295000 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.225000 0.945000 14.625000 1.295000 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.815000 0.945000 15.215000 1.295000 ;
    END
  END S[7]
  PIN S[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 4.145000 2.205000 4.495000 ;
    END
  END S[8]
  PIN S[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.395000 4.145000 2.795000 4.495000 ;
    END
  END S[9]
  PIN S[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.945000 4.145000 6.345000 4.495000 ;
    END
  END S[10]
  PIN S[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 4.145000 6.935000 4.495000 ;
    END
  END S[11]
  PIN S[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.085000 4.145000 10.485000 4.495000 ;
    END
  END S[12]
  PIN S[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.675000 4.145000 11.075000 4.495000 ;
    END
  END S[13]
  PIN S[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.225000 4.145000 14.625000 4.495000 ;
    END
  END S[14]
  PIN S[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.815000 4.145000 15.215000 4.495000 ;
    END
  END S[15]
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  1.005000 1.755000  1.295000 1.800000 ;
        RECT  1.005000 1.800000 16.015000 1.940000 ;
        RECT  1.005000 1.940000  1.295000 1.985000 ;
        RECT  1.005000 3.455000  1.295000 3.500000 ;
        RECT  1.005000 3.500000 16.015000 3.640000 ;
        RECT  1.005000 3.640000  1.295000 3.685000 ;
        RECT  3.305000 1.755000  3.595000 1.800000 ;
        RECT  3.305000 1.940000  3.595000 1.985000 ;
        RECT  3.305000 3.455000  3.595000 3.500000 ;
        RECT  3.305000 3.640000  3.595000 3.685000 ;
        RECT  5.145000 1.755000  5.435000 1.800000 ;
        RECT  5.145000 1.940000  5.435000 1.985000 ;
        RECT  5.145000 3.455000  5.435000 3.500000 ;
        RECT  5.145000 3.640000  5.435000 3.685000 ;
        RECT  7.445000 1.755000  7.735000 1.800000 ;
        RECT  7.445000 1.940000  7.735000 1.985000 ;
        RECT  7.445000 3.455000  7.735000 3.500000 ;
        RECT  7.445000 3.640000  7.735000 3.685000 ;
        RECT  9.285000 1.755000  9.575000 1.800000 ;
        RECT  9.285000 1.940000  9.575000 1.985000 ;
        RECT  9.285000 3.455000  9.575000 3.500000 ;
        RECT  9.285000 3.640000  9.575000 3.685000 ;
        RECT 11.585000 1.755000 11.875000 1.800000 ;
        RECT 11.585000 1.940000 11.875000 1.985000 ;
        RECT 11.585000 3.455000 11.875000 3.500000 ;
        RECT 11.585000 3.640000 11.875000 3.685000 ;
        RECT 13.425000 1.755000 13.715000 1.800000 ;
        RECT 13.425000 1.940000 13.715000 1.985000 ;
        RECT 13.425000 3.455000 13.715000 3.500000 ;
        RECT 13.425000 3.640000 13.715000 3.685000 ;
        RECT 15.725000 1.755000 16.015000 1.800000 ;
        RECT 15.725000 1.940000 16.015000 1.985000 ;
        RECT 15.725000 3.455000 16.015000 3.500000 ;
        RECT 15.725000 3.640000 16.015000 3.685000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 17.020000 0.240000 ;
        RECT 0.000000  5.200000 17.020000 5.680000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 17.020000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 17.020000 0.085000 ;
      RECT  0.000000  2.635000  0.920000 2.805000 ;
      RECT  0.000000  5.355000 17.020000 5.525000 ;
      RECT  0.095000  1.495000  0.425000 2.635000 ;
      RECT  0.095000  2.805000  0.425000 3.945000 ;
      RECT  0.130000  0.085000  0.390000 0.885000 ;
      RECT  0.130000  4.555000  0.390000 5.355000 ;
      RECT  0.900000  0.835000  1.290000 1.005000 ;
      RECT  0.900000  1.005000  1.070000 1.755000 ;
      RECT  0.900000  1.755000  1.295000 1.805000 ;
      RECT  0.900000  1.805000  1.420000 1.985000 ;
      RECT  0.900000  3.455000  1.420000 3.635000 ;
      RECT  0.900000  3.635000  1.295000 3.685000 ;
      RECT  0.900000  3.685000  1.070000 4.435000 ;
      RECT  0.900000  4.435000  1.290000 4.605000 ;
      RECT  1.045000  0.330000  1.290000 0.835000 ;
      RECT  1.045000  4.605000  1.290000 5.110000 ;
      RECT  1.090000  1.985000  1.420000 2.465000 ;
      RECT  1.090000  2.465000  1.295000 2.975000 ;
      RECT  1.090000  2.975000  1.420000 3.455000 ;
      RECT  1.240000  1.175000  1.630000 1.465000 ;
      RECT  1.240000  1.465000  1.940000 1.505000 ;
      RECT  1.240000  3.935000  1.940000 3.975000 ;
      RECT  1.240000  3.975000  1.630000 4.265000 ;
      RECT  1.460000  0.585000  1.900000 0.755000 ;
      RECT  1.460000  0.755000  1.630000 1.175000 ;
      RECT  1.460000  1.505000  1.940000 1.635000 ;
      RECT  1.460000  3.805000  1.940000 3.935000 ;
      RECT  1.460000  4.265000  1.630000 4.685000 ;
      RECT  1.460000  4.685000  1.900000 4.855000 ;
      RECT  1.465000  2.635000  3.135000 2.805000 ;
      RECT  1.610000  1.635000  1.940000 2.465000 ;
      RECT  1.610000  2.975000  1.940000 3.805000 ;
      RECT  1.650000  0.330000  1.900000 0.585000 ;
      RECT  1.650000  4.855000  1.900000 5.110000 ;
      RECT  2.135000  0.085000  2.465000 0.660000 ;
      RECT  2.135000  1.465000  2.465000 2.635000 ;
      RECT  2.135000  2.805000  2.465000 3.975000 ;
      RECT  2.135000  4.780000  2.465000 5.355000 ;
      RECT  2.660000  1.465000  3.360000 1.505000 ;
      RECT  2.660000  1.505000  3.140000 1.635000 ;
      RECT  2.660000  1.635000  2.990000 2.465000 ;
      RECT  2.660000  2.975000  2.990000 3.805000 ;
      RECT  2.660000  3.805000  3.140000 3.935000 ;
      RECT  2.660000  3.935000  3.360000 3.975000 ;
      RECT  2.700000  0.330000  2.950000 0.585000 ;
      RECT  2.700000  0.585000  3.140000 0.755000 ;
      RECT  2.700000  4.685000  3.140000 4.855000 ;
      RECT  2.700000  4.855000  2.950000 5.110000 ;
      RECT  2.970000  0.755000  3.140000 1.175000 ;
      RECT  2.970000  1.175000  3.360000 1.465000 ;
      RECT  2.970000  3.975000  3.360000 4.265000 ;
      RECT  2.970000  4.265000  3.140000 4.685000 ;
      RECT  3.180000  1.805000  3.700000 1.985000 ;
      RECT  3.180000  1.985000  3.510000 2.465000 ;
      RECT  3.180000  2.975000  3.510000 3.455000 ;
      RECT  3.180000  3.455000  3.700000 3.635000 ;
      RECT  3.305000  1.755000  3.700000 1.805000 ;
      RECT  3.305000  2.465000  3.510000 2.975000 ;
      RECT  3.305000  3.635000  3.700000 3.685000 ;
      RECT  3.310000  0.330000  3.555000 0.835000 ;
      RECT  3.310000  0.835000  3.700000 1.005000 ;
      RECT  3.310000  4.435000  3.700000 4.605000 ;
      RECT  3.310000  4.605000  3.555000 5.110000 ;
      RECT  3.530000  1.005000  3.700000 1.755000 ;
      RECT  3.530000  3.685000  3.700000 4.435000 ;
      RECT  3.680000  2.635000  5.060000 2.805000 ;
      RECT  4.175000  1.495000  4.565000 2.635000 ;
      RECT  4.175000  2.805000  4.565000 3.945000 ;
      RECT  4.210000  0.085000  4.530000 0.885000 ;
      RECT  4.210000  4.555000  4.530000 5.355000 ;
      RECT  5.040000  0.835000  5.430000 1.005000 ;
      RECT  5.040000  1.005000  5.210000 1.755000 ;
      RECT  5.040000  1.755000  5.435000 1.805000 ;
      RECT  5.040000  1.805000  5.560000 1.985000 ;
      RECT  5.040000  3.455000  5.560000 3.635000 ;
      RECT  5.040000  3.635000  5.435000 3.685000 ;
      RECT  5.040000  3.685000  5.210000 4.435000 ;
      RECT  5.040000  4.435000  5.430000 4.605000 ;
      RECT  5.185000  0.330000  5.430000 0.835000 ;
      RECT  5.185000  4.605000  5.430000 5.110000 ;
      RECT  5.230000  1.985000  5.560000 2.465000 ;
      RECT  5.230000  2.465000  5.435000 2.975000 ;
      RECT  5.230000  2.975000  5.560000 3.455000 ;
      RECT  5.380000  1.175000  5.770000 1.465000 ;
      RECT  5.380000  1.465000  6.080000 1.505000 ;
      RECT  5.380000  3.935000  6.080000 3.975000 ;
      RECT  5.380000  3.975000  5.770000 4.265000 ;
      RECT  5.600000  0.585000  6.040000 0.755000 ;
      RECT  5.600000  0.755000  5.770000 1.175000 ;
      RECT  5.600000  1.505000  6.080000 1.635000 ;
      RECT  5.600000  3.805000  6.080000 3.935000 ;
      RECT  5.600000  4.265000  5.770000 4.685000 ;
      RECT  5.600000  4.685000  6.040000 4.855000 ;
      RECT  5.605000  2.635000  7.275000 2.805000 ;
      RECT  5.750000  1.635000  6.080000 2.465000 ;
      RECT  5.750000  2.975000  6.080000 3.805000 ;
      RECT  5.790000  0.330000  6.040000 0.585000 ;
      RECT  5.790000  4.855000  6.040000 5.110000 ;
      RECT  6.275000  0.085000  6.605000 0.660000 ;
      RECT  6.275000  1.465000  6.605000 2.635000 ;
      RECT  6.275000  2.805000  6.605000 3.975000 ;
      RECT  6.275000  4.780000  6.605000 5.355000 ;
      RECT  6.800000  1.465000  7.500000 1.505000 ;
      RECT  6.800000  1.505000  7.280000 1.635000 ;
      RECT  6.800000  1.635000  7.130000 2.465000 ;
      RECT  6.800000  2.975000  7.130000 3.805000 ;
      RECT  6.800000  3.805000  7.280000 3.935000 ;
      RECT  6.800000  3.935000  7.500000 3.975000 ;
      RECT  6.840000  0.330000  7.090000 0.585000 ;
      RECT  6.840000  0.585000  7.280000 0.755000 ;
      RECT  6.840000  4.685000  7.280000 4.855000 ;
      RECT  6.840000  4.855000  7.090000 5.110000 ;
      RECT  7.110000  0.755000  7.280000 1.175000 ;
      RECT  7.110000  1.175000  7.500000 1.465000 ;
      RECT  7.110000  3.975000  7.500000 4.265000 ;
      RECT  7.110000  4.265000  7.280000 4.685000 ;
      RECT  7.320000  1.805000  7.840000 1.985000 ;
      RECT  7.320000  1.985000  7.650000 2.465000 ;
      RECT  7.320000  2.975000  7.650000 3.455000 ;
      RECT  7.320000  3.455000  7.840000 3.635000 ;
      RECT  7.445000  1.755000  7.840000 1.805000 ;
      RECT  7.445000  2.465000  7.650000 2.975000 ;
      RECT  7.445000  3.635000  7.840000 3.685000 ;
      RECT  7.450000  0.330000  7.695000 0.835000 ;
      RECT  7.450000  0.835000  7.840000 1.005000 ;
      RECT  7.450000  4.435000  7.840000 4.605000 ;
      RECT  7.450000  4.605000  7.695000 5.110000 ;
      RECT  7.670000  1.005000  7.840000 1.755000 ;
      RECT  7.670000  3.685000  7.840000 4.435000 ;
      RECT  7.820000  2.635000  9.200000 2.805000 ;
      RECT  8.315000  1.495000  8.705000 2.635000 ;
      RECT  8.315000  2.805000  8.705000 3.945000 ;
      RECT  8.350000  0.085000  8.670000 0.885000 ;
      RECT  8.350000  4.555000  8.670000 5.355000 ;
      RECT  9.180000  0.835000  9.570000 1.005000 ;
      RECT  9.180000  1.005000  9.350000 1.755000 ;
      RECT  9.180000  1.755000  9.575000 1.805000 ;
      RECT  9.180000  1.805000  9.700000 1.985000 ;
      RECT  9.180000  3.455000  9.700000 3.635000 ;
      RECT  9.180000  3.635000  9.575000 3.685000 ;
      RECT  9.180000  3.685000  9.350000 4.435000 ;
      RECT  9.180000  4.435000  9.570000 4.605000 ;
      RECT  9.325000  0.330000  9.570000 0.835000 ;
      RECT  9.325000  4.605000  9.570000 5.110000 ;
      RECT  9.370000  1.985000  9.700000 2.465000 ;
      RECT  9.370000  2.465000  9.575000 2.975000 ;
      RECT  9.370000  2.975000  9.700000 3.455000 ;
      RECT  9.520000  1.175000  9.910000 1.465000 ;
      RECT  9.520000  1.465000 10.220000 1.505000 ;
      RECT  9.520000  3.935000 10.220000 3.975000 ;
      RECT  9.520000  3.975000  9.910000 4.265000 ;
      RECT  9.740000  0.585000 10.180000 0.755000 ;
      RECT  9.740000  0.755000  9.910000 1.175000 ;
      RECT  9.740000  1.505000 10.220000 1.635000 ;
      RECT  9.740000  3.805000 10.220000 3.935000 ;
      RECT  9.740000  4.265000  9.910000 4.685000 ;
      RECT  9.740000  4.685000 10.180000 4.855000 ;
      RECT  9.745000  2.635000 11.415000 2.805000 ;
      RECT  9.890000  1.635000 10.220000 2.465000 ;
      RECT  9.890000  2.975000 10.220000 3.805000 ;
      RECT  9.930000  0.330000 10.180000 0.585000 ;
      RECT  9.930000  4.855000 10.180000 5.110000 ;
      RECT 10.415000  0.085000 10.745000 0.660000 ;
      RECT 10.415000  1.465000 10.745000 2.635000 ;
      RECT 10.415000  2.805000 10.745000 3.975000 ;
      RECT 10.415000  4.780000 10.745000 5.355000 ;
      RECT 10.940000  1.465000 11.640000 1.505000 ;
      RECT 10.940000  1.505000 11.420000 1.635000 ;
      RECT 10.940000  1.635000 11.270000 2.465000 ;
      RECT 10.940000  2.975000 11.270000 3.805000 ;
      RECT 10.940000  3.805000 11.420000 3.935000 ;
      RECT 10.940000  3.935000 11.640000 3.975000 ;
      RECT 10.980000  0.330000 11.230000 0.585000 ;
      RECT 10.980000  0.585000 11.420000 0.755000 ;
      RECT 10.980000  4.685000 11.420000 4.855000 ;
      RECT 10.980000  4.855000 11.230000 5.110000 ;
      RECT 11.250000  0.755000 11.420000 1.175000 ;
      RECT 11.250000  1.175000 11.640000 1.465000 ;
      RECT 11.250000  3.975000 11.640000 4.265000 ;
      RECT 11.250000  4.265000 11.420000 4.685000 ;
      RECT 11.460000  1.805000 11.980000 1.985000 ;
      RECT 11.460000  1.985000 11.790000 2.465000 ;
      RECT 11.460000  2.975000 11.790000 3.455000 ;
      RECT 11.460000  3.455000 11.980000 3.635000 ;
      RECT 11.585000  1.755000 11.980000 1.805000 ;
      RECT 11.585000  2.465000 11.790000 2.975000 ;
      RECT 11.585000  3.635000 11.980000 3.685000 ;
      RECT 11.590000  0.330000 11.835000 0.835000 ;
      RECT 11.590000  0.835000 11.980000 1.005000 ;
      RECT 11.590000  4.435000 11.980000 4.605000 ;
      RECT 11.590000  4.605000 11.835000 5.110000 ;
      RECT 11.810000  1.005000 11.980000 1.755000 ;
      RECT 11.810000  3.685000 11.980000 4.435000 ;
      RECT 11.960000  2.635000 13.340000 2.805000 ;
      RECT 12.455000  1.495000 12.845000 2.635000 ;
      RECT 12.455000  2.805000 12.845000 3.945000 ;
      RECT 12.490000  0.085000 12.810000 0.885000 ;
      RECT 12.490000  4.555000 12.810000 5.355000 ;
      RECT 13.320000  0.835000 13.710000 1.005000 ;
      RECT 13.320000  1.005000 13.490000 1.755000 ;
      RECT 13.320000  1.755000 13.715000 1.805000 ;
      RECT 13.320000  1.805000 13.840000 1.985000 ;
      RECT 13.320000  3.455000 13.840000 3.635000 ;
      RECT 13.320000  3.635000 13.715000 3.685000 ;
      RECT 13.320000  3.685000 13.490000 4.435000 ;
      RECT 13.320000  4.435000 13.710000 4.605000 ;
      RECT 13.465000  0.330000 13.710000 0.835000 ;
      RECT 13.465000  4.605000 13.710000 5.110000 ;
      RECT 13.510000  1.985000 13.840000 2.465000 ;
      RECT 13.510000  2.465000 13.715000 2.975000 ;
      RECT 13.510000  2.975000 13.840000 3.455000 ;
      RECT 13.660000  1.175000 14.050000 1.465000 ;
      RECT 13.660000  1.465000 14.360000 1.505000 ;
      RECT 13.660000  3.935000 14.360000 3.975000 ;
      RECT 13.660000  3.975000 14.050000 4.265000 ;
      RECT 13.880000  0.585000 14.320000 0.755000 ;
      RECT 13.880000  0.755000 14.050000 1.175000 ;
      RECT 13.880000  1.505000 14.360000 1.635000 ;
      RECT 13.880000  3.805000 14.360000 3.935000 ;
      RECT 13.880000  4.265000 14.050000 4.685000 ;
      RECT 13.880000  4.685000 14.320000 4.855000 ;
      RECT 13.885000  2.635000 15.555000 2.805000 ;
      RECT 14.030000  1.635000 14.360000 2.465000 ;
      RECT 14.030000  2.975000 14.360000 3.805000 ;
      RECT 14.070000  0.330000 14.320000 0.585000 ;
      RECT 14.070000  4.855000 14.320000 5.110000 ;
      RECT 14.555000  0.085000 14.885000 0.660000 ;
      RECT 14.555000  1.465000 14.885000 2.635000 ;
      RECT 14.555000  2.805000 14.885000 3.975000 ;
      RECT 14.555000  4.780000 14.885000 5.355000 ;
      RECT 15.080000  1.465000 15.780000 1.505000 ;
      RECT 15.080000  1.505000 15.560000 1.635000 ;
      RECT 15.080000  1.635000 15.410000 2.465000 ;
      RECT 15.080000  2.975000 15.410000 3.805000 ;
      RECT 15.080000  3.805000 15.560000 3.935000 ;
      RECT 15.080000  3.935000 15.780000 3.975000 ;
      RECT 15.120000  0.330000 15.370000 0.585000 ;
      RECT 15.120000  0.585000 15.560000 0.755000 ;
      RECT 15.120000  4.685000 15.560000 4.855000 ;
      RECT 15.120000  4.855000 15.370000 5.110000 ;
      RECT 15.390000  0.755000 15.560000 1.175000 ;
      RECT 15.390000  1.175000 15.780000 1.465000 ;
      RECT 15.390000  3.975000 15.780000 4.265000 ;
      RECT 15.390000  4.265000 15.560000 4.685000 ;
      RECT 15.600000  1.805000 16.120000 1.985000 ;
      RECT 15.600000  1.985000 15.930000 2.465000 ;
      RECT 15.600000  2.975000 15.930000 3.455000 ;
      RECT 15.600000  3.455000 16.120000 3.635000 ;
      RECT 15.725000  1.755000 16.120000 1.805000 ;
      RECT 15.725000  2.465000 15.930000 2.975000 ;
      RECT 15.725000  3.635000 16.120000 3.685000 ;
      RECT 15.730000  0.330000 15.975000 0.835000 ;
      RECT 15.730000  0.835000 16.120000 1.005000 ;
      RECT 15.730000  4.435000 16.120000 4.605000 ;
      RECT 15.730000  4.605000 15.975000 5.110000 ;
      RECT 15.950000  1.005000 16.120000 1.755000 ;
      RECT 15.950000  3.685000 16.120000 4.435000 ;
      RECT 16.100000  2.635000 17.020000 2.805000 ;
      RECT 16.595000  1.495000 16.925000 2.635000 ;
      RECT 16.595000  2.805000 16.925000 3.945000 ;
      RECT 16.630000  0.085000 16.890000 0.885000 ;
      RECT 16.630000  4.555000 16.890000 5.355000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.145000  5.355000  0.315000 5.525000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.605000  5.355000  0.775000 5.525000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  1.785000  1.235000 1.955000 ;
      RECT  1.065000  3.485000  1.235000 3.655000 ;
      RECT  1.065000  5.355000  1.235000 5.525000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.525000  5.355000  1.695000 5.525000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  1.985000  5.355000  2.155000 5.525000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.445000  5.355000  2.615000 5.525000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  2.905000  5.355000  3.075000 5.525000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  1.785000  3.535000 1.955000 ;
      RECT  3.365000  3.485000  3.535000 3.655000 ;
      RECT  3.365000  5.355000  3.535000 5.525000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  3.825000  5.355000  3.995000 5.525000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.285000  5.355000  4.455000 5.525000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.745000  5.355000  4.915000 5.525000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  3.485000  5.375000 3.655000 ;
      RECT  5.205000  5.355000  5.375000 5.525000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.665000  5.355000  5.835000 5.525000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.125000  5.355000  6.295000 5.525000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.585000  5.355000  6.755000 5.525000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.045000  5.355000  7.215000 5.525000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  1.785000  7.675000 1.955000 ;
      RECT  7.505000  3.485000  7.675000 3.655000 ;
      RECT  7.505000  5.355000  7.675000 5.525000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  7.965000  5.355000  8.135000 5.525000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.425000  5.355000  8.595000 5.525000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.885000  5.355000  9.055000 5.525000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  1.785000  9.515000 1.955000 ;
      RECT  9.345000  3.485000  9.515000 3.655000 ;
      RECT  9.345000  5.355000  9.515000 5.525000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT  9.805000  5.355000  9.975000 5.525000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.265000  5.355000 10.435000 5.525000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.725000  5.355000 10.895000 5.525000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.185000  5.355000 11.355000 5.525000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  1.785000 11.815000 1.955000 ;
      RECT 11.645000  3.485000 11.815000 3.655000 ;
      RECT 11.645000  5.355000 11.815000 5.525000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.105000  5.355000 12.275000 5.525000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 12.565000  5.355000 12.735000 5.525000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.025000  5.355000 13.195000 5.525000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  1.785000 13.655000 1.955000 ;
      RECT 13.485000  3.485000 13.655000 3.655000 ;
      RECT 13.485000  5.355000 13.655000 5.525000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 13.945000  5.355000 14.115000 5.525000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.405000  5.355000 14.575000 5.525000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 14.865000  5.355000 15.035000 5.525000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.325000  5.355000 15.495000 5.525000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  1.785000 15.955000 1.955000 ;
      RECT 15.785000  3.485000 15.955000 3.655000 ;
      RECT 15.785000  5.355000 15.955000 5.525000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.245000  5.355000 16.415000 5.525000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
      RECT 16.705000  5.355000 16.875000 5.525000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb16to1_1


MACRO sky130_fd_sc_hdll__and4bb_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.995000 0.330000 1.635000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 0.765000 4.525000 1.305000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.270000 0.420000 3.535000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.705000 0.425000 4.005000 1.405000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.255000 1.340000 1.545000 ;
        RECT 1.065000 1.545000 1.420000 1.715000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.720000 0.805000 ;
      RECT 0.175000  1.885000 2.075000 2.055000 ;
      RECT 0.175000  2.055000 0.345000 2.465000 ;
      RECT 0.500000  0.805000 0.720000 1.885000 ;
      RECT 0.515000  0.085000 0.895000 0.465000 ;
      RECT 0.515000  2.255000 0.895000 2.635000 ;
      RECT 1.510000  0.085000 1.890000 0.465000 ;
      RECT 1.515000  0.635000 2.605000 0.805000 ;
      RECT 1.515000  0.805000 1.735000 1.325000 ;
      RECT 1.640000  2.255000 2.310000 2.635000 ;
      RECT 1.905000  0.995000 2.215000 1.325000 ;
      RECT 1.905000  1.325000 2.075000 1.885000 ;
      RECT 2.145000  0.255000 2.315000 0.635000 ;
      RECT 2.385000  0.805000 2.605000 1.915000 ;
      RECT 2.385000  1.915000 3.715000 2.085000 ;
      RECT 2.595000  2.085000 2.765000 2.465000 ;
      RECT 2.795000  1.400000 3.015000 1.575000 ;
      RECT 2.795000  1.575000 4.105000 1.745000 ;
      RECT 2.935000  2.255000 3.325000 2.635000 ;
      RECT 3.545000  2.085000 3.715000 2.465000 ;
      RECT 3.885000  1.745000 4.105000 1.915000 ;
      RECT 3.885000  1.915000 4.915000 2.085000 ;
      RECT 4.105000  2.255000 4.435000 2.635000 ;
      RECT 4.185000  0.085000 4.435000 0.585000 ;
      RECT 4.655000  0.255000 4.915000 0.585000 ;
      RECT 4.655000  2.085000 4.915000 2.465000 ;
      RECT 4.745000  0.585000 4.915000 1.915000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4bb_2


MACRO sky130_fd_sc_hdll__and4bb_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.935000 0.995000 6.345000 1.620000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.765000 0.830000 1.635000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 0.640000 3.840000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.995000 3.195000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.650000 2.280000 0.820000 ;
        RECT 1.010000 0.820000 1.340000 1.545000 ;
        RECT 1.010000 1.545000 2.360000 1.715000 ;
        RECT 1.170000 0.255000 1.340000 0.650000 ;
        RECT 2.110000 0.255000 2.280000 0.650000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.260000 1.915000 ;
      RECT 0.085000  1.915000 4.940000 2.085000 ;
      RECT 0.085000  2.085000 0.345000 2.465000 ;
      RECT 0.515000  2.255000 0.895000 2.635000 ;
      RECT 0.620000  0.085000 0.950000 0.470000 ;
      RECT 1.510000  0.085000 1.890000 0.470000 ;
      RECT 1.510000  1.075000 2.700000 1.245000 ;
      RECT 1.510000  2.255000 1.890000 2.635000 ;
      RECT 2.450000  2.255000 2.830000 2.635000 ;
      RECT 2.470000  0.085000 2.800000 0.445000 ;
      RECT 2.530000  0.615000 3.195000 0.785000 ;
      RECT 2.530000  0.785000 2.700000 1.075000 ;
      RECT 2.530000  1.245000 2.700000 1.545000 ;
      RECT 2.530000  1.545000 4.550000 1.715000 ;
      RECT 2.975000  0.300000 5.060000 0.470000 ;
      RECT 2.975000  0.470000 3.195000 0.615000 ;
      RECT 3.680000  2.255000 4.010000 2.635000 ;
      RECT 4.080000  0.995000 4.300000 1.205000 ;
      RECT 4.080000  1.205000 4.940000 1.375000 ;
      RECT 4.710000  0.470000 5.060000 0.810000 ;
      RECT 4.770000  1.375000 4.940000 1.915000 ;
      RECT 4.810000  2.255000 5.820000 2.635000 ;
      RECT 5.360000  0.655000 6.265000 0.825000 ;
      RECT 5.360000  0.825000 5.530000 1.915000 ;
      RECT 5.360000  1.915000 6.265000 2.085000 ;
      RECT 5.385000  0.085000 5.715000 0.465000 ;
      RECT 6.095000  0.255000 6.265000 0.655000 ;
      RECT 6.095000  2.085000 6.265000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4bb_4


MACRO sky130_fd_sc_hdll__and4bb_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.625000 0.815000 1.955000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 0.765000 0.785000 0.945000 ;
        RECT 0.525000 0.945000 1.165000 1.115000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875000 0.415000 3.175000 1.635000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.345000 0.420000 3.640000 1.635000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.250000 0.255000 4.510000 0.825000 ;
        RECT 4.250000 1.445000 4.510000 2.465000 ;
        RECT 4.285000 0.825000 4.510000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.285000 ;
      RECT 0.085000  1.285000 1.235000 1.455000 ;
      RECT 0.085000  1.455000 0.255000 2.135000 ;
      RECT 0.085000  2.135000 0.345000 2.465000 ;
      RECT 0.575000  0.085000 0.955000 0.465000 ;
      RECT 0.575000  2.255000 0.955000 2.635000 ;
      RECT 1.015000  1.455000 1.235000 1.575000 ;
      RECT 1.015000  1.575000 1.645000 1.745000 ;
      RECT 1.165000  1.915000 1.985000 2.085000 ;
      RECT 1.165000  2.085000 1.375000 2.465000 ;
      RECT 1.185000  0.255000 2.665000 0.425000 ;
      RECT 1.185000  0.425000 1.585000 0.755000 ;
      RECT 1.415000  0.755000 1.585000 1.235000 ;
      RECT 1.415000  1.235000 1.985000 1.405000 ;
      RECT 1.625000  2.255000 1.955000 2.635000 ;
      RECT 1.755000  0.595000 2.325000 0.925000 ;
      RECT 1.815000  1.405000 1.985000 1.915000 ;
      RECT 2.155000  0.925000 2.325000 1.915000 ;
      RECT 2.155000  1.915000 3.980000 2.085000 ;
      RECT 2.185000  2.085000 2.355000 2.465000 ;
      RECT 2.495000  0.425000 2.665000 1.325000 ;
      RECT 2.550000  2.255000 2.930000 2.635000 ;
      RECT 3.210000  2.085000 3.380000 2.465000 ;
      RECT 3.700000  2.255000 4.030000 2.635000 ;
      RECT 3.810000  0.085000 3.980000 0.545000 ;
      RECT 3.810000  0.995000 4.115000 1.325000 ;
      RECT 3.810000  1.325000 3.980000 1.915000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4bb_1


MACRO sky130_fd_sc_hdll__or4b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.630000 0.995000 3.075000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.660000 2.125000 2.860000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.620000 0.995000 2.410000 1.615000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.755000 0.425000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.463700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.620000 0.415000 3.995000 0.760000 ;
        RECT 3.620000 1.495000 3.995000 2.465000 ;
        RECT 3.725000 0.760000 3.995000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.085000 0.425000 0.585000 ;
      RECT 0.085000  1.560000 0.425000 2.635000 ;
      RECT 0.645000  0.305000 0.890000 0.995000 ;
      RECT 0.645000  0.995000 1.300000 1.325000 ;
      RECT 0.645000  1.325000 0.885000 1.920000 ;
      RECT 1.080000  1.495000 1.400000 1.785000 ;
      RECT 1.080000  1.785000 2.860000 1.955000 ;
      RECT 1.085000  0.085000 1.415000 0.585000 ;
      RECT 1.665000  0.305000 1.835000 0.655000 ;
      RECT 1.665000  0.655000 3.415000 0.825000 ;
      RECT 2.010000  0.085000 2.390000 0.485000 ;
      RECT 2.610000  0.305000 2.780000 0.655000 ;
      RECT 2.690000  1.495000 3.415000 1.665000 ;
      RECT 2.690000  1.665000 2.860000 1.785000 ;
      RECT 2.950000  0.085000 3.380000 0.485000 ;
      RECT 3.080000  1.835000 3.360000 2.635000 ;
      RECT 3.245000  0.825000 3.415000 0.995000 ;
      RECT 3.245000  0.995000 3.505000 1.325000 ;
      RECT 3.245000  1.325000 3.415000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4b_1


MACRO sky130_fd_sc_hdll__or4b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.905000 1.075000 2.520000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.185000 2.125000 2.920000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.800000 1.075000 3.900000 1.275000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.435000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 0.260000 1.350000 0.790000 ;
        RECT 1.020000 0.790000 1.235000 1.495000 ;
        RECT 1.020000 1.495000 1.350000 1.825000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.325000 0.350000 0.735000 ;
      RECT 0.085000  0.735000 0.815000 0.905000 ;
      RECT 0.085000  1.605000 0.815000 1.890000 ;
      RECT 0.510000  1.890000 0.815000 1.995000 ;
      RECT 0.510000  1.995000 1.865000 2.165000 ;
      RECT 0.515000  2.335000 0.895000 2.635000 ;
      RECT 0.645000  0.905000 0.815000 1.605000 ;
      RECT 0.680000  0.085000 0.850000 0.565000 ;
      RECT 1.405000  0.960000 1.735000 1.325000 ;
      RECT 1.520000  1.325000 1.735000 1.445000 ;
      RECT 1.520000  1.445000 3.910000 1.615000 ;
      RECT 1.535000  0.085000 1.965000 0.485000 ;
      RECT 1.540000  1.785000 3.330000 1.955000 ;
      RECT 1.540000  1.955000 1.865000 1.995000 ;
      RECT 1.565000  0.700000 3.305000 0.870000 ;
      RECT 1.565000  0.870000 1.735000 0.960000 ;
      RECT 1.630000  2.335000 1.965000 2.635000 ;
      RECT 2.185000  0.270000 2.355000 0.700000 ;
      RECT 2.585000  0.085000 2.915000 0.485000 ;
      RECT 3.135000  0.270000 3.305000 0.700000 ;
      RECT 3.160000  1.955000 3.330000 2.215000 ;
      RECT 3.160000  2.215000 3.695000 2.385000 ;
      RECT 3.525000  0.085000 3.905000 0.585000 ;
      RECT 3.525000  1.615000 3.910000 1.780000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4b_2


MACRO sky130_fd_sc_hdll__or4b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.520000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875000 0.995000 3.175000 1.445000 ;
        RECT 2.875000 1.445000 3.440000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 0.995000 2.705000 2.375000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 0.995000 2.185000 2.375000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.995000 0.445000 1.955000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.695000 1.455000 5.415000 1.625000 ;
        RECT 3.695000 1.625000 3.945000 2.465000 ;
        RECT 3.735000 0.255000 3.985000 0.725000 ;
        RECT 3.735000 0.725000 5.415000 0.905000 ;
        RECT 4.545000 0.255000 4.925000 0.725000 ;
        RECT 4.635000 1.625000 4.885000 2.465000 ;
        RECT 5.175000 0.905000 5.415000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.825000 ;
      RECT 0.085000  2.135000 0.365000 2.635000 ;
      RECT 0.645000  0.435000 0.835000 0.995000 ;
      RECT 0.645000  0.995000 1.265000 1.325000 ;
      RECT 0.645000  1.325000 0.835000 2.455000 ;
      RECT 1.085000  0.085000 1.335000 0.585000 ;
      RECT 1.085000  1.575000 1.725000 1.745000 ;
      RECT 1.085000  1.745000 1.415000 2.450000 ;
      RECT 1.505000  0.655000 3.515000 0.825000 ;
      RECT 1.505000  0.825000 1.725000 1.575000 ;
      RECT 1.715000  0.305000 1.885000 0.655000 ;
      RECT 2.085000  0.085000 2.465000 0.485000 ;
      RECT 2.685000  0.305000 2.855000 0.655000 ;
      RECT 3.125000  0.085000 3.505000 0.485000 ;
      RECT 3.170000  1.795000 3.420000 2.635000 ;
      RECT 3.345000  0.825000 3.515000 1.075000 ;
      RECT 3.345000  1.075000 4.955000 1.245000 ;
      RECT 4.165000  1.795000 4.415000 2.635000 ;
      RECT 4.205000  0.085000 4.375000 0.555000 ;
      RECT 5.105000  1.795000 5.355000 2.635000 ;
      RECT 5.145000  0.085000 5.315000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4b_4


MACRO sky130_fd_sc_hdll__inv_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  1.840000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 0.435000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 0.255000 0.905000 0.885000 ;
        RECT 0.525000 1.485000 0.905000 2.465000 ;
        RECT 0.605000 0.885000 0.905000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.125000  0.085000 0.355000 0.905000 ;
      RECT 0.125000  1.495000 0.355000 2.635000 ;
      RECT 1.125000  0.085000 1.335000 0.905000 ;
      RECT 1.125000  1.495000 1.335000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_2


MACRO sky130_fd_sc_hdll__inv_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  1.380000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.075000 0.650000 1.315000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.770000 0.255000 1.285000 0.885000 ;
        RECT 0.770000 1.485000 1.285000 2.465000 ;
        RECT 0.995000 0.885000 1.285000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.320000  0.085000 0.550000 0.905000 ;
      RECT 0.340000  1.495000 0.550000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_1


MACRO sky130_fd_sc_hdll__inv_12
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  3.330000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.680000 1.075000 5.800000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.020500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 6.320000 0.905000 ;
        RECT 0.085000 0.905000 0.510000 1.495000 ;
        RECT 0.085000 1.495000 6.320000 1.665000 ;
        RECT 0.680000 0.255000 1.060000 0.715000 ;
        RECT 0.680000 1.665000 1.060000 2.465000 ;
        RECT 1.620000 0.255000 2.000000 0.715000 ;
        RECT 1.620000 1.665000 2.000000 2.465000 ;
        RECT 2.560000 0.255000 2.940000 0.715000 ;
        RECT 2.560000 1.665000 2.940000 2.465000 ;
        RECT 3.500000 0.255000 3.880000 0.715000 ;
        RECT 3.500000 1.665000 3.880000 2.465000 ;
        RECT 4.440000 0.255000 4.820000 0.715000 ;
        RECT 4.440000 1.665000 4.820000 2.465000 ;
        RECT 5.380000 0.255000 5.760000 0.715000 ;
        RECT 5.380000 1.665000 5.760000 2.465000 ;
        RECT 5.970000 0.905000 6.320000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.255000  0.085000 0.510000 0.545000 ;
      RECT 0.255000  1.835000 0.510000 2.635000 ;
      RECT 1.280000  0.085000 1.450000 0.545000 ;
      RECT 1.280000  1.835000 1.450000 2.635000 ;
      RECT 2.220000  0.085000 2.390000 0.545000 ;
      RECT 2.220000  1.835000 2.390000 2.635000 ;
      RECT 3.160000  0.085000 3.330000 0.545000 ;
      RECT 3.160000  1.835000 3.330000 2.635000 ;
      RECT 4.100000  0.085000 4.270000 0.545000 ;
      RECT 4.100000  1.835000 4.270000 2.635000 ;
      RECT 5.040000  0.085000 5.210000 0.545000 ;
      RECT 5.040000  1.835000 5.210000 2.635000 ;
      RECT 5.960000  0.085000 6.230000 0.545000 ;
      RECT 5.975000  1.835000 6.230000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_12


MACRO sky130_fd_sc_hdll__inv_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.885000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 0.255000 0.945000 0.725000 ;
        RECT 0.565000 0.725000 2.665000 0.905000 ;
        RECT 0.565000 1.495000 2.665000 1.665000 ;
        RECT 0.565000 1.665000 0.945000 2.465000 ;
        RECT 1.505000 0.255000 1.885000 0.725000 ;
        RECT 1.505000 1.665000 2.665000 1.685000 ;
        RECT 1.505000 1.685000 1.885000 2.465000 ;
        RECT 2.395000 0.905000 2.665000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.130000  0.085000 0.395000 0.545000 ;
      RECT 0.130000  1.495000 0.395000 2.635000 ;
      RECT 1.165000  0.085000 1.335000 0.545000 ;
      RECT 1.165000  1.835000 1.335000 2.635000 ;
      RECT 2.105000  0.085000 2.355000 0.550000 ;
      RECT 2.105000  2.175000 2.315000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_4


MACRO sky130_fd_sc_hdll__inv_6
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.285000 1.075000 2.695000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.494000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.495000 3.265000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.465000 ;
        RECT 0.645000 0.255000 0.815000 0.725000 ;
        RECT 0.645000 0.725000 3.265000 0.905000 ;
        RECT 1.455000 1.665000 1.835000 2.465000 ;
        RECT 1.585000 0.255000 1.755000 0.725000 ;
        RECT 2.395000 1.665000 3.265000 1.685000 ;
        RECT 2.395000 1.685000 2.775000 2.465000 ;
        RECT 2.525000 0.255000 2.695000 0.725000 ;
        RECT 2.865000 0.905000 3.265000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.130000  0.085000 0.395000 0.545000 ;
      RECT 0.175000  1.495000 0.345000 2.635000 ;
      RECT 1.115000  0.085000 1.285000 0.545000 ;
      RECT 1.115000  1.835000 1.285000 2.635000 ;
      RECT 2.055000  0.085000 2.225000 0.545000 ;
      RECT 2.055000  1.835000 2.225000 2.635000 ;
      RECT 2.865000  0.085000 3.165000 0.550000 ;
      RECT 2.995000  2.175000 3.165000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_6


MACRO sky130_fd_sc_hdll__inv_16
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.280000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  4.440000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 6.125000 1.315000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.984000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 0.255000 0.960000 0.715000 ;
        RECT 0.580000 0.715000 7.540000 0.905000 ;
        RECT 0.580000 1.495000 7.540000 1.665000 ;
        RECT 0.580000 1.665000 0.960000 2.465000 ;
        RECT 1.520000 0.255000 1.900000 0.715000 ;
        RECT 1.520000 1.665000 1.900000 2.465000 ;
        RECT 2.460000 0.255000 2.840000 0.715000 ;
        RECT 2.460000 1.665000 2.840000 2.465000 ;
        RECT 3.400000 0.255000 3.780000 0.715000 ;
        RECT 3.400000 1.665000 3.780000 2.465000 ;
        RECT 4.340000 0.255000 4.720000 0.715000 ;
        RECT 4.340000 1.665000 4.720000 2.465000 ;
        RECT 5.280000 0.255000 5.660000 0.715000 ;
        RECT 5.280000 1.665000 5.660000 2.465000 ;
        RECT 6.220000 0.255000 6.600000 0.715000 ;
        RECT 6.220000 1.665000 6.600000 2.465000 ;
        RECT 7.015000 0.905000 7.540000 1.495000 ;
        RECT 7.160000 0.255000 7.540000 0.715000 ;
        RECT 7.160000 1.665000 7.540000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.180000  0.085000 0.410000 0.885000 ;
      RECT 0.200000  1.485000 0.410000 2.635000 ;
      RECT 1.180000  0.085000 1.350000 0.545000 ;
      RECT 1.180000  1.835000 1.350000 2.635000 ;
      RECT 2.120000  0.085000 2.290000 0.545000 ;
      RECT 2.120000  1.835000 2.290000 2.635000 ;
      RECT 3.060000  0.085000 3.230000 0.545000 ;
      RECT 3.060000  1.835000 3.230000 2.635000 ;
      RECT 4.000000  0.085000 4.170000 0.545000 ;
      RECT 4.000000  1.835000 4.170000 2.635000 ;
      RECT 4.940000  0.085000 5.110000 0.545000 ;
      RECT 4.940000  1.835000 5.110000 2.635000 ;
      RECT 5.880000  0.085000 6.050000 0.545000 ;
      RECT 5.880000  1.835000 6.050000 2.635000 ;
      RECT 6.820000  0.085000 6.990000 0.545000 ;
      RECT 6.820000  1.835000 6.990000 2.635000 ;
      RECT 7.760000  0.085000 7.970000 0.885000 ;
      RECT 7.760000  1.835000 7.970000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_16


MACRO sky130_fd_sc_hdll__inv_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.680000 1.075000 3.885000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 4.505000 0.905000 ;
        RECT 0.085000 0.905000 0.430000 1.495000 ;
        RECT 0.085000 1.495000 4.505000 1.665000 ;
        RECT 0.680000 0.255000 1.060000 0.715000 ;
        RECT 0.680000 1.665000 1.060000 2.465000 ;
        RECT 1.620000 0.255000 2.000000 0.715000 ;
        RECT 1.620000 1.665000 2.000000 2.465000 ;
        RECT 2.560000 0.255000 2.940000 0.715000 ;
        RECT 2.560000 1.665000 2.940000 2.465000 ;
        RECT 3.500000 0.255000 3.880000 0.715000 ;
        RECT 3.500000 1.665000 3.880000 2.465000 ;
        RECT 4.185000 0.905000 4.505000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.255000  0.085000 0.510000 0.545000 ;
      RECT 0.255000  1.835000 0.510000 2.635000 ;
      RECT 1.280000  0.085000 1.450000 0.545000 ;
      RECT 1.280000  1.835000 1.450000 2.635000 ;
      RECT 2.220000  0.085000 2.390000 0.545000 ;
      RECT 2.220000  1.835000 2.390000 2.635000 ;
      RECT 3.160000  0.085000 3.330000 0.545000 ;
      RECT 3.160000  1.835000 3.330000 2.635000 ;
      RECT 4.100000  0.085000 4.405000 0.545000 ;
      RECT 4.100000  1.835000 4.400000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_8


MACRO sky130_fd_sc_hdll__a211oi_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.280000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 1.035000 3.305000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.035000 1.535000 1.445000 ;
        RECT 0.100000 1.445000 3.975000 1.625000 ;
        RECT 3.595000 1.035000 3.975000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.225000 1.415000 4.515000 1.460000 ;
        RECT 4.225000 1.460000 7.570000 1.600000 ;
        RECT 4.225000 1.600000 4.515000 1.645000 ;
        RECT 7.280000 1.415000 7.570000 1.460000 ;
        RECT 7.280000 1.600000 7.570000 1.645000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.550000 1.035000 7.050000 1.275000 ;
        RECT 6.830000 1.275000 7.050000 1.695000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.985000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 0.675000 3.680000 0.695000 ;
        RECT 1.925000 0.695000 8.160000 0.825000 ;
        RECT 1.925000 0.825000 7.055000 0.865000 ;
        RECT 4.275000 0.255000 4.645000 0.615000 ;
        RECT 4.275000 0.615000 5.595000 0.625000 ;
        RECT 4.275000 0.625000 8.160000 0.695000 ;
        RECT 5.425000 0.255000 5.595000 0.615000 ;
        RECT 5.720000 1.865000 8.160000 2.085000 ;
        RECT 6.365000 0.255000 6.535000 0.615000 ;
        RECT 6.365000 0.615000 8.160000 0.625000 ;
        RECT 7.680000 1.495000 8.160000 1.865000 ;
        RECT 7.905000 0.825000 8.160000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.095000  0.085000 0.395000 0.585000 ;
      RECT 0.095000  1.795000 4.105000 2.085000 ;
      RECT 0.095000  2.085000 0.345000 2.465000 ;
      RECT 0.515000  2.255000 0.895000 2.635000 ;
      RECT 0.615000  0.530000 0.825000 0.695000 ;
      RECT 0.615000  0.695000 1.755000 0.865000 ;
      RECT 1.000000  0.085000 1.285000 0.525000 ;
      RECT 1.115000  2.085000 4.105000 2.105000 ;
      RECT 1.115000  2.105000 1.285000 2.465000 ;
      RECT 1.455000  0.255000 3.715000 0.505000 ;
      RECT 1.455000  0.505000 1.755000 0.695000 ;
      RECT 1.455000  2.275000 1.835000 2.635000 ;
      RECT 2.055000  2.105000 2.225000 2.465000 ;
      RECT 2.395000  2.275000 2.775000 2.635000 ;
      RECT 2.995000  2.105000 3.165000 2.465000 ;
      RECT 3.335000  2.275000 3.715000 2.635000 ;
      RECT 3.935000  0.085000 4.105000 0.525000 ;
      RECT 3.935000  2.105000 4.105000 2.255000 ;
      RECT 3.935000  2.255000 8.070000 2.465000 ;
      RECT 4.145000  1.035000 5.305000 1.275000 ;
      RECT 4.145000  1.275000 4.960000 1.615000 ;
      RECT 4.275000  1.785000 5.460000 2.085000 ;
      RECT 4.865000  0.085000 5.195000 0.445000 ;
      RECT 5.130000  1.445000 6.610000 1.695000 ;
      RECT 5.130000  1.695000 5.460000 1.785000 ;
      RECT 5.815000  0.085000 6.145000 0.445000 ;
      RECT 6.755000  0.085000 7.085000 0.445000 ;
      RECT 7.300000  0.995000 7.735000 1.325000 ;
      RECT 7.300000  1.325000 7.510000 1.655000 ;
      RECT 7.665000  0.085000 8.070000 0.445000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  1.445000 4.455000 1.615000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.340000  1.445000 7.510000 1.615000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211oi_4


MACRO sky130_fd_sc_hdll__a211oi_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.810000 1.035000 3.570000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.890000 1.035000 4.915000 1.285000 ;
        RECT 4.685000 1.285000 4.915000 1.655000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.035000 1.935000 1.285000 ;
        RECT 1.065000 1.285000 1.285000 1.615000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.995000 0.405000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.008500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 0.255000 0.885000 0.655000 ;
        RECT 0.575000 0.655000 3.395000 0.855000 ;
        RECT 0.575000 0.855000 0.895000 2.115000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.145000  0.085000 0.395000 0.815000 ;
      RECT 0.145000  1.785000 0.405000 2.285000 ;
      RECT 0.145000  2.285000 2.415000 2.455000 ;
      RECT 1.055000  0.085000 1.435000 0.475000 ;
      RECT 1.175000  1.785000 1.365000 2.255000 ;
      RECT 1.175000  2.255000 2.415000 2.285000 ;
      RECT 1.535000  1.455000 4.325000 1.655000 ;
      RECT 1.535000  1.655000 1.915000 2.075000 ;
      RECT 2.015000  0.085000 2.395000 0.475000 ;
      RECT 2.135000  1.835000 2.415000 2.255000 ;
      RECT 2.585000  0.265000 3.795000 0.475000 ;
      RECT 2.635000  1.835000 2.865000 2.635000 ;
      RECT 3.095000  1.655000 3.365000 2.465000 ;
      RECT 3.595000  1.835000 3.825000 2.635000 ;
      RECT 3.625000  0.475000 3.795000 0.635000 ;
      RECT 3.625000  0.635000 4.835000 0.855000 ;
      RECT 3.975000  0.085000 4.355000 0.455000 ;
      RECT 4.055000  1.655000 4.325000 2.465000 ;
      RECT 4.555000  1.835000 4.785000 2.635000 ;
      RECT 4.585000  0.265000 4.835000 0.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211oi_2


MACRO sky130_fd_sc_hdll__a211oi_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.265000 0.905000 0.995000 ;
        RECT 0.605000 0.995000 1.280000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.765000 0.435000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 0.995000 1.795000 2.455000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.980000 0.995000 2.265000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.870200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.155000 0.265000 1.340000 0.625000 ;
        RECT 1.155000 0.625000 2.650000 0.815000 ;
        RECT 1.965000 1.785000 2.650000 2.455000 ;
        RECT 2.255000 0.265000 2.480000 0.625000 ;
        RECT 2.435000 0.815000 2.650000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.085000 0.425000 0.595000 ;
      RECT 0.125000  1.525000 1.330000 1.725000 ;
      RECT 0.125000  1.725000 0.375000 2.455000 ;
      RECT 0.545000  1.905000 0.925000 2.635000 ;
      RECT 1.145000  1.725000 1.330000 2.455000 ;
      RECT 1.550000  0.085000 1.930000 0.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211oi_1


MACRO sky130_fd_sc_hdll__dlrtp_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.820000 BY  2.720000 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.955000 1.765000 1.325000 ;
    END
  END D
  PIN GATE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.435000 1.625000 ;
    END
  END GATE
  PIN Q
    ANTENNADIFFAREA  0.931000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.815000 0.255000 6.195000 0.735000 ;
        RECT 5.815000 0.735000 7.085000 0.905000 ;
        RECT 5.815000 2.255000 6.145000 2.465000 ;
        RECT 5.845000 1.875000 6.145000 2.255000 ;
        RECT 5.895000 1.495000 7.085000 1.665000 ;
        RECT 5.895000 1.665000 6.145000 1.875000 ;
        RECT 6.405000 0.905000 7.085000 1.055000 ;
        RECT 6.405000 1.055000 7.265000 1.325000 ;
        RECT 6.405000 1.325000 7.085000 1.495000 ;
        RECT 6.755000 0.255000 7.085000 0.735000 ;
        RECT 6.755000 1.665000 7.085000 2.465000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.890000 0.995000 5.385000 1.325000 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  1.795000 0.775000 1.965000 ;
      RECT 0.085000  1.965000 0.395000 2.465000 ;
      RECT 0.225000  0.280000 0.395000 0.635000 ;
      RECT 0.225000  0.635000 0.775000 0.805000 ;
      RECT 0.565000  0.085000 0.895000 0.465000 ;
      RECT 0.565000  2.135000 0.895000 2.635000 ;
      RECT 0.605000  0.805000 0.775000 1.070000 ;
      RECT 0.605000  1.070000 0.895000 1.400000 ;
      RECT 0.605000  1.400000 0.775000 1.795000 ;
      RECT 1.065000  0.280000 1.235000 1.685000 ;
      RECT 1.065000  1.685000 1.335000 2.465000 ;
      RECT 1.555000  1.495000 2.115000 1.665000 ;
      RECT 1.555000  1.665000 1.885000 2.465000 ;
      RECT 1.660000  0.345000 1.855000 0.615000 ;
      RECT 1.660000  0.615000 2.115000 0.765000 ;
      RECT 1.660000  0.765000 2.535000 0.785000 ;
      RECT 1.945000  0.785000 2.535000 1.095000 ;
      RECT 1.945000  1.095000 2.115000 1.495000 ;
      RECT 2.025000  0.085000 2.355000 0.445000 ;
      RECT 2.055000  1.835000 2.325000 2.635000 ;
      RECT 2.445000  1.265000 2.955000 1.685000 ;
      RECT 2.780000  0.735000 3.295000 1.095000 ;
      RECT 3.020000  2.165000 3.850000 2.385000 ;
      RECT 3.040000  0.280000 3.660000 0.565000 ;
      RECT 3.125000  1.095000 3.295000 1.575000 ;
      RECT 3.125000  1.575000 3.510000 1.995000 ;
      RECT 3.490000  0.565000 3.660000 0.995000 ;
      RECT 3.490000  0.995000 4.380000 1.165000 ;
      RECT 3.680000  1.165000 4.380000 1.325000 ;
      RECT 3.680000  1.325000 3.850000 2.165000 ;
      RECT 3.870000  0.085000 4.200000 0.610000 ;
      RECT 4.020000  1.535000 5.725000 1.705000 ;
      RECT 4.020000  1.705000 5.175000 1.865000 ;
      RECT 4.020000  2.135000 4.705000 2.635000 ;
      RECT 4.455000  0.255000 4.785000 0.825000 ;
      RECT 4.550000  0.825000 4.720000 1.535000 ;
      RECT 4.875000  1.865000 5.175000 2.435000 ;
      RECT 5.315000  0.085000 5.645000 0.825000 ;
      RECT 5.345000  1.875000 5.675000 2.150000 ;
      RECT 5.345000  2.150000 5.645000 2.635000 ;
      RECT 5.555000  1.075000 6.235000 1.325000 ;
      RECT 5.555000  1.325000 5.725000 1.535000 ;
      RECT 6.315000  1.835000 6.585000 2.635000 ;
      RECT 6.375000  0.085000 6.585000 0.565000 ;
      RECT 7.255000  0.085000 7.465000 0.885000 ;
      RECT 7.255000  1.495000 7.510000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  1.445000 0.775000 1.615000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.115000  1.785000 1.285000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.725000  1.445000 2.895000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.280000  1.785000 3.450000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 0.545000 1.415000 0.835000 1.460000 ;
      RECT 0.545000 1.460000 2.955000 1.600000 ;
      RECT 0.545000 1.600000 0.835000 1.645000 ;
      RECT 1.055000 1.755000 1.345000 1.800000 ;
      RECT 1.055000 1.800000 3.510000 1.940000 ;
      RECT 1.055000 1.940000 1.345000 1.985000 ;
      RECT 2.665000 1.415000 2.955000 1.460000 ;
      RECT 2.665000 1.600000 2.955000 1.645000 ;
      RECT 3.220000 1.755000 3.510000 1.800000 ;
      RECT 3.220000 1.940000 3.510000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtp_4


MACRO sky130_fd_sc_hdll__dlrtp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.955000 1.765000 1.325000 ;
    END
  END D
  PIN GATE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.435000 1.625000 ;
    END
  END GATE
  PIN Q
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.765000 0.255000 6.295000 0.495000 ;
        RECT 5.815000 2.255000 6.295000 2.465000 ;
        RECT 5.820000 0.495000 6.295000 0.885000 ;
        RECT 5.895000 1.495000 6.295000 2.255000 ;
        RECT 6.065000 0.885000 6.295000 1.495000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.890000 0.995000 5.385000 1.325000 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  1.795000 0.775000 1.965000 ;
      RECT 0.085000  1.965000 0.395000 2.465000 ;
      RECT 0.225000  0.280000 0.395000 0.635000 ;
      RECT 0.225000  0.635000 0.775000 0.805000 ;
      RECT 0.565000  0.085000 0.895000 0.465000 ;
      RECT 0.565000  2.135000 0.895000 2.635000 ;
      RECT 0.605000  0.805000 0.775000 1.070000 ;
      RECT 0.605000  1.070000 0.895000 1.400000 ;
      RECT 0.605000  1.400000 0.775000 1.795000 ;
      RECT 1.065000  0.280000 1.235000 1.685000 ;
      RECT 1.065000  1.685000 1.335000 2.465000 ;
      RECT 1.555000  1.495000 2.115000 1.665000 ;
      RECT 1.555000  1.665000 1.885000 2.465000 ;
      RECT 1.660000  0.345000 1.855000 0.615000 ;
      RECT 1.660000  0.615000 2.115000 0.765000 ;
      RECT 1.660000  0.765000 2.535000 0.785000 ;
      RECT 1.945000  0.785000 2.535000 1.095000 ;
      RECT 1.945000  1.095000 2.115000 1.495000 ;
      RECT 2.025000  0.085000 2.355000 0.445000 ;
      RECT 2.055000  1.835000 2.325000 2.635000 ;
      RECT 2.445000  1.265000 2.955000 1.685000 ;
      RECT 2.780000  0.735000 3.295000 1.095000 ;
      RECT 3.020000  2.165000 3.850000 2.385000 ;
      RECT 3.040000  0.280000 3.660000 0.565000 ;
      RECT 3.125000  1.095000 3.295000 1.575000 ;
      RECT 3.125000  1.575000 3.510000 1.995000 ;
      RECT 3.490000  0.565000 3.660000 0.995000 ;
      RECT 3.490000  0.995000 4.380000 1.165000 ;
      RECT 3.680000  1.165000 4.380000 1.325000 ;
      RECT 3.680000  1.325000 3.850000 2.165000 ;
      RECT 3.870000  0.085000 4.200000 0.610000 ;
      RECT 4.020000  1.535000 5.725000 1.705000 ;
      RECT 4.020000  1.705000 5.170000 1.865000 ;
      RECT 4.050000  2.135000 4.635000 2.635000 ;
      RECT 4.455000  0.255000 4.785000 0.825000 ;
      RECT 4.550000  0.825000 4.720000 1.535000 ;
      RECT 4.885000  1.865000 5.170000 2.465000 ;
      RECT 5.320000  0.085000 5.595000 0.625000 ;
      RECT 5.320000  0.625000 5.650000 0.825000 ;
      RECT 5.345000  1.885000 5.675000 2.150000 ;
      RECT 5.345000  2.150000 5.645000 2.635000 ;
      RECT 5.555000  1.055000 5.895000 1.325000 ;
      RECT 5.555000  1.325000 5.725000 1.535000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  1.445000 0.775000 1.615000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.115000  1.785000 1.285000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.725000  1.445000 2.895000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.280000  1.785000 3.450000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.545000 1.415000 0.835000 1.460000 ;
      RECT 0.545000 1.460000 2.955000 1.600000 ;
      RECT 0.545000 1.600000 0.835000 1.645000 ;
      RECT 1.055000 1.755000 1.345000 1.800000 ;
      RECT 1.055000 1.800000 3.510000 1.940000 ;
      RECT 1.055000 1.940000 1.345000 1.985000 ;
      RECT 2.665000 1.415000 2.955000 1.460000 ;
      RECT 2.665000 1.600000 2.955000 1.645000 ;
      RECT 3.220000 1.755000 3.510000 1.800000 ;
      RECT 3.220000 1.940000 3.510000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtp_1


MACRO sky130_fd_sc_hdll__dlrtp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.900000 BY  2.720000 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.955000 1.765000 1.325000 ;
    END
  END D
  PIN GATE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.435000 1.625000 ;
    END
  END GATE
  PIN Q
    ANTENNADIFFAREA  0.465500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.815000 0.255000 6.205000 0.825000 ;
        RECT 5.815000 2.255000 6.205000 2.455000 ;
        RECT 5.895000 1.495000 6.205000 2.255000 ;
        RECT 6.035000 0.825000 6.205000 1.055000 ;
        RECT 6.035000 1.055000 6.435000 1.325000 ;
        RECT 6.035000 1.325000 6.205000 1.495000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.890000 0.995000 5.385000 1.325000 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.085000  1.795000 0.775000 1.965000 ;
      RECT 0.085000  1.965000 0.395000 2.465000 ;
      RECT 0.225000  0.280000 0.395000 0.635000 ;
      RECT 0.225000  0.635000 0.775000 0.805000 ;
      RECT 0.565000  0.085000 0.895000 0.465000 ;
      RECT 0.565000  2.135000 0.895000 2.635000 ;
      RECT 0.605000  0.805000 0.775000 1.070000 ;
      RECT 0.605000  1.070000 0.895000 1.400000 ;
      RECT 0.605000  1.400000 0.775000 1.795000 ;
      RECT 1.065000  0.280000 1.235000 1.685000 ;
      RECT 1.065000  1.685000 1.335000 2.465000 ;
      RECT 1.555000  1.495000 2.115000 1.665000 ;
      RECT 1.555000  1.665000 1.885000 2.465000 ;
      RECT 1.660000  0.345000 1.855000 0.615000 ;
      RECT 1.660000  0.615000 2.115000 0.765000 ;
      RECT 1.660000  0.765000 2.535000 0.785000 ;
      RECT 1.945000  0.785000 2.535000 1.095000 ;
      RECT 1.945000  1.095000 2.115000 1.495000 ;
      RECT 2.025000  0.085000 2.355000 0.445000 ;
      RECT 2.055000  1.835000 2.325000 2.635000 ;
      RECT 2.445000  1.265000 2.955000 1.685000 ;
      RECT 2.780000  0.735000 3.295000 1.095000 ;
      RECT 3.020000  2.165000 3.850000 2.385000 ;
      RECT 3.040000  0.280000 3.660000 0.565000 ;
      RECT 3.125000  1.095000 3.295000 1.575000 ;
      RECT 3.125000  1.575000 3.510000 1.995000 ;
      RECT 3.490000  0.565000 3.660000 0.995000 ;
      RECT 3.490000  0.995000 4.380000 1.165000 ;
      RECT 3.680000  1.165000 4.380000 1.325000 ;
      RECT 3.680000  1.325000 3.850000 2.165000 ;
      RECT 3.870000  0.085000 4.200000 0.610000 ;
      RECT 4.020000  1.535000 5.725000 1.705000 ;
      RECT 4.020000  1.705000 5.170000 1.865000 ;
      RECT 4.050000  2.135000 4.635000 2.635000 ;
      RECT 4.455000  0.255000 4.785000 0.825000 ;
      RECT 4.550000  0.825000 4.720000 1.535000 ;
      RECT 4.885000  1.865000 5.170000 2.465000 ;
      RECT 5.315000  0.085000 5.645000 0.825000 ;
      RECT 5.345000  1.885000 5.675000 2.150000 ;
      RECT 5.345000  2.150000 5.645000 2.635000 ;
      RECT 5.555000  0.995000 5.865000 1.325000 ;
      RECT 5.555000  1.325000 5.725000 1.535000 ;
      RECT 6.375000  0.085000 6.585000 0.885000 ;
      RECT 6.375000  1.495000 6.580000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  1.445000 0.775000 1.615000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.115000  1.785000 1.285000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.725000  1.445000 2.895000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.280000  1.785000 3.450000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
    LAYER met1 ;
      RECT 0.545000 1.415000 0.835000 1.460000 ;
      RECT 0.545000 1.460000 2.955000 1.600000 ;
      RECT 0.545000 1.600000 0.835000 1.645000 ;
      RECT 1.055000 1.755000 1.345000 1.800000 ;
      RECT 1.055000 1.800000 3.510000 1.940000 ;
      RECT 1.055000 1.940000 1.345000 1.985000 ;
      RECT 2.665000 1.415000 2.955000 1.460000 ;
      RECT 2.665000 1.600000 2.955000 1.645000 ;
      RECT 3.220000 1.755000 3.510000 1.800000 ;
      RECT 3.220000 1.940000 3.510000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtp_2


MACRO sky130_fd_sc_hdll__o21ai_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.995000 0.410000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 0.995000 1.075000 1.325000 ;
        RECT 0.580000 1.325000 0.835000 2.375000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.223500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655000 1.295000 2.215000 1.655000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.506200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.505000 1.415000 2.465000 ;
        RECT 1.245000 0.955000 2.110000 1.125000 ;
        RECT 1.245000 1.125000 1.415000 1.505000 ;
        RECT 1.645000 0.275000 2.110000 0.955000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.090000  0.265000 0.380000 0.615000 ;
      RECT 0.090000  0.615000 1.405000 0.785000 ;
      RECT 0.090000  1.495000 0.410000 2.635000 ;
      RECT 0.625000  0.085000 1.005000 0.445000 ;
      RECT 1.175000  0.310000 1.405000 0.615000 ;
      RECT 1.645000  1.835000 2.110000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ai_1


MACRO sky130_fd_sc_hdll__o21ai_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.015000 1.625000 1.320000 ;
        RECT 0.625000 1.320000 1.625000 1.515000 ;
        RECT 0.625000 1.515000 4.095000 1.685000 ;
        RECT 3.795000 0.990000 4.095000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.185000 1.070000 3.625000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.305000 1.015000 5.600000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.661500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.855000 5.700000 2.025000 ;
        RECT 4.335000 1.445000 6.330000 1.700000 ;
        RECT 4.335000 1.700000 5.700000 1.855000 ;
        RECT 4.430000 0.615000 6.330000 0.845000 ;
        RECT 4.530000 2.025000 5.700000 2.085000 ;
        RECT 4.530000 2.085000 4.740000 2.465000 ;
        RECT 5.510000 2.085000 5.700000 2.465000 ;
        RECT 5.920000 0.845000 6.330000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.120000  0.615000 4.260000 0.820000 ;
      RECT 0.120000  1.820000 0.405000 2.635000 ;
      RECT 0.550000  0.085000 0.930000 0.445000 ;
      RECT 0.625000  1.915000 1.820000 2.085000 ;
      RECT 0.625000  2.085000 0.860000 2.465000 ;
      RECT 1.030000  2.255000 1.410000 2.635000 ;
      RECT 1.510000  0.085000 1.890000 0.445000 ;
      RECT 1.630000  2.085000 1.820000 2.275000 ;
      RECT 1.630000  2.275000 3.810000 2.465000 ;
      RECT 2.470000  0.085000 2.850000 0.445000 ;
      RECT 3.430000  0.085000 3.810000 0.445000 ;
      RECT 4.030000  0.255000 6.250000 0.445000 ;
      RECT 4.030000  0.445000 4.260000 0.615000 ;
      RECT 4.030000  2.195000 4.310000 2.635000 ;
      RECT 4.910000  2.255000 5.290000 2.635000 ;
      RECT 5.870000  1.880000 6.250000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ai_4


MACRO sky130_fd_sc_hdll__o21ai_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 1.055000 0.450000 1.445000 ;
        RECT 0.120000 1.445000 2.295000 1.615000 ;
        RECT 1.750000 1.075000 2.295000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.670000 1.075000 1.570000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.280000 0.765000 3.570000 1.400000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.814500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.095000 1.785000 3.110000 1.965000 ;
        RECT 1.095000 1.965000 1.395000 2.125000 ;
        RECT 2.695000 0.595000 3.110000 1.785000 ;
        RECT 2.695000 1.965000 3.110000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.105000  0.255000 0.435000 0.715000 ;
      RECT 0.105000  0.715000 2.465000 0.885000 ;
      RECT 0.105000  1.785000 0.435000 2.635000 ;
      RECT 0.655000  1.785000 0.875000 2.295000 ;
      RECT 0.655000  2.295000 1.865000 2.465000 ;
      RECT 0.665000  0.085000 0.835000 0.545000 ;
      RECT 1.015000  0.255000 1.395000 0.715000 ;
      RECT 1.675000  0.085000 1.845000 0.545000 ;
      RECT 1.675000  2.135000 1.865000 2.295000 ;
      RECT 2.060000  2.175000 2.440000 2.635000 ;
      RECT 2.135000  0.255000 3.530000 0.425000 ;
      RECT 2.135000  0.425000 2.465000 0.715000 ;
      RECT 3.280000  0.425000 3.530000 0.595000 ;
      RECT 3.280000  1.570000 3.530000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ai_2


MACRO sky130_fd_sc_hdll__nand4_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.740000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.115000 1.075000 8.510000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.250000 1.075000 6.115000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.190000 1.075000 4.025000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.835000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.736000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.445000 8.055000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.465000 ;
        RECT 1.455000 1.665000 1.835000 2.465000 ;
        RECT 2.395000 1.665000 2.775000 2.465000 ;
        RECT 3.335000 1.665000 3.715000 2.465000 ;
        RECT 4.795000 1.665000 5.175000 2.465000 ;
        RECT 5.735000 1.665000 6.115000 2.465000 ;
        RECT 6.545000 0.655000 8.055000 0.905000 ;
        RECT 6.545000 0.905000 6.825000 1.445000 ;
        RECT 6.735000 1.665000 7.115000 2.465000 ;
        RECT 7.675000 1.665000 8.055000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.090000  0.255000 0.345000 0.655000 ;
      RECT 0.090000  0.655000 2.225000 0.905000 ;
      RECT 0.090000  1.445000 0.345000 2.635000 ;
      RECT 0.515000  0.085000 0.895000 0.485000 ;
      RECT 1.115000  0.255000 1.285000 0.655000 ;
      RECT 1.115000  1.835000 1.285000 2.635000 ;
      RECT 1.455000  0.085000 1.835000 0.485000 ;
      RECT 2.055000  0.255000 4.185000 0.485000 ;
      RECT 2.055000  0.485000 2.225000 0.655000 ;
      RECT 2.055000  1.835000 2.225000 2.635000 ;
      RECT 2.395000  0.655000 6.115000 0.905000 ;
      RECT 2.995000  1.835000 3.165000 2.635000 ;
      RECT 3.935000  1.835000 4.625000 2.635000 ;
      RECT 4.375000  0.255000 8.530000 0.485000 ;
      RECT 5.395000  1.835000 5.565000 2.635000 ;
      RECT 6.370000  1.835000 6.540000 2.635000 ;
      RECT 7.335000  1.835000 7.505000 2.635000 ;
      RECT 8.275000  0.485000 8.530000 0.905000 ;
      RECT 8.275000  1.445000 8.535000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4_4


MACRO sky130_fd_sc_hdll__nand4_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.175000 0.995000 2.640000 1.665000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 0.300000 1.415000 0.825000 ;
        RECT 1.245000 0.825000 1.415000 0.995000 ;
        RECT 1.245000 0.995000 1.605000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.300000 0.860000 0.995000 ;
        RECT 0.595000 0.995000 1.075000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.995000 0.395000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.867500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.495000 1.945000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.465000 ;
        RECT 1.535000 1.665000 1.865000 2.465000 ;
        RECT 1.670000 0.255000 2.415000 0.825000 ;
        RECT 1.775000 0.825000 1.945000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.090000  0.085000 0.425000 0.825000 ;
      RECT 1.115000  1.835000 1.285000 2.635000 ;
      RECT 2.115000  1.835000 2.395000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4_1


MACRO sky130_fd_sc_hdll__nand4_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.615000 1.075000 4.945000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435000 1.075000 3.380000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.850000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.895000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.368000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.445000 4.325000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.465000 ;
        RECT 1.455000 1.665000 1.835000 2.465000 ;
        RECT 2.555000 1.665000 2.935000 2.465000 ;
        RECT 3.720000 1.055000 4.325000 1.445000 ;
        RECT 3.945000 0.635000 4.325000 1.055000 ;
        RECT 3.945000 1.665000 4.325000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 1.285000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.645000  0.085000 0.815000 0.545000 ;
      RECT 0.985000  0.255000 2.325000 0.465000 ;
      RECT 0.985000  0.465000 1.285000 0.735000 ;
      RECT 1.115000  1.835000 1.285000 2.635000 ;
      RECT 1.455000  0.635000 3.385000 0.905000 ;
      RECT 2.055000  1.835000 2.385000 2.635000 ;
      RECT 2.515000  0.255000 4.875000 0.465000 ;
      RECT 3.295000  1.835000 3.675000 2.635000 ;
      RECT 3.605000  0.465000 3.775000 0.885000 ;
      RECT 4.545000  0.465000 4.875000 0.905000 ;
      RECT 4.545000  1.445000 4.875000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4_2


MACRO sky130_fd_sc_hdll__sedfxbp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  16.56000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795000 0.765000 2.155000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 0.765000 2.765000 1.185000 ;
        RECT 2.325000 1.185000 2.525000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.320000 0.255000 15.700000 2.420000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.935000 1.065000 13.430000 1.300000 ;
        RECT 12.935000 1.300000 13.315000 2.465000 ;
        RECT 13.100000 0.255000 13.430000 1.065000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.445000 1.105000 6.950000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.605000 1.105000 5.885000 1.615000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 16.560000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 16.560000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.560000 0.085000 ;
      RECT  0.000000  2.635000 16.560000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.895000 0.805000 ;
      RECT  0.175000  1.795000  0.895000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.515000  2.135000  0.895000 2.635000 ;
      RECT  0.665000  0.805000  0.895000 1.795000 ;
      RECT  1.115000  0.345000  1.285000 2.465000 ;
      RECT  1.455000  0.255000  1.885000 0.515000 ;
      RECT  1.455000  0.515000  1.625000 1.890000 ;
      RECT  1.455000  1.890000  1.885000 2.465000 ;
      RECT  2.385000  0.085000  2.765000 0.515000 ;
      RECT  2.385000  1.890000  2.765000 2.635000 ;
      RECT  2.695000  1.355000  3.285000 1.720000 ;
      RECT  2.955000  1.720000  3.285000 2.425000 ;
      RECT  2.980000  0.255000  3.205000 0.845000 ;
      RECT  2.980000  0.845000  3.885000 1.175000 ;
      RECT  2.980000  1.175000  3.285000 1.355000 ;
      RECT  3.385000  0.085000  3.765000 0.610000 ;
      RECT  3.515000  1.825000  3.710000 2.635000 ;
      RECT  4.105000  0.685000  4.275000 1.320000 ;
      RECT  4.105000  1.320000  4.525000 1.650000 ;
      RECT  4.425000  1.820000  4.865000 2.020000 ;
      RECT  4.425000  2.020000  4.805000 2.465000 ;
      RECT  4.445000  0.255000  4.765000 0.980000 ;
      RECT  4.445000  0.980000  4.865000 1.150000 ;
      RECT  4.695000  1.150000  4.865000 1.820000 ;
      RECT  4.995000  0.255000  5.195000 0.645000 ;
      RECT  4.995000  0.645000  5.255000 0.825000 ;
      RECT  5.035000  2.210000  5.365000 2.465000 ;
      RECT  5.085000  0.825000  5.255000 1.785000 ;
      RECT  5.085000  1.785000  5.365000 2.210000 ;
      RECT  5.365000  0.255000  6.225000 0.515000 ;
      RECT  5.790000  1.835000  7.370000 2.005000 ;
      RECT  5.790000  2.005000  6.130000 2.465000 ;
      RECT  5.895000  0.515000  6.225000 0.935000 ;
      RECT  6.055000  0.935000  6.225000 1.835000 ;
      RECT  6.350000  2.175000  6.695000 2.635000 ;
      RECT  6.445000  0.085000  6.695000 0.905000 ;
      RECT  7.120000  1.355000  7.370000 1.835000 ;
      RECT  7.300000  0.255000  7.920000 0.565000 ;
      RECT  7.300000  0.565000  7.710000 1.185000 ;
      RECT  7.460000  2.150000  7.790000 2.465000 ;
      RECT  7.540000  1.185000  7.710000 1.865000 ;
      RECT  7.540000  1.865000  7.790000 2.150000 ;
      RECT  7.880000  1.125000  8.115000 1.720000 ;
      RECT  7.900000  0.735000  8.455000 0.955000 ;
      RECT  8.000000  2.175000  9.190000 2.375000 ;
      RECT  8.140000  0.255000  8.865000 0.565000 ;
      RECT  8.285000  0.955000  8.455000 1.655000 ;
      RECT  8.285000  1.655000  8.800000 2.005000 ;
      RECT  8.695000  0.565000  8.865000 1.315000 ;
      RECT  8.695000  1.315000  9.595000 1.485000 ;
      RECT  8.970000  1.485000  9.595000 1.575000 ;
      RECT  8.970000  1.575000  9.190000 2.175000 ;
      RECT  9.055000  0.765000 10.220000 1.045000 ;
      RECT  9.055000  1.045000 10.730000 1.065000 ;
      RECT  9.055000  1.065000  9.305000 1.095000 ;
      RECT  9.180000  0.085000  9.575000 0.560000 ;
      RECT  9.360000  1.835000  9.595000 2.635000 ;
      RECT  9.425000  1.245000  9.595000 1.315000 ;
      RECT  9.765000  0.255000 10.220000 0.765000 ;
      RECT  9.765000  1.065000 10.730000 1.375000 ;
      RECT  9.765000  1.375000 10.145000 2.465000 ;
      RECT 10.355000  2.105000 10.645000 2.635000 ;
      RECT 10.450000  0.085000 10.725000 0.615000 ;
      RECT 11.125000  1.245000 11.365000 1.965000 ;
      RECT 11.260000  2.165000 12.375000 2.355000 ;
      RECT 11.390000  0.705000 11.905000 1.035000 ;
      RECT 11.410000  0.330000 12.375000 0.535000 ;
      RECT 11.535000  1.035000 11.905000 1.995000 ;
      RECT 12.125000  0.535000 12.375000 2.165000 ;
      RECT 12.595000  1.495000 12.765000 2.635000 ;
      RECT 12.630000  0.085000 12.880000 0.900000 ;
      RECT 13.535000  1.465000 13.785000 2.635000 ;
      RECT 13.650000  0.085000 13.900000 0.900000 ;
      RECT 13.955000  1.575000 14.185000 2.010000 ;
      RECT 14.070000  0.890000 14.695000 1.220000 ;
      RECT 14.355000  0.255000 14.695000 0.890000 ;
      RECT 14.355000  1.220000 14.695000 2.465000 ;
      RECT 14.915000  0.085000 15.150000 0.900000 ;
      RECT 14.915000  1.465000 15.150000 2.635000 ;
      RECT 15.920000  0.085000 16.180000 0.900000 ;
      RECT 15.920000  1.465000 16.180000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.685000  1.785000  0.855000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.115000  1.445000  1.285000 1.615000 ;
      RECT  1.455000  0.425000  1.625000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.105000  0.765000  4.275000 0.935000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.535000  0.425000  4.705000 0.595000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.015000  0.425000  5.185000 0.595000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.315000  0.425000  7.485000 0.595000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.910000  1.445000  8.080000 1.615000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.345000  1.785000  8.515000 1.955000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.160000  1.785000 11.330000 1.955000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.630000  1.445000 11.800000 1.615000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.165000  1.785000 12.335000 1.955000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 13.985000  1.785000 14.155000 1.955000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.445000  0.765000 14.615000 0.935000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
    LAYER met1 ;
      RECT  0.625000 1.755000  0.915000 1.800000 ;
      RECT  0.625000 1.800000 11.415000 1.940000 ;
      RECT  0.625000 1.940000  0.915000 1.985000 ;
      RECT  1.005000 1.415000  1.345000 1.460000 ;
      RECT  1.005000 1.460000 11.885000 1.600000 ;
      RECT  1.005000 1.600000  1.345000 1.645000 ;
      RECT  1.395000 0.395000  4.765000 0.580000 ;
      RECT  1.395000 0.580000  1.685000 0.625000 ;
      RECT  4.045000 0.735000  4.335000 0.780000 ;
      RECT  4.045000 0.780000 14.675000 0.920000 ;
      RECT  4.045000 0.920000  4.335000 0.965000 ;
      RECT  4.425000 0.580000  4.765000 0.625000 ;
      RECT  4.905000 0.395000  7.545000 0.580000 ;
      RECT  4.905000 0.580000  5.245000 0.625000 ;
      RECT  7.205000 0.580000  7.545000 0.625000 ;
      RECT  7.825000 1.415000  8.165000 1.460000 ;
      RECT  7.825000 1.600000  8.165000 1.645000 ;
      RECT  8.285000 1.755000  8.625000 1.800000 ;
      RECT  8.285000 1.940000  8.625000 1.985000 ;
      RECT 11.075000 1.755000 11.415000 1.800000 ;
      RECT 11.075000 1.940000 11.415000 1.985000 ;
      RECT 11.545000 1.415000 11.885000 1.460000 ;
      RECT 11.545000 1.600000 11.885000 1.645000 ;
      RECT 12.105000 1.755000 12.395000 1.800000 ;
      RECT 12.105000 1.800000 14.215000 1.940000 ;
      RECT 12.105000 1.940000 12.395000 1.985000 ;
      RECT 13.925000 1.755000 14.215000 1.800000 ;
      RECT 13.925000 1.940000 14.215000 1.985000 ;
      RECT 14.385000 0.735000 14.675000 0.780000 ;
      RECT 14.385000 0.920000 14.675000 0.965000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sedfxbp_2


MACRO sky130_fd_sc_hdll__sedfxbp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  15.18000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795000 0.765000 2.155000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 0.765000 2.765000 1.185000 ;
        RECT 2.325000 1.185000 2.525000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.513200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.655000 0.255000 15.070000 2.420000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.960000 0.255000 13.315000 2.465000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.445000 1.105000 6.950000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.605000 1.105000 5.885000 1.615000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.180000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 15.180000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.180000 0.085000 ;
      RECT  0.000000  2.635000 15.180000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.895000 0.805000 ;
      RECT  0.175000  1.795000  0.895000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.515000  2.135000  0.895000 2.635000 ;
      RECT  0.665000  0.805000  0.895000 1.795000 ;
      RECT  1.115000  0.345000  1.285000 2.465000 ;
      RECT  1.455000  0.255000  1.885000 0.515000 ;
      RECT  1.455000  0.515000  1.625000 1.890000 ;
      RECT  1.455000  1.890000  1.885000 2.465000 ;
      RECT  2.385000  0.085000  2.765000 0.515000 ;
      RECT  2.385000  1.890000  2.765000 2.635000 ;
      RECT  2.695000  1.355000  3.285000 1.720000 ;
      RECT  2.955000  1.720000  3.285000 2.425000 ;
      RECT  2.980000  0.255000  3.205000 0.845000 ;
      RECT  2.980000  0.845000  3.885000 1.175000 ;
      RECT  2.980000  1.175000  3.285000 1.355000 ;
      RECT  3.385000  0.085000  3.765000 0.610000 ;
      RECT  3.515000  1.825000  3.710000 2.635000 ;
      RECT  4.105000  0.685000  4.275000 1.320000 ;
      RECT  4.105000  1.320000  4.525000 1.650000 ;
      RECT  4.425000  1.820000  4.865000 2.020000 ;
      RECT  4.425000  2.020000  4.805000 2.465000 ;
      RECT  4.445000  0.255000  4.765000 0.980000 ;
      RECT  4.445000  0.980000  4.865000 1.150000 ;
      RECT  4.695000  1.150000  4.865000 1.820000 ;
      RECT  4.995000  0.255000  5.195000 0.645000 ;
      RECT  4.995000  0.645000  5.255000 0.825000 ;
      RECT  5.035000  2.210000  5.365000 2.465000 ;
      RECT  5.085000  0.825000  5.255000 1.785000 ;
      RECT  5.085000  1.785000  5.365000 2.210000 ;
      RECT  5.365000  0.255000  6.225000 0.515000 ;
      RECT  5.790000  1.835000  7.370000 2.005000 ;
      RECT  5.790000  2.005000  6.130000 2.465000 ;
      RECT  5.895000  0.515000  6.225000 0.935000 ;
      RECT  6.055000  0.935000  6.225000 1.835000 ;
      RECT  6.350000  2.175000  6.695000 2.635000 ;
      RECT  6.445000  0.085000  6.695000 0.905000 ;
      RECT  7.120000  1.355000  7.370000 1.835000 ;
      RECT  7.300000  0.255000  7.920000 0.565000 ;
      RECT  7.300000  0.565000  7.710000 1.185000 ;
      RECT  7.460000  2.150000  7.790000 2.465000 ;
      RECT  7.540000  1.185000  7.710000 1.865000 ;
      RECT  7.540000  1.865000  7.790000 2.150000 ;
      RECT  7.880000  1.125000  8.115000 1.720000 ;
      RECT  7.900000  0.735000  8.455000 0.955000 ;
      RECT  8.000000  2.175000  9.190000 2.375000 ;
      RECT  8.140000  0.255000  8.865000 0.565000 ;
      RECT  8.285000  0.955000  8.455000 1.655000 ;
      RECT  8.285000  1.655000  8.800000 2.005000 ;
      RECT  8.695000  0.565000  8.865000 1.315000 ;
      RECT  8.695000  1.315000  9.595000 1.485000 ;
      RECT  8.970000  1.485000  9.595000 1.575000 ;
      RECT  8.970000  1.575000  9.190000 2.175000 ;
      RECT  9.055000  0.765000 10.220000 1.045000 ;
      RECT  9.055000  1.045000 10.730000 1.065000 ;
      RECT  9.055000  1.065000  9.305000 1.095000 ;
      RECT  9.180000  0.085000  9.575000 0.560000 ;
      RECT  9.360000  1.835000  9.595000 2.635000 ;
      RECT  9.425000  1.245000  9.595000 1.315000 ;
      RECT  9.765000  0.255000 10.220000 0.765000 ;
      RECT  9.765000  1.065000 10.730000 1.375000 ;
      RECT  9.765000  1.375000 10.145000 2.465000 ;
      RECT 10.355000  2.105000 10.645000 2.635000 ;
      RECT 10.450000  0.085000 10.725000 0.615000 ;
      RECT 11.125000  1.245000 11.365000 1.965000 ;
      RECT 11.260000  2.165000 12.375000 2.355000 ;
      RECT 11.375000  0.705000 11.905000 1.035000 ;
      RECT 11.410000  0.330000 12.375000 0.535000 ;
      RECT 11.535000  1.035000 11.905000 1.995000 ;
      RECT 12.125000  0.535000 12.375000 2.165000 ;
      RECT 12.545000  0.085000 12.790000 0.900000 ;
      RECT 12.595000  1.495000 12.765000 2.635000 ;
      RECT 13.485000  0.890000 13.945000 1.220000 ;
      RECT 13.605000  0.255000 13.945000 0.890000 ;
      RECT 13.605000  1.220000 13.945000 2.465000 ;
      RECT 14.115000  1.070000 14.445000 1.295000 ;
      RECT 14.165000  0.085000 14.400000 0.900000 ;
      RECT 14.165000  1.465000 14.400000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.685000  1.785000  0.855000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.115000  1.445000  1.285000 1.615000 ;
      RECT  1.455000  0.425000  1.625000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.105000  0.765000  4.275000 0.935000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.535000  0.425000  4.705000 0.595000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.015000  0.425000  5.185000 0.595000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.315000  0.425000  7.485000 0.595000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.910000  1.445000  8.080000 1.615000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.345000  1.785000  8.515000 1.955000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.160000  1.785000 11.330000 1.955000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.630000  1.445000 11.800000 1.615000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.165000  1.105000 12.335000 1.275000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.700000  0.765000 13.870000 0.935000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.195000  1.105000 14.365000 1.275000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
    LAYER met1 ;
      RECT  0.625000 1.755000  0.915000 1.800000 ;
      RECT  0.625000 1.800000 11.415000 1.940000 ;
      RECT  0.625000 1.940000  0.915000 1.985000 ;
      RECT  1.005000 1.415000  1.345000 1.460000 ;
      RECT  1.005000 1.460000 11.885000 1.600000 ;
      RECT  1.005000 1.600000  1.345000 1.645000 ;
      RECT  1.395000 0.395000  4.765000 0.580000 ;
      RECT  1.395000 0.580000  1.685000 0.625000 ;
      RECT  4.045000 0.735000  4.335000 0.780000 ;
      RECT  4.045000 0.780000 13.930000 0.920000 ;
      RECT  4.045000 0.920000  4.335000 0.965000 ;
      RECT  4.425000 0.580000  4.765000 0.625000 ;
      RECT  4.905000 0.395000  7.545000 0.580000 ;
      RECT  4.905000 0.580000  5.245000 0.625000 ;
      RECT  7.205000 0.580000  7.545000 0.625000 ;
      RECT  7.825000 1.415000  8.165000 1.460000 ;
      RECT  7.825000 1.600000  8.165000 1.645000 ;
      RECT  8.285000 1.755000  8.625000 1.800000 ;
      RECT  8.285000 1.940000  8.625000 1.985000 ;
      RECT 11.075000 1.755000 11.415000 1.800000 ;
      RECT 11.075000 1.940000 11.415000 1.985000 ;
      RECT 11.545000 1.415000 11.885000 1.460000 ;
      RECT 11.545000 1.600000 11.885000 1.645000 ;
      RECT 12.105000 1.075000 12.395000 1.120000 ;
      RECT 12.105000 1.120000 14.425000 1.260000 ;
      RECT 12.105000 1.260000 12.395000 1.305000 ;
      RECT 13.640000 0.735000 13.930000 0.780000 ;
      RECT 13.640000 0.920000 13.930000 0.965000 ;
      RECT 14.135000 1.075000 14.425000 1.120000 ;
      RECT 14.135000 1.260000 14.425000 1.305000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sedfxbp_1


MACRO sky130_fd_sc_hdll__or3_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.995000 1.490000 1.325000 ;
        RECT 0.605000 1.325000 0.845000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 2.125000 1.375000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.430000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.810200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.340000 0.415000 2.615000 0.760000 ;
        RECT 2.340000 1.495000 2.615000 2.465000 ;
        RECT 2.445000 0.760000 2.615000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.100000  0.305000 0.355000 0.655000 ;
      RECT 0.100000  0.655000 1.975000 0.825000 ;
      RECT 0.105000  1.495000 0.430000 1.785000 ;
      RECT 0.105000  1.785000 1.375000 1.955000 ;
      RECT 0.525000  0.085000 0.905000 0.485000 ;
      RECT 1.125000  0.305000 1.295000 0.655000 ;
      RECT 1.205000  1.495000 1.975000 1.665000 ;
      RECT 1.205000  1.665000 1.375000 1.785000 ;
      RECT 1.465000  0.085000 1.895000 0.485000 ;
      RECT 1.595000  1.835000 1.875000 2.635000 ;
      RECT 1.805000  0.825000 1.975000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3_1


MACRO sky130_fd_sc_hdll__or3_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.995000 1.580000 1.325000 ;
        RECT 0.555000 1.325000 0.880000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 2.125000 1.380000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.385000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.330000 0.415000 2.655000 0.760000 ;
        RECT 2.330000 1.495000 2.655000 2.465000 ;
        RECT 2.470000 0.760000 2.655000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.105000  0.305000 0.360000 0.655000 ;
      RECT 0.105000  0.655000 2.110000 0.825000 ;
      RECT 0.105000  1.495000 0.385000 1.785000 ;
      RECT 0.105000  1.785000 1.370000 1.955000 ;
      RECT 0.530000  0.085000 0.910000 0.485000 ;
      RECT 1.130000  0.305000 1.300000 0.655000 ;
      RECT 1.200000  1.495000 2.110000 1.665000 ;
      RECT 1.200000  1.665000 1.370000 1.785000 ;
      RECT 1.470000  0.085000 2.090000 0.485000 ;
      RECT 1.600000  1.835000 2.070000 2.635000 ;
      RECT 1.890000  0.825000 2.110000 0.995000 ;
      RECT 1.890000  0.995000 2.300000 1.325000 ;
      RECT 1.890000  1.325000 2.110000 1.495000 ;
      RECT 2.825000  0.085000 3.115000 0.915000 ;
      RECT 2.825000  1.430000 3.115000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3_2


MACRO sky130_fd_sc_hdll__or3_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.325000 1.075000 1.850000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 1.075000 1.155000 1.325000 ;
        RECT 0.595000 1.325000 0.830000 2.050000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.455000 0.265000 2.835000 0.735000 ;
        RECT 2.455000 0.735000 4.455000 0.905000 ;
        RECT 2.545000 1.445000 4.455000 1.615000 ;
        RECT 2.545000 1.615000 2.795000 2.465000 ;
        RECT 3.395000 0.265000 3.775000 0.735000 ;
        RECT 3.485000 1.615000 3.735000 2.465000 ;
        RECT 4.115000 0.905000 4.455000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.255000 0.425000 0.725000 ;
      RECT 0.085000  0.725000 2.240000 0.905000 ;
      RECT 0.085000  1.495000 0.425000 2.295000 ;
      RECT 0.085000  2.295000 1.365000 2.465000 ;
      RECT 0.645000  0.085000 0.815000 0.555000 ;
      RECT 0.985000  0.255000 1.365000 0.725000 ;
      RECT 1.100000  1.495000 2.240000 1.665000 ;
      RECT 1.100000  1.665000 1.365000 2.295000 ;
      RECT 1.585000  0.085000 2.285000 0.555000 ;
      RECT 1.585000  1.835000 2.285000 2.635000 ;
      RECT 2.020000  0.905000 2.240000 1.075000 ;
      RECT 2.020000  1.075000 3.945000 1.245000 ;
      RECT 2.020000  1.245000 2.240000 1.495000 ;
      RECT 3.015000  1.795000 3.265000 2.635000 ;
      RECT 3.055000  0.085000 3.225000 0.555000 ;
      RECT 3.955000  1.795000 4.205000 2.635000 ;
      RECT 3.995000  0.085000 4.165000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3_4


MACRO sky130_fd_sc_hdll__or3b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.800000 0.995000 3.110000 1.700000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.330000 0.995000 3.570000 1.700000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.640000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.285000 1.430000 0.735000 ;
        RECT 1.010000 0.735000 2.240000 0.905000 ;
        RECT 1.010000 0.905000 1.270000 1.415000 ;
        RECT 1.010000 1.415000 2.420000 1.700000 ;
        RECT 2.005000 0.255000 2.240000 0.735000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.290000 0.345000 0.735000 ;
      RECT 0.085000  0.735000 0.815000 0.905000 ;
      RECT 0.085000  1.810000 0.815000 1.870000 ;
      RECT 0.085000  1.870000 4.030000 2.040000 ;
      RECT 0.085000  2.040000 0.345000 2.220000 ;
      RECT 0.600000  2.210000 0.960000 2.635000 ;
      RECT 0.645000  0.905000 0.815000 1.810000 ;
      RECT 0.670000  0.085000 0.840000 0.565000 ;
      RECT 1.440000  1.075000 2.615000 1.245000 ;
      RECT 1.520000  2.210000 1.900000 2.635000 ;
      RECT 1.650000  0.085000 1.820000 0.565000 ;
      RECT 2.445000  0.655000 4.455000 0.825000 ;
      RECT 2.445000  0.825000 2.615000 1.075000 ;
      RECT 2.455000  2.210000 2.845000 2.635000 ;
      RECT 2.460000  0.085000 2.840000 0.485000 ;
      RECT 3.400000  0.085000 3.840000 0.485000 ;
      RECT 3.860000  0.995000 4.030000 1.870000 ;
      RECT 3.870000  2.210000 4.455000 2.425000 ;
      RECT 4.250000  0.825000 4.455000 2.210000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3b_4


MACRO sky130_fd_sc_hdll__or3b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 1.075000 2.540000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195000 2.125000 3.545000 2.365000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.640000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.741200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 0.265000 1.385000 0.595000 ;
        RECT 0.985000 0.595000 1.235000 1.495000 ;
        RECT 0.985000 1.495000 1.430000 1.700000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.290000 0.345000 0.735000 ;
      RECT 0.085000  0.735000 0.815000 0.905000 ;
      RECT 0.085000  1.810000 0.815000 1.870000 ;
      RECT 0.085000  1.870000 3.020000 1.955000 ;
      RECT 0.085000  1.955000 1.980000 2.040000 ;
      RECT 0.085000  2.040000 0.345000 2.220000 ;
      RECT 0.600000  2.210000 0.960000 2.635000 ;
      RECT 0.645000  0.085000 0.815000 0.565000 ;
      RECT 0.645000  0.905000 0.815000 1.810000 ;
      RECT 1.485000  0.735000 3.545000 0.825000 ;
      RECT 1.485000  0.825000 2.535000 0.905000 ;
      RECT 1.485000  0.905000 1.655000 1.325000 ;
      RECT 1.685000  2.210000 2.015000 2.635000 ;
      RECT 1.810000  1.785000 3.020000 1.870000 ;
      RECT 1.865000  0.085000 2.035000 0.565000 ;
      RECT 2.365000  0.305000 2.535000 0.655000 ;
      RECT 2.365000  0.655000 3.545000 0.735000 ;
      RECT 2.740000  0.085000 3.070000 0.485000 ;
      RECT 2.850000  0.995000 3.200000 1.325000 ;
      RECT 2.850000  1.325000 3.020000 1.785000 ;
      RECT 3.240000  0.305000 3.545000 0.655000 ;
      RECT 3.240000  1.495000 3.545000 1.925000 ;
      RECT 3.375000  0.825000 3.545000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3b_2


MACRO sky130_fd_sc_hdll__or3b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 2.465000 1.325000 ;
        RECT 1.525000 1.325000 1.770000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 2.125000 2.350000 2.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.325000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.463700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.110000 0.415000 3.535000 0.760000 ;
        RECT 3.110000 1.495000 3.535000 2.465000 ;
        RECT 3.215000 0.760000 3.535000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.905000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.515000  0.485000 0.895000 0.905000 ;
      RECT 0.645000  0.905000 0.895000 0.995000 ;
      RECT 0.645000  0.995000 1.270000 1.325000 ;
      RECT 0.645000  1.325000 0.815000 1.885000 ;
      RECT 1.075000  0.255000 1.335000 0.655000 ;
      RECT 1.075000  0.655000 2.890000 0.825000 ;
      RECT 1.075000  1.495000 1.335000 1.785000 ;
      RECT 1.075000  1.785000 2.350000 1.955000 ;
      RECT 1.505000  0.085000 1.885000 0.485000 ;
      RECT 2.105000  0.305000 2.275000 0.655000 ;
      RECT 2.180000  1.495000 2.890000 1.665000 ;
      RECT 2.180000  1.665000 2.350000 1.785000 ;
      RECT 2.445000  0.085000 2.870000 0.485000 ;
      RECT 2.570000  1.835000 2.850000 2.635000 ;
      RECT 2.720000  0.825000 2.890000 0.995000 ;
      RECT 2.720000  0.995000 2.995000 1.325000 ;
      RECT 2.720000  1.325000 2.890000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3b_1


MACRO sky130_fd_sc_hdll__a2bb2oi_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.475000 1.075000 4.470000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.720000 1.075000 5.435000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.640000 1.445000 ;
        RECT 0.110000 1.445000 2.095000 1.615000 ;
        RECT 1.715000 1.075000 2.095000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 1.075000 1.445000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.738500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 0.645000 1.365000 0.725000 ;
        RECT 0.985000 0.725000 2.775000 0.905000 ;
        RECT 2.395000 0.255000 2.775000 0.725000 ;
        RECT 2.445000 0.905000 2.775000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.135000  1.785000 2.265000 1.955000 ;
      RECT 0.135000  1.955000 0.385000 2.465000 ;
      RECT 0.175000  0.085000 0.345000 0.895000 ;
      RECT 0.515000  0.255000 1.835000 0.475000 ;
      RECT 0.515000  0.475000 0.815000 0.895000 ;
      RECT 0.605000  2.135000 0.855000 2.635000 ;
      RECT 1.075000  1.955000 1.325000 2.465000 ;
      RECT 1.545000  2.135000 1.795000 2.635000 ;
      RECT 2.015000  1.955000 2.265000 2.295000 ;
      RECT 2.015000  2.295000 3.205000 2.465000 ;
      RECT 2.055000  0.085000 2.225000 0.555000 ;
      RECT 2.955000  1.795000 3.205000 2.295000 ;
      RECT 2.995000  0.085000 3.685000 0.555000 ;
      RECT 2.995000  0.995000 3.285000 1.325000 ;
      RECT 3.115000  0.725000 5.175000 0.905000 ;
      RECT 3.115000  0.905000 3.285000 0.995000 ;
      RECT 3.115000  1.325000 3.285000 1.445000 ;
      RECT 3.115000  1.445000 5.135000 1.615000 ;
      RECT 3.475000  1.785000 4.665000 1.965000 ;
      RECT 3.475000  1.965000 3.725000 2.465000 ;
      RECT 3.855000  0.255000 4.235000 0.725000 ;
      RECT 3.945000  2.135000 4.195000 2.635000 ;
      RECT 4.415000  1.965000 4.665000 2.295000 ;
      RECT 4.415000  2.295000 5.605000 2.465000 ;
      RECT 4.455000  0.085000 4.625000 0.555000 ;
      RECT 4.795000  0.255000 5.175000 0.725000 ;
      RECT 4.885000  1.615000 5.135000 2.125000 ;
      RECT 5.355000  1.455000 5.605000 2.295000 ;
      RECT 5.395000  0.085000 5.565000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2oi_2


MACRO sky130_fd_sc_hdll__a2bb2oi_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.995000 0.520000 1.615000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.775000 1.010000 1.340000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.885000 0.995000 3.225000 1.615000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385000 0.995000 2.615000 1.615000 ;
        RECT 2.445000 0.425000 2.615000 0.995000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.530000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 1.785000 2.155000 1.955000 ;
        RECT 1.520000 1.955000 1.885000 2.465000 ;
        RECT 1.985000 0.255000 2.275000 0.825000 ;
        RECT 1.985000 0.825000 2.155000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
        RECT 0.095000  0.085000 0.425000 0.825000 ;
        RECT 1.045000  0.085000 1.715000 0.490000 ;
        RECT 3.005000  0.085000 3.385000 0.825000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
        RECT 0.095000 1.805000 0.425000 2.635000 ;
        RECT 2.665000 2.135000 2.915000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.645000 0.255000 0.815000 0.660000 ;
      RECT 0.645000 0.660000 1.815000 0.830000 ;
      RECT 0.925000 1.445000 1.815000 1.615000 ;
      RECT 0.925000 1.615000 1.305000 2.465000 ;
      RECT 1.645000 0.830000 1.815000 1.445000 ;
      RECT 2.055000 2.235000 2.495000 2.465000 ;
      RECT 2.325000 1.785000 3.390000 1.955000 ;
      RECT 2.325000 1.955000 2.495000 2.235000 ;
      RECT 3.135000 1.955000 3.390000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2oi_1


MACRO sky130_fd_sc_hdll__a2bb2oi_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.58000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.545000 1.075000 8.070000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.440000 1.075000 9.965000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 1.705000 1.285000 ;
        RECT 1.535000 1.285000 1.705000 1.445000 ;
        RECT 1.535000 1.445000 3.975000 1.615000 ;
        RECT 3.595000 1.075000 3.975000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.875000 1.075000 3.425000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.477000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 0.645000 3.295000 0.725000 ;
        RECT 1.925000 0.725000 5.595000 0.905000 ;
        RECT 4.145000 0.905000 4.365000 1.415000 ;
        RECT 4.145000 1.415000 5.515000 1.615000 ;
        RECT 4.275000 0.275000 4.655000 0.725000 ;
        RECT 4.365000 1.615000 4.615000 2.125000 ;
        RECT 5.215000 0.275000 5.595000 0.725000 ;
        RECT 5.245000 1.615000 5.515000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.085000  1.455000  1.315000 1.625000 ;
      RECT  0.085000  1.625000  0.425000 2.465000 ;
      RECT  0.175000  0.085000  0.345000 0.895000 ;
      RECT  0.515000  0.255000  0.895000 0.725000 ;
      RECT  0.515000  0.725000  1.755000 0.905000 ;
      RECT  0.645000  1.795000  0.855000 2.635000 ;
      RECT  1.075000  1.625000  1.315000 1.795000 ;
      RECT  1.075000  1.795000  4.145000 1.965000 ;
      RECT  1.075000  1.965000  1.315000 2.465000 ;
      RECT  1.115000  0.085000  1.285000 0.555000 ;
      RECT  1.455000  0.255000  3.715000 0.475000 ;
      RECT  1.455000  0.475000  1.755000 0.725000 ;
      RECT  1.545000  2.135000  1.795000 2.635000 ;
      RECT  2.015000  1.965000  2.265000 2.465000 ;
      RECT  2.485000  2.135000  2.735000 2.635000 ;
      RECT  2.955000  1.965000  3.205000 2.465000 ;
      RECT  3.425000  2.135000  3.675000 2.635000 ;
      RECT  3.895000  1.965000  4.145000 2.295000 ;
      RECT  3.895000  2.295000  6.065000 2.465000 ;
      RECT  3.935000  0.085000  4.105000 0.555000 ;
      RECT  4.535000  1.075000  6.325000 1.245000 ;
      RECT  4.835000  1.795000  5.075000 2.295000 ;
      RECT  4.875000  0.085000  5.045000 0.555000 ;
      RECT  5.685000  1.455000  6.065000 2.295000 ;
      RECT  5.815000  0.085000  6.505000 0.555000 ;
      RECT  6.155000  0.735000 10.460000 0.905000 ;
      RECT  6.155000  0.905000  6.325000 1.075000 ;
      RECT  6.255000  1.455000  8.425000 1.625000 ;
      RECT  6.255000  1.625000  6.585000 2.465000 ;
      RECT  6.675000  0.255000  7.055000 0.725000 ;
      RECT  6.675000  0.725000  9.875000 0.735000 ;
      RECT  6.805000  1.795000  7.015000 2.635000 ;
      RECT  7.240000  1.625000  7.480000 2.465000 ;
      RECT  7.275000  0.085000  7.445000 0.555000 ;
      RECT  7.615000  0.255000  7.995000 0.725000 ;
      RECT  7.705000  1.795000  7.955000 2.635000 ;
      RECT  8.175000  1.625000  8.425000 2.295000 ;
      RECT  8.175000  2.295000 10.310000 2.465000 ;
      RECT  8.215000  0.085000  8.385000 0.555000 ;
      RECT  8.555000  0.255000  8.935000 0.725000 ;
      RECT  8.645000  1.455000 10.460000 1.625000 ;
      RECT  8.645000  1.625000  8.895000 2.125000 ;
      RECT  9.115000  1.795000  9.365000 2.295000 ;
      RECT  9.155000  0.085000  9.325000 0.555000 ;
      RECT  9.495000  0.255000  9.875000 0.725000 ;
      RECT  9.585000  1.625000  9.835000 2.125000 ;
      RECT 10.060000  1.795000 10.310000 2.295000 ;
      RECT 10.095000  0.085000 10.265000 0.555000 ;
      RECT 10.135000  0.905000 10.460000 1.455000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2oi_4


MACRO sky130_fd_sc_hdll__nor3b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 0.995000 1.815000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 0.995000 1.305000 1.615000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.995000 2.335000 1.615000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  0.759000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.605000 0.655000 ;
        RECT 0.085000 0.655000 1.545000 0.825000 ;
        RECT 0.085000 0.825000 0.255000 1.445000 ;
        RECT 0.085000 1.445000 0.545000 2.455000 ;
        RECT 1.375000 0.310000 1.545000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.425000  1.075000 0.885000 1.245000 ;
      RECT 0.715000  1.245000 0.885000 1.785000 ;
      RECT 0.715000  1.785000 2.675000 1.955000 ;
      RECT 0.775000  0.085000 1.155000 0.485000 ;
      RECT 1.715000  0.085000 2.095000 0.825000 ;
      RECT 1.715000  2.125000 2.095000 2.635000 ;
      RECT 2.380000  0.405000 2.550000 0.655000 ;
      RECT 2.380000  0.655000 2.675000 0.825000 ;
      RECT 2.505000  0.825000 2.675000 1.785000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3b_1


MACRO sky130_fd_sc_hdll__nor3b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.015000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.235000 1.075000 2.200000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.330000 1.075000 4.915000 1.285000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  0.979000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 3.355000 0.905000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 2.870000 0.905000 3.355000 2.045000 ;
        RECT 2.935000 0.255000 3.355000 0.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 2.325000 1.625000 ;
      RECT 0.090000  1.625000 0.405000 2.465000 ;
      RECT 0.625000  1.795000 0.875000 2.635000 ;
      RECT 1.095000  1.625000 1.345000 2.465000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 1.565000  1.795000 1.815000 2.275000 ;
      RECT 1.565000  2.275000 3.780000 2.465000 ;
      RECT 1.995000  1.625000 2.325000 2.035000 ;
      RECT 2.075000  0.085000 2.765000 0.555000 ;
      RECT 3.535000  1.075000 4.160000 1.285000 ;
      RECT 3.535000  1.455000 3.780000 2.275000 ;
      RECT 3.575000  0.085000 3.780000 0.895000 ;
      RECT 3.990000  0.380000 4.345000 0.905000 ;
      RECT 3.990000  0.905000 4.160000 1.075000 ;
      RECT 3.990000  1.285000 4.160000 1.455000 ;
      RECT 3.990000  1.455000 4.345000 1.870000 ;
      RECT 4.565000  0.085000 4.855000 0.825000 ;
      RECT 4.565000  1.540000 4.815000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3b_2


MACRO sky130_fd_sc_hdll__nor3b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.360000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.210000 1.075000 2.770000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.285000 1.075000 4.700000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.445000 1.285000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  1.925500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 0.255000 1.385000 0.725000 ;
        RECT 1.005000 0.725000 7.245000 0.905000 ;
        RECT 1.945000 0.255000 2.325000 0.725000 ;
        RECT 3.405000 0.255000 3.785000 0.725000 ;
        RECT 4.345000 0.255000 4.725000 0.725000 ;
        RECT 5.285000 0.255000 5.665000 0.725000 ;
        RECT 5.375000 1.455000 7.245000 1.625000 ;
        RECT 5.375000 1.625000 5.625000 2.125000 ;
        RECT 6.225000 0.255000 6.605000 0.725000 ;
        RECT 6.315000 1.625000 6.565000 2.125000 ;
        RECT 6.905000 0.905000 7.245000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.110000  0.255000 0.445000 0.735000 ;
      RECT 0.110000  0.735000 0.835000 0.905000 ;
      RECT 0.110000  1.455000 5.155000 1.625000 ;
      RECT 0.110000  1.625000 0.405000 2.465000 ;
      RECT 0.625000  1.795000 0.875000 2.635000 ;
      RECT 0.665000  0.085000 0.835000 0.555000 ;
      RECT 0.665000  0.905000 0.835000 1.455000 ;
      RECT 1.095000  1.795000 4.685000 1.965000 ;
      RECT 1.095000  1.965000 1.345000 2.465000 ;
      RECT 1.565000  2.135000 1.815000 2.635000 ;
      RECT 1.605000  0.085000 1.775000 0.555000 ;
      RECT 2.035000  1.965000 2.285000 2.465000 ;
      RECT 2.505000  2.135000 2.755000 2.635000 ;
      RECT 2.545000  0.085000 3.235000 0.555000 ;
      RECT 3.025000  2.135000 3.275000 2.295000 ;
      RECT 3.025000  2.295000 7.035000 2.465000 ;
      RECT 3.495000  1.965000 3.745000 2.125000 ;
      RECT 3.965000  2.135000 4.215000 2.295000 ;
      RECT 4.005000  0.085000 4.175000 0.555000 ;
      RECT 4.435000  1.965000 4.685000 2.125000 ;
      RECT 4.905000  1.795000 5.155000 2.295000 ;
      RECT 4.945000  0.085000 5.115000 0.555000 ;
      RECT 4.985000  1.075000 6.720000 1.285000 ;
      RECT 4.985000  1.285000 5.155000 1.455000 ;
      RECT 5.845000  1.795000 6.095000 2.295000 ;
      RECT 5.885000  0.085000 6.055000 0.555000 ;
      RECT 6.785000  1.795000 7.035000 2.295000 ;
      RECT 6.825000  0.085000 6.995000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3b_4


MACRO sky130_fd_sc_hdll__o2bb2a_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.820000 1.075000 1.320000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 0.380000 1.300000 0.735000 ;
        RECT 1.015000 0.735000 1.715000 0.905000 ;
        RECT 1.490000 0.905000 1.715000 1.100000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.705000 1.075000 4.055000 1.645000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.720000 1.075000 3.535000 1.325000 ;
        RECT 3.335000 1.325000 3.535000 2.425000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.471500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 0.825000 ;
        RECT 0.085000 0.825000 0.260000 1.795000 ;
        RECT 0.085000 1.795000 0.345000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.430000  0.995000 0.650000 1.445000 ;
      RECT 0.430000  1.445000 0.875000 1.615000 ;
      RECT 0.515000  2.235000 0.895000 2.635000 ;
      RECT 0.670000  0.085000 0.840000 0.750000 ;
      RECT 0.705000  1.615000 0.875000 1.885000 ;
      RECT 0.705000  1.885000 2.935000 2.055000 ;
      RECT 1.045000  1.495000 2.160000 1.715000 ;
      RECT 1.560000  0.395000 2.055000 0.565000 ;
      RECT 1.865000  2.235000 2.265000 2.635000 ;
      RECT 1.885000  0.565000 2.055000 1.355000 ;
      RECT 1.885000  1.355000 2.160000 1.495000 ;
      RECT 2.225000  0.320000 2.475000 0.690000 ;
      RECT 2.305000  0.690000 2.475000 1.075000 ;
      RECT 2.305000  1.075000 2.500000 1.245000 ;
      RECT 2.330000  1.245000 2.500000 1.495000 ;
      RECT 2.330000  1.495000 2.935000 1.885000 ;
      RECT 2.555000  2.055000 2.935000 2.290000 ;
      RECT 2.695000  0.320000 2.945000 0.725000 ;
      RECT 2.695000  0.725000 4.055000 0.905000 ;
      RECT 3.135000  0.085000 3.485000 0.555000 ;
      RECT 3.665000  0.320000 4.055000 0.725000 ;
      RECT 3.705000  1.815000 4.055000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2a_1


MACRO sky130_fd_sc_hdll__o2bb2a_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.075000 1.835000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 0.380000 1.885000 0.735000 ;
        RECT 1.520000 0.735000 2.225000 0.905000 ;
        RECT 2.005000 0.905000 2.225000 1.100000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.000000 1.075000 4.465000 1.645000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.220000 1.075000 3.825000 1.325000 ;
        RECT 3.655000 1.325000 3.825000 1.915000 ;
        RECT 3.655000 1.915000 3.995000 2.425000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.920000 0.825000 ;
        RECT 0.535000 0.825000 0.755000 1.795000 ;
        RECT 0.535000 1.795000 0.840000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.110000  0.085000 0.365000 0.910000 ;
      RECT 0.110000  1.410000 0.365000 2.635000 ;
      RECT 0.925000  0.995000 1.145000 1.445000 ;
      RECT 0.925000  1.445000 1.370000 1.615000 ;
      RECT 1.010000  2.235000 1.390000 2.635000 ;
      RECT 1.135000  0.085000 1.305000 0.750000 ;
      RECT 1.200000  1.615000 1.370000 1.885000 ;
      RECT 1.200000  1.885000 3.435000 2.055000 ;
      RECT 1.540000  1.495000 2.660000 1.715000 ;
      RECT 2.055000  0.395000 2.565000 0.565000 ;
      RECT 2.360000  2.235000 2.765000 2.635000 ;
      RECT 2.395000  0.565000 2.565000 1.355000 ;
      RECT 2.395000  1.355000 2.660000 1.495000 ;
      RECT 2.735000  0.320000 2.980000 0.690000 ;
      RECT 2.810000  0.690000 2.980000 1.075000 ;
      RECT 2.810000  1.075000 3.000000 1.245000 ;
      RECT 2.830000  1.245000 3.000000 1.495000 ;
      RECT 2.830000  1.495000 3.435000 1.885000 ;
      RECT 3.035000  2.055000 3.435000 2.425000 ;
      RECT 3.205000  0.320000 3.435000 0.725000 ;
      RECT 3.205000  0.725000 4.405000 0.905000 ;
      RECT 3.675000  0.085000 3.845000 0.555000 ;
      RECT 4.015000  0.320000 4.405000 0.725000 ;
      RECT 4.165000  1.815000 4.480000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2a_2


MACRO sky130_fd_sc_hdll__o2bb2a_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.820000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.615000 1.075000 3.995000 1.445000 ;
        RECT 3.615000 1.445000 5.465000 1.615000 ;
        RECT 5.055000 1.075000 5.465000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 1.075000 4.885000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.625000 1.445000 ;
        RECT 0.085000 1.445000 2.095000 1.615000 ;
        RECT 1.715000 1.075000 2.095000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 1.075000 1.445000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.735000 0.275000 6.115000 0.725000 ;
        RECT 5.735000 0.725000 7.710000 0.905000 ;
        RECT 5.825000 1.785000 7.015000 1.955000 ;
        RECT 5.825000 1.955000 6.075000 2.465000 ;
        RECT 6.675000 0.275000 7.055000 0.725000 ;
        RECT 6.765000 1.415000 7.710000 1.655000 ;
        RECT 6.765000 1.655000 7.015000 1.785000 ;
        RECT 6.765000 1.955000 7.015000 2.465000 ;
        RECT 7.405000 0.905000 7.710000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.095000  0.255000 0.425000 0.725000 ;
      RECT 0.095000  0.725000 1.365000 0.735000 ;
      RECT 0.095000  0.735000 2.225000 0.905000 ;
      RECT 0.140000  1.795000 0.345000 2.635000 ;
      RECT 0.605000  1.785000 0.855000 2.295000 ;
      RECT 0.605000  2.295000 1.795000 2.465000 ;
      RECT 0.645000  0.085000 0.815000 0.555000 ;
      RECT 0.985000  0.255000 1.365000 0.725000 ;
      RECT 1.075000  1.785000 2.865000 1.955000 ;
      RECT 1.075000  1.955000 1.325000 2.125000 ;
      RECT 1.545000  2.125000 1.795000 2.295000 ;
      RECT 1.585000  0.085000 1.755000 0.555000 ;
      RECT 1.925000  0.255000 3.245000 0.475000 ;
      RECT 1.925000  0.475000 2.225000 0.735000 ;
      RECT 2.015000  2.125000 2.265000 2.635000 ;
      RECT 2.265000  1.075000 2.695000 1.415000 ;
      RECT 2.265000  1.415000 2.865000 1.785000 ;
      RECT 2.395000  0.645000 2.775000 0.815000 ;
      RECT 2.395000  0.815000 2.695000 1.075000 ;
      RECT 2.485000  1.955000 2.865000 1.965000 ;
      RECT 2.485000  1.965000 2.775000 2.465000 ;
      RECT 2.865000  1.075000 3.445000 1.245000 ;
      RECT 2.995000  2.135000 3.725000 2.635000 ;
      RECT 3.255000  0.725000 4.705000 0.905000 ;
      RECT 3.255000  0.905000 3.445000 1.075000 ;
      RECT 3.255000  1.245000 3.445000 1.785000 ;
      RECT 3.255000  1.785000 5.135000 1.965000 ;
      RECT 3.515000  0.085000 3.685000 0.555000 ;
      RECT 3.855000  0.305000 5.175000 0.475000 ;
      RECT 3.945000  1.965000 4.195000 2.125000 ;
      RECT 4.325000  0.645000 4.705000 0.725000 ;
      RECT 4.415000  2.135000 4.665000 2.635000 ;
      RECT 4.885000  1.965000 5.135000 2.465000 ;
      RECT 4.925000  0.475000 5.175000 0.895000 ;
      RECT 5.355000  1.795000 5.605000 2.635000 ;
      RECT 5.395000  0.085000 5.565000 0.895000 ;
      RECT 5.665000  1.075000 7.085000 1.245000 ;
      RECT 5.665000  1.245000 6.005000 1.615000 ;
      RECT 6.295000  2.165000 6.545000 2.635000 ;
      RECT 6.335000  0.085000 6.505000 0.555000 ;
      RECT 7.235000  1.825000 7.485000 2.635000 ;
      RECT 7.275000  0.085000 7.445000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.695000  1.435000 2.865000 1.605000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.725000  1.445000 5.895000 1.615000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 2.635000 1.385000 2.975000 1.460000 ;
      RECT 2.635000 1.460000 5.960000 1.600000 ;
      RECT 2.635000 1.600000 2.975000 1.635000 ;
      RECT 5.665000 1.395000 5.960000 1.460000 ;
      RECT 5.665000 1.600000 5.960000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2a_4


MACRO sky130_fd_sc_hdll__o21bai_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 1.075000 4.455000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.175000 1.075000 3.390000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.480000 1.325000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.788000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.185000 1.445000 2.900000 1.615000 ;
        RECT 1.185000 1.615000 1.355000 2.465000 ;
        RECT 1.510000 0.645000 2.005000 1.445000 ;
        RECT 2.655000 1.615000 2.900000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.180000  0.085000 0.350000 0.825000 ;
      RECT 0.180000  1.495000 0.915000 1.665000 ;
      RECT 0.180000  1.665000 0.350000 1.915000 ;
      RECT 0.635000  1.875000 0.965000 2.635000 ;
      RECT 0.650000  0.445000 0.820000 1.075000 ;
      RECT 0.650000  1.075000 1.340000 1.245000 ;
      RECT 0.650000  1.245000 0.915000 1.495000 ;
      RECT 1.060000  0.255000 2.475000 0.475000 ;
      RECT 1.060000  0.475000 1.340000 0.905000 ;
      RECT 1.620000  1.795000 1.870000 2.635000 ;
      RECT 2.105000  1.795000 2.435000 2.295000 ;
      RECT 2.105000  2.295000 3.335000 2.465000 ;
      RECT 2.225000  0.475000 2.475000 0.725000 ;
      RECT 2.225000  0.725000 4.380000 0.905000 ;
      RECT 2.695000  0.085000 2.865000 0.555000 ;
      RECT 3.035000  0.255000 3.415000 0.725000 ;
      RECT 3.165000  1.455000 4.380000 1.665000 ;
      RECT 3.165000  1.665000 3.335000 2.295000 ;
      RECT 3.505000  1.835000 3.885000 2.635000 ;
      RECT 3.635000  0.085000 3.805000 0.555000 ;
      RECT 3.975000  0.265000 4.380000 0.725000 ;
      RECT 4.105000  1.665000 4.380000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21bai_2


MACRO sky130_fd_sc_hdll__o21bai_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.360000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.145000 1.075000 7.250000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.075000 4.975000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.510000 1.285000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.576000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.455000 4.765000 1.625000 ;
        RECT 1.035000 1.625000 1.375000 2.465000 ;
        RECT 1.520000 0.645000 2.925000 0.815000 ;
        RECT 2.065000 1.625000 2.315000 2.465000 ;
        RECT 2.695000 0.815000 2.925000 1.075000 ;
        RECT 2.695000 1.075000 3.195000 1.445000 ;
        RECT 2.695000 1.445000 4.765000 1.455000 ;
        RECT 3.575000 1.625000 3.825000 2.125000 ;
        RECT 4.515000 1.625000 4.765000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.145000  1.455000 0.850000 1.625000 ;
      RECT 0.145000  1.625000 0.475000 2.435000 ;
      RECT 0.225000  0.085000 0.395000 0.895000 ;
      RECT 0.565000  0.290000 0.945000 0.895000 ;
      RECT 0.680000  0.895000 0.945000 1.075000 ;
      RECT 0.680000  1.075000 2.525000 1.285000 ;
      RECT 0.680000  1.285000 0.850000 1.455000 ;
      RECT 0.695000  1.795000 0.865000 2.635000 ;
      RECT 1.180000  0.305000 3.395000 0.475000 ;
      RECT 1.595000  1.795000 1.845000 2.635000 ;
      RECT 2.535000  1.795000 2.785000 2.635000 ;
      RECT 3.025000  1.795000 3.355000 2.295000 ;
      RECT 3.025000  2.295000 5.235000 2.465000 ;
      RECT 3.145000  0.475000 3.395000 0.725000 ;
      RECT 3.145000  0.725000 7.155000 0.905000 ;
      RECT 3.615000  0.085000 3.785000 0.555000 ;
      RECT 3.955000  0.255000 4.335000 0.725000 ;
      RECT 4.045000  1.795000 4.295000 2.295000 ;
      RECT 4.555000  0.085000 4.725000 0.555000 ;
      RECT 4.895000  0.255000 5.275000 0.725000 ;
      RECT 4.985000  1.455000 7.115000 1.625000 ;
      RECT 4.985000  1.625000 5.235000 2.295000 ;
      RECT 5.455000  1.795000 5.705000 2.635000 ;
      RECT 5.495000  0.085000 5.665000 0.555000 ;
      RECT 5.835000  0.255000 6.215000 0.725000 ;
      RECT 5.925000  1.625000 6.175000 2.465000 ;
      RECT 6.395000  1.795000 6.645000 2.635000 ;
      RECT 6.435000  0.085000 6.605000 0.555000 ;
      RECT 6.775000  0.255000 7.155000 0.725000 ;
      RECT 6.865000  1.625000 7.115000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21bai_4


MACRO sky130_fd_sc_hdll__o21bai_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365000 1.075000 2.925000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.675000 1.075000 2.195000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.535000 1.345000 ;
        RECT 0.085000 1.345000 0.355000 2.445000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.521500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.235000 0.255000 1.455000 1.445000 ;
        RECT 1.235000 1.445000 2.155000 1.625000 ;
        RECT 1.635000 1.625000 2.155000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.360000 0.825000 ;
      RECT 0.525000  1.535000 1.065000 1.705000 ;
      RECT 0.525000  1.705000 0.850000 2.210000 ;
      RECT 0.675000  0.495000 0.940000 0.825000 ;
      RECT 0.770000  0.825000 0.940000 0.995000 ;
      RECT 0.770000  0.995000 1.065000 1.535000 ;
      RECT 1.070000  1.875000 1.400000 2.635000 ;
      RECT 1.640000  0.255000 1.970000 0.735000 ;
      RECT 1.640000  0.735000 2.915000 0.905000 ;
      RECT 2.195000  0.085000 2.365000 0.555000 ;
      RECT 2.470000  1.535000 3.060000 2.635000 ;
      RECT 2.535000  0.270000 2.915000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21bai_1


MACRO sky130_fd_sc_hdll__xor3_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.660000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.005000 1.075000 8.695000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.735900 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.085000 0.995000 7.305000 1.445000 ;
        RECT 7.085000 1.445000 7.715000 1.725000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 0.995000 2.645000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.472000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.590000 0.925000 ;
        RECT 0.085000 0.925000 0.400000 1.440000 ;
        RECT 0.085000 1.440000 0.610000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.800000  0.695000 1.450000 0.865000 ;
      RECT 0.800000  0.865000 1.000000 1.875000 ;
      RECT 0.800000  1.875000 1.570000 2.045000 ;
      RECT 0.810000  0.085000 1.060000 0.525000 ;
      RECT 0.830000  2.215000 1.165000 2.635000 ;
      RECT 1.230000  0.255000 2.890000 0.425000 ;
      RECT 1.230000  0.425000 1.450000 0.695000 ;
      RECT 1.235000  1.535000 2.985000 1.705000 ;
      RECT 1.350000  2.045000 1.570000 2.235000 ;
      RECT 1.350000  2.235000 3.045000 2.405000 ;
      RECT 1.620000  0.595000 1.790000 1.535000 ;
      RECT 1.970000  1.895000 3.375000 2.065000 ;
      RECT 2.070000  0.655000 3.280000 0.825000 ;
      RECT 2.490000  0.425000 2.890000 0.455000 ;
      RECT 2.815000  0.995000 3.140000 1.325000 ;
      RECT 2.815000  1.325000 2.985000 1.535000 ;
      RECT 3.060000  0.255000 3.960000 0.425000 ;
      RECT 3.060000  0.425000 3.280000 0.655000 ;
      RECT 3.205000  1.525000 3.735000 1.695000 ;
      RECT 3.205000  1.695000 3.375000 1.895000 ;
      RECT 3.310000  2.235000 3.715000 2.405000 ;
      RECT 3.450000  0.595000 3.620000 1.375000 ;
      RECT 3.450000  1.375000 3.735000 1.525000 ;
      RECT 3.545000  1.895000 4.820000 2.065000 ;
      RECT 3.545000  2.065000 3.715000 2.235000 ;
      RECT 3.790000  0.425000 3.960000 1.035000 ;
      RECT 3.790000  1.035000 4.075000 1.205000 ;
      RECT 3.885000  2.235000 4.215000 2.635000 ;
      RECT 3.905000  1.205000 4.075000 1.895000 ;
      RECT 4.130000  0.085000 4.300000 0.865000 ;
      RECT 4.305000  1.445000 4.820000 1.715000 ;
      RECT 4.530000  0.415000 4.820000 1.445000 ;
      RECT 4.650000  2.065000 4.820000 2.275000 ;
      RECT 4.650000  2.275000 7.945000 2.445000 ;
      RECT 4.995000  0.265000 5.410000 0.485000 ;
      RECT 4.995000  0.485000 5.215000 0.595000 ;
      RECT 4.995000  0.595000 5.165000 2.105000 ;
      RECT 5.335000  0.720000 5.800000 0.825000 ;
      RECT 5.335000  0.825000 5.605000 0.890000 ;
      RECT 5.335000  0.890000 5.505000 2.275000 ;
      RECT 5.385000  0.655000 5.800000 0.720000 ;
      RECT 5.630000  0.320000 5.800000 0.655000 ;
      RECT 5.745000  1.445000 6.575000 1.615000 ;
      RECT 5.745000  1.615000 6.160000 2.045000 ;
      RECT 5.760000  0.995000 6.185000 1.270000 ;
      RECT 5.970000  0.630000 6.185000 0.995000 ;
      RECT 6.405000  0.255000 7.600000 0.425000 ;
      RECT 6.405000  0.425000 6.575000 1.445000 ;
      RECT 6.745000  0.595000 6.915000 1.935000 ;
      RECT 6.745000  1.935000 9.565000 2.105000 ;
      RECT 7.085000  0.425000 7.600000 0.465000 ;
      RECT 7.475000  0.730000 7.680000 0.945000 ;
      RECT 7.475000  0.945000 7.785000 1.275000 ;
      RECT 7.935000  1.495000 9.115000 1.705000 ;
      RECT 7.975000  0.295000 8.265000 0.735000 ;
      RECT 7.975000  0.735000 9.115000 0.750000 ;
      RECT 8.015000  0.750000 9.115000 0.905000 ;
      RECT 8.355000  2.275000 9.050000 2.635000 ;
      RECT 8.485000  0.085000 8.935000 0.565000 ;
      RECT 8.945000  0.905000 9.115000 0.995000 ;
      RECT 8.945000  0.995000 9.225000 1.325000 ;
      RECT 8.945000  1.325000 9.115000 1.495000 ;
      RECT 9.030000  1.875000 9.565000 1.935000 ;
      RECT 9.265000  0.255000 9.565000 0.585000 ;
      RECT 9.270000  2.105000 9.565000 2.465000 ;
      RECT 9.395000  0.585000 9.565000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.565000  1.445000 3.735000 1.615000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.535000  0.765000 4.705000 0.935000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.045000  0.425000 5.215000 0.595000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.015000  0.765000 6.185000 0.935000 ;
      RECT 6.015000  1.445000 6.185000 1.615000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.495000  0.765000 7.665000 0.935000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.005000  0.425000 8.175000 0.595000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 3.505000 1.415000 3.795000 1.460000 ;
      RECT 3.505000 1.460000 6.245000 1.600000 ;
      RECT 3.505000 1.600000 3.795000 1.645000 ;
      RECT 4.475000 0.735000 4.765000 0.780000 ;
      RECT 4.475000 0.780000 7.725000 0.920000 ;
      RECT 4.475000 0.920000 4.765000 0.965000 ;
      RECT 4.985000 0.395000 5.275000 0.440000 ;
      RECT 4.985000 0.440000 8.235000 0.580000 ;
      RECT 4.985000 0.580000 5.275000 0.625000 ;
      RECT 5.955000 0.735000 6.245000 0.780000 ;
      RECT 5.955000 0.920000 6.245000 0.965000 ;
      RECT 5.955000 1.415000 6.245000 1.460000 ;
      RECT 5.955000 1.600000 6.245000 1.645000 ;
      RECT 7.435000 0.735000 7.725000 0.780000 ;
      RECT 7.435000 0.920000 7.725000 0.965000 ;
      RECT 7.945000 0.395000 8.235000 0.440000 ;
      RECT 7.945000 0.580000 8.235000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor3_1


MACRO sky130_fd_sc_hdll__xor3_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.660000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.300000 1.075000 8.760000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.735900 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.380000 0.995000 7.600000 1.445000 ;
        RECT 7.380000 1.445000 8.010000 1.665000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.255000 0.995000 2.940000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.517500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.330000 0.660000 0.930000 0.925000 ;
        RECT 0.330000 0.925000 0.695000 1.440000 ;
        RECT 0.330000 1.440000 0.905000 2.045000 ;
        RECT 0.655000 2.045000 0.905000 2.465000 ;
        RECT 0.680000 0.350000 0.930000 0.660000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.105000  0.085000 0.435000 0.465000 ;
      RECT 0.105000  2.215000 0.435000 2.635000 ;
      RECT 1.095000  0.995000 1.295000 1.325000 ;
      RECT 1.105000  0.085000 1.355000 0.525000 ;
      RECT 1.125000  0.695000 1.745000 0.865000 ;
      RECT 1.125000  0.865000 1.295000 0.995000 ;
      RECT 1.125000  1.325000 1.295000 1.875000 ;
      RECT 1.125000  1.875000 1.865000 2.045000 ;
      RECT 1.125000  2.215000 1.460000 2.635000 ;
      RECT 1.525000  0.255000 3.190000 0.425000 ;
      RECT 1.525000  0.425000 1.745000 0.695000 ;
      RECT 1.530000  1.535000 3.280000 1.705000 ;
      RECT 1.645000  2.045000 1.865000 2.235000 ;
      RECT 1.645000  2.235000 3.340000 2.405000 ;
      RECT 1.915000  0.595000 2.085000 1.535000 ;
      RECT 2.265000  1.895000 3.670000 2.065000 ;
      RECT 2.365000  0.655000 3.575000 0.825000 ;
      RECT 2.785000  0.425000 3.190000 0.455000 ;
      RECT 3.110000  0.995000 3.435000 1.325000 ;
      RECT 3.110000  1.325000 3.280000 1.535000 ;
      RECT 3.360000  0.255000 4.255000 0.425000 ;
      RECT 3.360000  0.425000 3.575000 0.655000 ;
      RECT 3.500000  1.525000 4.030000 1.695000 ;
      RECT 3.500000  1.695000 3.670000 1.895000 ;
      RECT 3.605000  2.235000 4.010000 2.405000 ;
      RECT 3.745000  0.595000 3.915000 1.375000 ;
      RECT 3.745000  1.375000 4.030000 1.525000 ;
      RECT 3.840000  1.895000 5.115000 2.065000 ;
      RECT 3.840000  2.065000 4.010000 2.235000 ;
      RECT 4.085000  0.425000 4.255000 1.035000 ;
      RECT 4.085000  1.035000 4.370000 1.205000 ;
      RECT 4.180000  2.235000 4.510000 2.635000 ;
      RECT 4.200000  1.205000 4.370000 1.895000 ;
      RECT 4.425000  0.085000 4.595000 0.865000 ;
      RECT 4.600000  1.445000 5.115000 1.715000 ;
      RECT 4.825000  0.415000 5.115000 1.445000 ;
      RECT 4.945000  2.065000 5.115000 2.275000 ;
      RECT 4.945000  2.275000 8.240000 2.445000 ;
      RECT 5.290000  0.265000 5.705000 0.485000 ;
      RECT 5.290000  0.485000 5.510000 0.595000 ;
      RECT 5.290000  0.595000 5.460000 2.105000 ;
      RECT 5.630000  0.720000 6.095000 0.825000 ;
      RECT 5.630000  0.825000 5.900000 0.890000 ;
      RECT 5.630000  0.890000 5.800000 2.275000 ;
      RECT 5.680000  0.655000 6.095000 0.720000 ;
      RECT 5.925000  0.320000 6.095000 0.655000 ;
      RECT 6.040000  1.445000 6.870000 1.615000 ;
      RECT 6.040000  1.615000 6.455000 2.045000 ;
      RECT 6.055000  0.995000 6.480000 1.270000 ;
      RECT 6.265000  0.630000 6.480000 0.995000 ;
      RECT 6.700000  0.255000 7.895000 0.425000 ;
      RECT 6.700000  0.425000 6.870000 1.445000 ;
      RECT 7.040000  0.595000 7.210000 1.935000 ;
      RECT 7.040000  1.935000 9.550000 2.105000 ;
      RECT 7.380000  0.425000 7.895000 0.465000 ;
      RECT 7.770000  0.730000 7.975000 0.945000 ;
      RECT 7.770000  0.945000 8.090000 1.275000 ;
      RECT 8.230000  1.495000 9.100000 1.705000 ;
      RECT 8.270000  0.295000 8.560000 0.735000 ;
      RECT 8.270000  0.735000 9.100000 0.750000 ;
      RECT 8.310000  0.750000 9.100000 0.905000 ;
      RECT 8.650000  2.275000 9.035000 2.635000 ;
      RECT 8.780000  0.085000 8.950000 0.565000 ;
      RECT 8.930000  0.905000 9.100000 0.995000 ;
      RECT 8.930000  0.995000 9.210000 1.325000 ;
      RECT 8.930000  1.325000 9.100000 1.495000 ;
      RECT 9.015000  1.875000 9.550000 1.935000 ;
      RECT 9.250000  0.255000 9.550000 0.585000 ;
      RECT 9.255000  2.105000 9.550000 2.465000 ;
      RECT 9.380000  0.585000 9.550000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 3.860000  1.445000 4.030000 1.615000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 4.830000  0.765000 5.000000 0.935000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.340000  0.425000 5.510000 0.595000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.310000  0.765000 6.480000 0.935000 ;
      RECT 6.310000  1.445000 6.480000 1.615000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.790000  0.765000 7.960000 0.935000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.300000  0.425000 8.470000 0.595000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 3.800000 1.415000 4.090000 1.460000 ;
      RECT 3.800000 1.460000 6.540000 1.600000 ;
      RECT 3.800000 1.600000 4.090000 1.645000 ;
      RECT 4.770000 0.735000 5.060000 0.780000 ;
      RECT 4.770000 0.780000 8.020000 0.920000 ;
      RECT 4.770000 0.920000 5.060000 0.965000 ;
      RECT 5.280000 0.395000 5.570000 0.440000 ;
      RECT 5.280000 0.440000 8.530000 0.580000 ;
      RECT 5.280000 0.580000 5.570000 0.625000 ;
      RECT 6.250000 0.735000 6.540000 0.780000 ;
      RECT 6.250000 0.920000 6.540000 0.965000 ;
      RECT 6.250000 1.415000 6.540000 1.460000 ;
      RECT 6.250000 1.600000 6.540000 1.645000 ;
      RECT 7.730000 0.735000 8.020000 0.780000 ;
      RECT 7.730000 0.920000 8.020000 0.965000 ;
      RECT 8.240000 0.395000 8.530000 0.440000 ;
      RECT 8.240000 0.580000 8.530000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor3_2


MACRO sky130_fd_sc_hdll__xor3_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.58000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.175000 1.075000 9.635000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.735900 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.255000 0.995000 8.475000 1.445000 ;
        RECT 8.255000 1.445000 8.640000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.130000 0.995000 3.815000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.645000 0.350000 0.815000 0.660000 ;
        RECT 0.645000 0.660000 1.755000 0.925000 ;
        RECT 0.745000 1.440000 1.570000 1.455000 ;
        RECT 0.745000 1.455000 1.855000 2.045000 ;
        RECT 0.745000 2.045000 0.915000 2.465000 ;
        RECT 1.205000 0.925000 1.570000 1.440000 ;
        RECT 1.585000 0.350000 1.755000 0.660000 ;
        RECT 1.685000 2.045000 1.855000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.175000  0.085000  0.345000 0.545000 ;
      RECT  0.275000  2.135000  0.445000 2.635000 ;
      RECT  0.985000  0.085000  1.365000 0.465000 ;
      RECT  1.135000  2.215000  1.465000 2.635000 ;
      RECT  2.020000  0.965000  2.245000 1.325000 ;
      RECT  2.055000  0.085000  2.225000 0.525000 ;
      RECT  2.075000  0.695000  2.565000 0.865000 ;
      RECT  2.075000  0.865000  2.245000 0.965000 ;
      RECT  2.075000  1.325000  2.245000 1.875000 ;
      RECT  2.075000  1.875000  2.795000 2.045000 ;
      RECT  2.075000  2.215000  2.405000 2.635000 ;
      RECT  2.395000  0.255000  4.060000 0.425000 ;
      RECT  2.395000  0.425000  2.565000 0.695000 ;
      RECT  2.570000  1.535000  4.155000 1.705000 ;
      RECT  2.575000  2.045000  2.795000 2.235000 ;
      RECT  2.575000  2.235000  4.215000 2.405000 ;
      RECT  2.790000  0.595000  2.960000 1.535000 ;
      RECT  3.140000  1.895000  4.545000 2.065000 ;
      RECT  3.240000  0.655000  4.450000 0.825000 ;
      RECT  3.660000  0.425000  4.060000 0.455000 ;
      RECT  3.985000  0.995000  4.405000 1.325000 ;
      RECT  3.985000  1.325000  4.155000 1.535000 ;
      RECT  4.230000  0.255000  5.130000 0.425000 ;
      RECT  4.230000  0.425000  4.450000 0.655000 ;
      RECT  4.375000  1.525000  4.905000 1.695000 ;
      RECT  4.375000  1.695000  4.545000 1.895000 ;
      RECT  4.480000  2.235000  4.885000 2.405000 ;
      RECT  4.620000  0.595000  4.790000 1.375000 ;
      RECT  4.620000  1.375000  4.905000 1.525000 ;
      RECT  4.715000  1.895000  5.990000 2.065000 ;
      RECT  4.715000  2.065000  4.885000 2.235000 ;
      RECT  4.960000  0.425000  5.130000 1.035000 ;
      RECT  4.960000  1.035000  5.215000 1.040000 ;
      RECT  4.960000  1.040000  5.230000 1.045000 ;
      RECT  4.960000  1.045000  5.240000 1.050000 ;
      RECT  4.960000  1.050000  5.245000 1.205000 ;
      RECT  5.055000  2.235000  5.385000 2.635000 ;
      RECT  5.075000  1.205000  5.245000 1.895000 ;
      RECT  5.300000  0.085000  5.470000 0.885000 ;
      RECT  5.475000  1.445000  5.990000 1.715000 ;
      RECT  5.700000  0.415000  5.990000 1.445000 ;
      RECT  5.820000  2.065000  5.990000 2.275000 ;
      RECT  5.820000  2.275000  9.115000 2.445000 ;
      RECT  6.165000  0.265000  6.580000 0.485000 ;
      RECT  6.165000  0.485000  6.385000 0.595000 ;
      RECT  6.165000  0.595000  6.335000 2.105000 ;
      RECT  6.525000  0.720000  6.970000 0.825000 ;
      RECT  6.525000  0.825000  6.775000 0.890000 ;
      RECT  6.525000  0.890000  6.695000 2.275000 ;
      RECT  6.555000  0.655000  6.970000 0.720000 ;
      RECT  6.800000  0.320000  6.970000 0.655000 ;
      RECT  6.915000  1.445000  7.745000 1.615000 ;
      RECT  6.915000  1.615000  7.330000 2.045000 ;
      RECT  6.930000  0.995000  7.355000 1.270000 ;
      RECT  7.140000  0.630000  7.355000 0.995000 ;
      RECT  7.575000  0.255000  8.770000 0.425000 ;
      RECT  7.575000  0.425000  7.745000 1.445000 ;
      RECT  7.915000  0.595000  8.085000 1.935000 ;
      RECT  7.915000  1.935000 10.425000 2.105000 ;
      RECT  8.255000  0.425000  8.770000 0.465000 ;
      RECT  8.645000  0.730000  8.850000 0.945000 ;
      RECT  8.645000  0.945000  8.955000 1.275000 ;
      RECT  9.105000  1.495000  9.975000 1.705000 ;
      RECT  9.145000  0.295000  9.435000 0.735000 ;
      RECT  9.145000  0.735000  9.975000 0.750000 ;
      RECT  9.185000  0.750000  9.975000 0.905000 ;
      RECT  9.615000  2.275000  9.945000 2.635000 ;
      RECT  9.695000  0.085000  9.865000 0.565000 ;
      RECT  9.805000  0.905000  9.975000 0.995000 ;
      RECT  9.805000  0.995000 10.035000 1.325000 ;
      RECT  9.805000  1.325000  9.975000 1.495000 ;
      RECT  9.890000  1.875000 10.425000 1.935000 ;
      RECT 10.165000  0.255000 10.425000 0.585000 ;
      RECT 10.165000  2.105000 10.425000 2.465000 ;
      RECT 10.255000  0.585000 10.425000 1.875000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.735000  1.445000  4.905000 1.615000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.705000  0.765000  5.875000 0.935000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.215000  0.425000  6.385000 0.595000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.185000  0.765000  7.355000 0.935000 ;
      RECT  7.185000  1.445000  7.355000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.665000  0.765000  8.835000 0.935000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.175000  0.425000  9.345000 0.595000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 4.675000 1.415000 4.965000 1.460000 ;
      RECT 4.675000 1.460000 7.415000 1.600000 ;
      RECT 4.675000 1.600000 4.965000 1.645000 ;
      RECT 5.645000 0.735000 5.985000 0.780000 ;
      RECT 5.645000 0.780000 8.895000 0.920000 ;
      RECT 5.645000 0.920000 5.985000 0.965000 ;
      RECT 6.155000 0.395000 6.445000 0.440000 ;
      RECT 6.155000 0.440000 9.405000 0.580000 ;
      RECT 6.155000 0.580000 6.445000 0.625000 ;
      RECT 7.125000 0.735000 7.415000 0.780000 ;
      RECT 7.125000 0.920000 7.415000 0.965000 ;
      RECT 7.125000 1.415000 7.415000 1.460000 ;
      RECT 7.125000 1.600000 7.415000 1.645000 ;
      RECT 8.605000 0.735000 8.895000 0.780000 ;
      RECT 8.605000 0.920000 8.895000 0.965000 ;
      RECT 9.115000 0.395000 9.405000 0.440000 ;
      RECT 9.115000 0.580000 9.405000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor3_4


MACRO sky130_fd_sc_hdll__decap_3
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  1.380000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.085000  0.085000 1.295000 0.835000 ;
      RECT 0.085000  0.835000 0.605000 1.375000 ;
      RECT 0.085000  1.545000 1.295000 2.635000 ;
      RECT 0.775000  1.005000 1.295000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__decap_3


MACRO sky130_fd_sc_hdll__decap_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 3.595000 0.855000 ;
      RECT 0.085000  0.855000 1.735000 1.375000 ;
      RECT 0.085000  1.545000 3.595000 2.635000 ;
      RECT 1.905000  1.025000 3.595000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__decap_8


MACRO sky130_fd_sc_hdll__decap_12
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.520000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.085000 5.430000 0.855000 ;
      RECT 0.085000  0.855000 2.665000 1.375000 ;
      RECT 0.085000  1.545000 5.430000 2.635000 ;
      RECT 2.835000  1.025000 5.430000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__decap_12


MACRO sky130_fd_sc_hdll__decap_6
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.085000 2.675000 0.855000 ;
      RECT 0.085000  0.855000 1.295000 1.375000 ;
      RECT 0.085000  1.545000 2.675000 2.635000 ;
      RECT 1.465000  1.025000 2.675000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__decap_6


MACRO sky130_fd_sc_hdll__decap_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  1.840000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.085000 1.755000 0.855000 ;
      RECT 0.085000  0.855000 0.835000 1.375000 ;
      RECT 0.085000  1.545000 1.755000 2.635000 ;
      RECT 1.005000  1.025000 1.755000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__decap_4


MACRO sky130_fd_sc_hdll__nor4_6
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  12.42000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505000 1.075000 2.875000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.325000 1.075000 5.695000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.665000 1.075000 9.035000 1.285000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.395000 1.075000 11.085000 1.285000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.976000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.585000 0.255000  0.915000 0.725000 ;
        RECT  0.585000 0.725000 11.835000 0.905000 ;
        RECT  1.525000 0.255000  1.855000 0.725000 ;
        RECT  2.465000 0.255000  2.795000 0.725000 ;
        RECT  3.405000 0.255000  3.735000 0.725000 ;
        RECT  4.345000 0.255000  4.675000 0.725000 ;
        RECT  5.285000 0.255000  5.615000 0.725000 ;
        RECT  6.745000 0.255000  7.075000 0.725000 ;
        RECT  7.685000 0.255000  8.015000 0.725000 ;
        RECT  8.625000 0.255000  8.955000 0.725000 ;
        RECT  9.565000 0.255000  9.895000 0.725000 ;
        RECT  9.605000 1.455000 11.835000 1.625000 ;
        RECT  9.605000 1.625000  9.855000 2.125000 ;
        RECT 10.505000 0.255000 10.835000 0.725000 ;
        RECT 10.545000 1.625000 10.795000 2.125000 ;
        RECT 11.445000 0.255000 11.835000 0.725000 ;
        RECT 11.445000 0.905000 11.835000 1.455000 ;
        RECT 11.445000 1.625000 11.835000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.115000  0.085000  0.415000 0.905000 ;
      RECT  0.115000  1.455000  3.225000 1.625000 ;
      RECT  0.115000  1.625000  0.405000 2.465000 ;
      RECT  0.625000  1.795000  0.875000 2.635000 ;
      RECT  1.085000  0.085000  1.355000 0.555000 ;
      RECT  1.095000  1.625000  1.345000 2.465000 ;
      RECT  1.565000  1.795000  1.815000 2.635000 ;
      RECT  2.025000  0.085000  2.295000 0.555000 ;
      RECT  2.035000  1.625000  2.285000 2.465000 ;
      RECT  2.505000  1.795000  2.755000 2.635000 ;
      RECT  2.965000  0.085000  3.235000 0.555000 ;
      RECT  2.975000  1.625000  3.225000 2.295000 ;
      RECT  2.975000  2.295000  6.085000 2.465000 ;
      RECT  3.445000  1.455000  8.915000 1.625000 ;
      RECT  3.445000  1.625000  3.695000 2.125000 ;
      RECT  3.905000  0.085000  4.175000 0.555000 ;
      RECT  3.915000  1.795000  4.165000 2.295000 ;
      RECT  4.385000  1.625000  4.635000 2.125000 ;
      RECT  4.845000  0.085000  5.115000 0.555000 ;
      RECT  4.855000  1.795000  5.105000 2.295000 ;
      RECT  5.325000  1.625000  5.575000 2.125000 ;
      RECT  5.785000  0.085000  6.575000 0.555000 ;
      RECT  5.795000  1.795000  6.085000 2.295000 ;
      RECT  6.275000  1.795000  6.565000 2.295000 ;
      RECT  6.275000  2.295000 12.255000 2.465000 ;
      RECT  6.785000  1.625000  7.035000 2.125000 ;
      RECT  7.245000  0.085000  7.515000 0.555000 ;
      RECT  7.255000  1.795000  7.505000 2.295000 ;
      RECT  7.725000  1.625000  7.975000 2.125000 ;
      RECT  8.185000  0.085000  8.455000 0.555000 ;
      RECT  8.195000  1.795000  8.445000 2.295000 ;
      RECT  8.665000  1.625000  8.915000 2.125000 ;
      RECT  9.125000  0.085000  9.395000 0.555000 ;
      RECT  9.135000  1.455000  9.385000 2.295000 ;
      RECT 10.065000  0.085000 10.335000 0.555000 ;
      RECT 10.075000  1.795000 10.325000 2.295000 ;
      RECT 11.005000  0.085000 11.275000 0.555000 ;
      RECT 11.015000  1.795000 11.265000 2.295000 ;
      RECT 12.005000  0.085000 12.255000 0.905000 ;
      RECT 12.005000  1.455000 12.255000 2.295000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_6


MACRO sky130_fd_sc_hdll__nor4_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.740000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.180000 1.075000 2.025000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 1.075000 4.470000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.695000 1.075000 6.305000 1.285000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.475000 1.075000 8.045000 1.285000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.374000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 8.630000 0.905000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 2.415000 0.255000 2.795000 0.725000 ;
        RECT 3.355000 0.255000 3.735000 0.725000 ;
        RECT 4.815000 0.255000 5.195000 0.725000 ;
        RECT 5.755000 0.255000 6.135000 0.725000 ;
        RECT 6.695000 0.255000 7.075000 0.725000 ;
        RECT 6.785000 1.455000 8.630000 1.625000 ;
        RECT 6.785000 1.625000 7.035000 2.125000 ;
        RECT 7.635000 0.255000 8.015000 0.725000 ;
        RECT 7.725000 1.625000 7.975000 2.125000 ;
        RECT 8.360000 0.905000 8.630000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 2.285000 1.625000 ;
      RECT 0.090000  1.625000 0.405000 2.465000 ;
      RECT 0.625000  1.795000 0.875000 2.635000 ;
      RECT 1.095000  1.625000 1.345000 2.465000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 1.565000  1.795000 1.815000 2.635000 ;
      RECT 2.035000  1.625000 2.285000 2.295000 ;
      RECT 2.035000  2.295000 4.220000 2.465000 ;
      RECT 2.075000  0.085000 2.245000 0.555000 ;
      RECT 2.505000  1.455000 6.095000 1.625000 ;
      RECT 2.505000  1.625000 2.755000 2.125000 ;
      RECT 2.975000  1.795000 3.225000 2.295000 ;
      RECT 3.015000  0.085000 3.185000 0.555000 ;
      RECT 3.445000  1.625000 3.695000 2.125000 ;
      RECT 3.915000  1.795000 4.220000 2.295000 ;
      RECT 3.955000  0.085000 4.645000 0.555000 ;
      RECT 4.405000  1.795000 4.685000 2.295000 ;
      RECT 4.405000  2.295000 8.445000 2.465000 ;
      RECT 4.905000  1.625000 5.155000 2.125000 ;
      RECT 5.375000  1.795000 5.625000 2.295000 ;
      RECT 5.415000  0.085000 5.585000 0.555000 ;
      RECT 5.845000  1.625000 6.095000 2.125000 ;
      RECT 6.315000  1.795000 6.565000 2.295000 ;
      RECT 6.355000  0.085000 6.525000 0.555000 ;
      RECT 7.255000  1.795000 7.505000 2.295000 ;
      RECT 7.295000  0.085000 7.465000 0.555000 ;
      RECT 8.195000  1.795000 8.445000 2.295000 ;
      RECT 8.235000  0.085000 8.405000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_4


MACRO sky130_fd_sc_hdll__nor4_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.655000 2.205000 1.665000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.995000 1.745000 2.450000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 0.995000 1.285000 2.450000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.745000 0.335000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.699000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.495000 0.775000 1.665000 ;
        RECT 0.090000 1.665000 0.425000 2.450000 ;
        RECT 0.515000 0.385000 0.815000 0.655000 ;
        RECT 0.515000 0.655000 1.765000 0.825000 ;
        RECT 0.515000 0.825000 0.775000 1.495000 ;
        RECT 1.595000 0.385000 1.765000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.575000 ;
      RECT 1.035000  0.085000 1.365000 0.485000 ;
      RECT 2.005000  0.085000 2.520000 0.485000 ;
      RECT 2.135000  1.835000 2.535000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_1


MACRO sky130_fd_sc_hdll__nor4_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  16.10000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.405000 1.075000 3.795000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.245000 1.075000 7.635000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.445000 1.075000 11.835000 1.285000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.985000 1.075000 15.355000 1.285000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  3.968000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.565000 0.255000  0.895000 0.725000 ;
        RECT  0.565000 0.725000 15.515000 0.905000 ;
        RECT  1.505000 0.255000  1.835000 0.725000 ;
        RECT  2.445000 0.255000  2.775000 0.725000 ;
        RECT  3.385000 0.255000  3.715000 0.725000 ;
        RECT  4.325000 0.255000  4.655000 0.725000 ;
        RECT  5.265000 0.255000  5.595000 0.725000 ;
        RECT  6.205000 0.255000  6.535000 0.725000 ;
        RECT  7.145000 0.255000  7.475000 0.725000 ;
        RECT  8.605000 0.255000  8.935000 0.725000 ;
        RECT  9.545000 0.255000  9.875000 0.725000 ;
        RECT 10.485000 0.255000 10.815000 0.725000 ;
        RECT 11.425000 0.255000 11.755000 0.725000 ;
        RECT 12.365000 0.255000 12.695000 0.725000 ;
        RECT 12.405000 0.905000 12.815000 1.455000 ;
        RECT 12.405000 1.455000 15.475000 1.625000 ;
        RECT 12.405000 1.625000 12.655000 2.125000 ;
        RECT 13.305000 0.255000 13.635000 0.725000 ;
        RECT 13.345000 1.625000 13.595000 2.125000 ;
        RECT 14.245000 0.255000 14.575000 0.725000 ;
        RECT 14.285000 1.625000 14.535000 2.125000 ;
        RECT 15.185000 0.255000 15.515000 0.725000 ;
        RECT 15.225000 1.625000 15.475000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 16.100000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 16.100000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.100000 0.085000 ;
      RECT  0.000000  2.635000 16.100000 2.805000 ;
      RECT  0.095000  1.455000  4.145000 1.625000 ;
      RECT  0.095000  1.625000  0.425000 2.465000 ;
      RECT  0.135000  0.085000  0.395000 0.905000 ;
      RECT  0.605000  1.795000  0.855000 2.635000 ;
      RECT  1.065000  0.085000  1.335000 0.555000 ;
      RECT  1.075000  1.625000  1.325000 2.465000 ;
      RECT  1.545000  1.795000  1.795000 2.635000 ;
      RECT  2.005000  0.085000  2.275000 0.555000 ;
      RECT  2.015000  1.625000  2.265000 2.465000 ;
      RECT  2.485000  1.795000  2.735000 2.635000 ;
      RECT  2.945000  0.085000  3.215000 0.555000 ;
      RECT  2.955000  1.625000  3.205000 2.465000 ;
      RECT  3.425000  1.795000  3.675000 2.635000 ;
      RECT  3.885000  0.085000  4.155000 0.555000 ;
      RECT  3.895000  1.625000  4.145000 2.295000 ;
      RECT  3.895000  2.295000  7.945000 2.465000 ;
      RECT  4.365000  1.455000 11.715000 1.625000 ;
      RECT  4.365000  1.625000  4.615000 2.125000 ;
      RECT  4.825000  0.085000  5.095000 0.555000 ;
      RECT  4.835000  1.795000  5.085000 2.295000 ;
      RECT  5.305000  1.625000  5.555000 2.125000 ;
      RECT  5.765000  0.085000  6.035000 0.555000 ;
      RECT  5.775000  1.795000  6.025000 2.295000 ;
      RECT  6.245000  1.625000  6.495000 2.125000 ;
      RECT  6.705000  0.085000  6.975000 0.555000 ;
      RECT  6.715000  1.795000  6.965000 2.295000 ;
      RECT  7.185000  1.625000  7.435000 2.125000 ;
      RECT  7.645000  0.085000  8.435000 0.555000 ;
      RECT  7.655000  1.795000  7.945000 2.295000 ;
      RECT  8.135000  1.795000  8.425000 2.295000 ;
      RECT  8.135000  2.295000 15.995000 2.465000 ;
      RECT  8.645000  1.625000  8.895000 2.125000 ;
      RECT  9.075000  1.795000  9.365000 2.295000 ;
      RECT  9.105000  0.085000  9.375000 0.555000 ;
      RECT  9.585000  1.625000  9.835000 2.125000 ;
      RECT 10.045000  0.085000 10.315000 0.555000 ;
      RECT 10.055000  1.795000 10.305000 2.295000 ;
      RECT 10.525000  1.625000 10.775000 2.125000 ;
      RECT 10.985000  0.085000 11.255000 0.555000 ;
      RECT 10.995000  1.795000 11.245000 2.295000 ;
      RECT 11.465000  1.625000 11.715000 2.125000 ;
      RECT 11.925000  0.085000 12.195000 0.555000 ;
      RECT 11.935000  1.455000 12.185000 2.295000 ;
      RECT 12.865000  0.085000 13.135000 0.555000 ;
      RECT 12.875000  1.795000 13.125000 2.295000 ;
      RECT 13.805000  0.085000 14.075000 0.555000 ;
      RECT 13.815000  1.795000 14.065000 2.295000 ;
      RECT 14.745000  0.085000 15.015000 0.555000 ;
      RECT 14.755000  1.795000 15.005000 2.295000 ;
      RECT 15.685000  0.085000 15.965000 0.905000 ;
      RECT 15.695000  1.465000 15.995000 2.295000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_8


MACRO sky130_fd_sc_hdll__nor4_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.200000 1.075000 1.015000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.235000 1.075000 2.140000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.410000 1.075000 3.355000 1.285000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.640000 1.075000 4.275000 1.285000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.252000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.570000 0.255000 0.950000 0.725000 ;
        RECT 0.570000 0.725000 4.950000 0.905000 ;
        RECT 1.510000 0.255000 1.890000 0.725000 ;
        RECT 3.010000 0.255000 3.390000 0.725000 ;
        RECT 3.950000 0.255000 4.330000 0.725000 ;
        RECT 4.040000 1.455000 4.950000 1.625000 ;
        RECT 4.040000 1.625000 4.290000 2.125000 ;
        RECT 4.615000 0.905000 4.950000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.150000  1.455000 2.285000 1.625000 ;
      RECT 0.150000  1.625000 0.405000 2.465000 ;
      RECT 0.625000  1.795000 0.875000 2.635000 ;
      RECT 1.095000  1.625000 1.345000 2.465000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 1.565000  1.795000 1.815000 2.295000 ;
      RECT 1.565000  2.295000 3.315000 2.465000 ;
      RECT 2.035000  1.625000 2.285000 2.125000 ;
      RECT 2.075000  0.085000 2.805000 0.555000 ;
      RECT 2.595000  1.455000 3.785000 1.625000 ;
      RECT 2.595000  1.625000 2.845000 2.125000 ;
      RECT 3.065000  1.795000 3.315000 2.295000 ;
      RECT 3.535000  1.625000 3.785000 2.295000 ;
      RECT 3.535000  2.295000 4.725000 2.465000 ;
      RECT 3.575000  0.085000 3.745000 0.555000 ;
      RECT 4.475000  1.795000 4.725000 2.295000 ;
      RECT 4.515000  0.085000 4.805000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_2


MACRO sky130_fd_sc_hdll__a22o_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.675000 1.820000 1.075000 ;
        RECT 1.525000 1.075000 1.940000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.160000 1.075000 2.615000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.815000 1.075000 1.340000 1.285000 ;
        RECT 1.065000 0.675000 1.340000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.625000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.150000 0.255000 3.560000 0.585000 ;
        RECT 3.150000 1.785000 3.560000 2.465000 ;
        RECT 3.240000 0.585000 3.560000 1.785000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.095000  0.085000 0.595000 0.850000 ;
      RECT 0.095000  1.455000 3.015000 1.625000 ;
      RECT 0.095000  1.625000 0.425000 2.295000 ;
      RECT 0.095000  2.295000 1.365000 2.465000 ;
      RECT 0.645000  1.795000 2.380000 2.035000 ;
      RECT 0.645000  2.035000 0.875000 2.125000 ;
      RECT 0.870000  0.255000 2.295000 0.505000 ;
      RECT 1.035000  2.255000 1.365000 2.295000 ;
      RECT 1.555000  2.215000 1.910000 2.635000 ;
      RECT 2.125000  0.505000 2.295000 0.735000 ;
      RECT 2.125000  0.735000 3.015000 0.905000 ;
      RECT 2.130000  2.035000 2.380000 2.465000 ;
      RECT 2.505000  0.085000 2.885000 0.565000 ;
      RECT 2.600000  1.875000 2.930000 2.635000 ;
      RECT 2.845000  0.905000 3.015000 1.455000 ;
      RECT 3.755000  0.085000 3.925000 0.985000 ;
      RECT 3.755000  1.445000 3.925000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22o_2


MACRO sky130_fd_sc_hdll__a22o_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.675000 1.745000 1.065000 ;
        RECT 1.525000 1.065000 2.085000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275000 0.980000 2.625000 1.285000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.815000 1.075000 1.285000 1.285000 ;
        RECT 1.065000 0.675000 1.285000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.625000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.670000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.275000 0.255000 3.535000 0.585000 ;
        RECT 3.275000 1.785000 3.535000 2.465000 ;
        RECT 3.365000 0.585000 3.535000 1.785000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.085000 0.595000 0.850000 ;
      RECT 0.090000  1.495000 3.035000 1.715000 ;
      RECT 0.090000  1.715000 0.345000 2.245000 ;
      RECT 0.090000  2.245000 0.425000 2.465000 ;
      RECT 0.565000  1.885000 2.395000 2.085000 ;
      RECT 0.870000  0.255000 2.280000 0.465000 ;
      RECT 1.540000  2.255000 1.895000 2.635000 ;
      RECT 2.065000  2.085000 2.395000 2.465000 ;
      RECT 2.110000  0.465000 2.280000 0.615000 ;
      RECT 2.110000  0.615000 3.035000 0.785000 ;
      RECT 2.585000  0.085000 2.915000 0.445000 ;
      RECT 2.585000  1.935000 2.915000 2.635000 ;
      RECT 2.865000  0.785000 3.035000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22o_1


MACRO sky130_fd_sc_hdll__a22o_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.900000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.350000 1.075000 5.895000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.750000 1.075000 5.130000 1.445000 ;
        RECT 4.750000 1.445000 6.285000 1.615000 ;
        RECT 6.115000 1.075000 6.815000 1.275000 ;
        RECT 6.115000 1.275000 6.285000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375000 1.075000 4.030000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.620000 1.075000 3.205000 1.445000 ;
        RECT 2.620000 1.445000 4.580000 1.615000 ;
        RECT 4.200000 1.075000 4.580000 1.445000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.725000 1.920000 0.905000 ;
        RECT 0.085000 0.905000 0.370000 1.445000 ;
        RECT 0.085000 1.445000 1.880000 1.615000 ;
        RECT 0.600000 0.265000 0.980000 0.725000 ;
        RECT 0.690000 1.615000 0.940000 2.465000 ;
        RECT 1.540000 0.255000 1.920000 0.725000 ;
        RECT 1.630000 1.615000 1.880000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.220000  1.825000 0.470000 2.635000 ;
      RECT 0.260000  0.085000 0.430000 0.555000 ;
      RECT 0.540000  1.075000 2.430000 1.275000 ;
      RECT 1.160000  1.795000 1.410000 2.635000 ;
      RECT 1.200000  0.085000 1.370000 0.555000 ;
      RECT 2.100000  1.275000 2.430000 1.785000 ;
      RECT 2.100000  1.785000 4.280000 1.955000 ;
      RECT 2.100000  2.125000 2.350000 2.635000 ;
      RECT 2.140000  0.085000 2.830000 0.555000 ;
      RECT 2.140000  0.735000 5.810000 0.905000 ;
      RECT 2.140000  0.905000 2.430000 1.075000 ;
      RECT 2.620000  2.125000 2.870000 2.295000 ;
      RECT 2.620000  2.295000 4.830000 2.465000 ;
      RECT 3.000000  0.255000 4.320000 0.475000 ;
      RECT 3.090000  1.955000 3.340000 2.125000 ;
      RECT 3.420000  0.645000 3.905000 0.735000 ;
      RECT 3.560000  2.125000 3.810000 2.295000 ;
      RECT 4.030000  1.955000 4.280000 2.125000 ;
      RECT 4.500000  1.785000 6.710000 1.955000 ;
      RECT 4.500000  1.955000 4.830000 2.295000 ;
      RECT 4.585000  0.085000 4.755000 0.555000 ;
      RECT 4.960000  0.255000 6.280000 0.475000 ;
      RECT 5.050000  2.125000 5.300000 2.635000 ;
      RECT 5.385000  0.645000 5.810000 0.735000 ;
      RECT 5.520000  1.955000 5.770000 2.465000 ;
      RECT 5.990000  2.125000 6.240000 2.635000 ;
      RECT 6.030000  0.475000 6.280000 0.895000 ;
      RECT 6.500000  0.085000 6.670000 0.895000 ;
      RECT 6.505000  1.455000 6.710000 1.785000 ;
      RECT 6.505000  1.955000 6.710000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22o_4


MACRO sky130_fd_sc_hdll__inputiso1p_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.440000 1.325000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.765000 1.315000 1.325000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.650500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.665000 0.255000 2.215000 0.825000 ;
        RECT 1.795000 1.845000 2.215000 2.465000 ;
        RECT 1.900000 0.825000 2.215000 1.845000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.150000  1.495000 1.705000 1.665000 ;
      RECT 0.150000  1.665000 0.540000 1.840000 ;
      RECT 0.190000  0.085000 0.430000 0.595000 ;
      RECT 0.610000  0.265000 0.940000 0.595000 ;
      RECT 0.610000  0.595000 0.830000 1.495000 ;
      RECT 1.185000  1.835000 1.515000 2.635000 ;
      RECT 1.220000  0.085000 1.435000 0.595000 ;
      RECT 1.535000  0.995000 1.705000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inputiso1p_1


MACRO sky130_fd_sc_hdll__a221oi_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.675000 2.350000 1.075000 ;
        RECT 1.985000 1.075000 2.425000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.670000 0.995000 3.075000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.325000 1.075000 1.815000 1.285000 ;
        RECT 1.525000 0.675000 1.815000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.075000 1.155000 1.285000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.435000 1.285000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.874500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.170000 0.255000 0.345000 0.735000 ;
        RECT 0.170000 0.735000 1.335000 0.905000 ;
        RECT 0.175000 1.455000 2.450000 1.495000 ;
        RECT 0.175000 1.495000 3.535000 1.625000 ;
        RECT 0.175000 1.625000 0.345000 2.465000 ;
        RECT 1.165000 0.255000 2.780000 0.505000 ;
        RECT 1.165000 0.505000 1.335000 0.735000 ;
        RECT 2.300000 1.625000 3.535000 1.665000 ;
        RECT 2.580000 0.505000 2.780000 0.655000 ;
        RECT 2.580000 0.655000 3.535000 0.825000 ;
        RECT 3.255000 0.825000 3.535000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.515000  0.085000 0.895000 0.565000 ;
      RECT 0.515000  1.795000 0.815000 2.295000 ;
      RECT 0.515000  2.295000 1.835000 2.465000 ;
      RECT 1.115000  1.795000 2.175000 1.835000 ;
      RECT 1.115000  1.835000 2.825000 2.045000 ;
      RECT 1.115000  2.045000 1.340000 2.125000 ;
      RECT 1.455000  2.255000 1.835000 2.295000 ;
      RECT 2.025000  2.215000 2.355000 2.635000 ;
      RECT 2.575000  2.045000 2.825000 2.465000 ;
      RECT 3.030000  0.085000 3.360000 0.485000 ;
      RECT 3.045000  1.875000 3.375000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a221oi_1


MACRO sky130_fd_sc_hdll__a221oi_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.58000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.145000 1.075000 8.755000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.585000 1.075000  6.965000 1.445000 ;
        RECT 6.585000 1.445000  9.135000 1.615000 ;
        RECT 8.965000 1.075000 10.400000 1.275000 ;
        RECT 8.965000 1.275000  9.135000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.335000 0.995000 5.885000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 0.995000 4.165000 1.325000 ;
        RECT 3.945000 1.325000 4.165000 1.445000 ;
        RECT 3.945000 1.445000 6.410000 1.615000 ;
        RECT 6.065000 1.075000 6.410000 1.445000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.435000 1.275000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.893000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 1.855000 0.905000 ;
        RECT 0.625000 1.445000 1.855000 1.615000 ;
        RECT 0.625000 1.615000 0.875000 2.125000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 1.565000 1.615000 1.815000 2.125000 ;
        RECT 1.655000 0.905000 1.855000 1.095000 ;
        RECT 1.655000 1.095000 3.595000 1.275000 ;
        RECT 1.655000 1.275000 1.855000 1.445000 ;
        RECT 3.375000 0.645000 6.280000 0.735000 ;
        RECT 3.375000 0.735000 8.585000 0.820000 ;
        RECT 3.375000 0.820000 3.595000 1.095000 ;
        RECT 6.110000 0.820000 7.130000 0.905000 ;
        RECT 6.960000 0.645000 8.585000 0.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.090000  1.445000  0.405000 2.295000 ;
      RECT  0.090000  2.295000  2.325000 2.465000 ;
      RECT  0.115000  0.085000  0.365000 0.895000 ;
      RECT  1.095000  1.785000  1.345000 2.295000 ;
      RECT  1.135000  0.085000  1.305000 0.555000 ;
      RECT  2.075000  0.085000  2.245000 0.645000 ;
      RECT  2.075000  0.645000  3.205000 0.925000 ;
      RECT  2.075000  1.445000  3.330000 1.615000 ;
      RECT  2.075000  1.615000  2.325000 2.295000 ;
      RECT  2.435000  0.255000  6.185000 0.425000 ;
      RECT  2.435000  0.425000  2.860000 0.475000 ;
      RECT  2.565000  1.795000  2.815000 2.215000 ;
      RECT  2.565000  2.215000  6.655000 2.465000 ;
      RECT  3.035000  0.595000  3.205000 0.645000 ;
      RECT  3.035000  1.615000  3.330000 1.835000 ;
      RECT  3.035000  1.835000  6.185000 2.045000 ;
      RECT  3.335000  0.425000  6.185000 0.475000 ;
      RECT  6.405000  1.785000  9.525000 2.045000 ;
      RECT  6.405000  2.045000  6.655000 2.215000 ;
      RECT  6.455000  0.085000  6.625000 0.555000 ;
      RECT  6.795000  0.255000  9.055000 0.475000 ;
      RECT  6.825000  2.215000  9.085000 2.635000 ;
      RECT  8.805000  0.475000  9.055000 0.725000 ;
      RECT  8.805000  0.725000  9.995000 0.905000 ;
      RECT  9.275000  0.085000  9.445000 0.555000 ;
      RECT  9.275000  2.045000  9.445000 2.465000 ;
      RECT  9.355000  1.445000 10.425000 1.615000 ;
      RECT  9.355000  1.615000  9.525000 1.785000 ;
      RECT  9.615000  0.255000  9.995000 0.725000 ;
      RECT  9.745000  1.795000  9.915000 2.635000 ;
      RECT 10.165000  0.085000 10.335000 0.905000 ;
      RECT 10.175000  1.615000 10.425000 2.465000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a221oi_4


MACRO sky130_fd_sc_hdll__a221oi_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.235000 1.075000 4.915000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.735000 1.075000 4.065000 1.445000 ;
        RECT 3.735000 1.445000 5.270000 1.615000 ;
        RECT 5.100000 1.075000 5.885000 1.275000 ;
        RECT 5.100000 1.275000 5.270000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.360000 1.075000 3.015000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.730000 1.075000 2.190000 1.445000 ;
        RECT 1.730000 1.445000 3.565000 1.615000 ;
        RECT 3.185000 1.075000 3.565000 1.445000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.420000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.979000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 0.305000 0.905000 0.725000 ;
        RECT 0.525000 0.725000 4.795000 0.865000 ;
        RECT 0.605000 0.865000 4.795000 0.905000 ;
        RECT 0.605000 0.905000 0.905000 2.125000 ;
        RECT 2.435000 0.645000 2.835000 0.725000 ;
        RECT 4.415000 0.645000 4.795000 0.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.090000  1.795000 0.435000 2.295000 ;
      RECT 0.090000  2.295000 1.375000 2.465000 ;
      RECT 0.105000  0.085000 0.355000 0.895000 ;
      RECT 1.125000  0.085000 1.815000 0.555000 ;
      RECT 1.125000  1.495000 1.375000 1.785000 ;
      RECT 1.125000  1.785000 3.265000 1.955000 ;
      RECT 1.125000  1.955000 1.375000 2.295000 ;
      RECT 1.605000  2.125000 1.855000 2.295000 ;
      RECT 1.605000  2.295000 3.775000 2.465000 ;
      RECT 1.985000  0.255000 3.305000 0.475000 ;
      RECT 2.075000  1.955000 2.325000 2.125000 ;
      RECT 2.545000  2.125000 2.795000 2.295000 ;
      RECT 3.015000  1.955000 3.265000 2.125000 ;
      RECT 3.525000  1.785000 5.695000 1.955000 ;
      RECT 3.525000  1.955000 3.775000 2.295000 ;
      RECT 3.570000  0.085000 3.740000 0.555000 ;
      RECT 3.945000  0.255000 5.265000 0.475000 ;
      RECT 4.035000  2.125000 4.285000 2.635000 ;
      RECT 4.505000  1.955000 4.755000 2.465000 ;
      RECT 4.975000  2.125000 5.225000 2.635000 ;
      RECT 5.015000  0.475000 5.265000 0.905000 ;
      RECT 5.485000  0.085000 5.655000 0.905000 ;
      RECT 5.490000  1.455000 5.695000 1.785000 ;
      RECT 5.490000  1.955000 5.695000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a221oi_2


MACRO sky130_fd_sc_hdll__xnor2_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.980000 1.075000 1.775000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.810000 1.445000 ;
        RECT 0.425000 1.445000 2.165000 1.615000 ;
        RECT 1.945000 1.075000 2.645000 1.245000 ;
        RECT 1.945000 1.245000 2.165000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.545000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515000 2.125000 2.895000 2.295000 ;
        RECT 2.725000 1.755000 3.595000 1.955000 ;
        RECT 2.725000 1.955000 2.895000 2.125000 ;
        RECT 3.175000 0.345000 3.595000 0.825000 ;
        RECT 3.355000 0.825000 3.595000 1.755000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.280000 0.550000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.785000 ;
      RECT 0.085000  1.785000 2.555000 1.955000 ;
      RECT 0.085000  2.125000 0.385000 2.635000 ;
      RECT 0.555000  1.955000 0.935000 2.465000 ;
      RECT 1.155000  0.085000 1.325000 0.905000 ;
      RECT 1.155000  2.125000 1.835000 2.635000 ;
      RECT 1.495000  0.255000 1.875000 0.655000 ;
      RECT 1.495000  0.655000 2.895000 0.825000 ;
      RECT 2.095000  0.085000 2.495000 0.475000 ;
      RECT 2.335000  1.415000 3.095000 1.585000 ;
      RECT 2.335000  1.585000 2.555000 1.785000 ;
      RECT 2.665000  0.255000 2.895000 0.655000 ;
      RECT 2.875000  0.995000 3.095000 1.415000 ;
      RECT 3.115000  2.125000 3.415000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor2_1


MACRO sky130_fd_sc_hdll__xnor2_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.075000 2.905000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485000 1.075000 1.010000 1.285000 ;
        RECT 0.840000 1.285000 1.010000 1.445000 ;
        RECT 0.840000 1.445000 3.350000 1.615000 ;
        RECT 3.180000 1.075000 4.305000 1.285000 ;
        RECT 3.180000 1.285000 3.350000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.953000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.075000 1.795000 5.745000 1.965000 ;
        RECT 4.075000 1.965000 4.285000 2.125000 ;
        RECT 4.985000 0.305000 6.340000 0.475000 ;
        RECT 5.495000 1.415000 6.340000 1.625000 ;
        RECT 5.495000 1.625000 5.745000 1.795000 ;
        RECT 5.495000 1.965000 5.745000 2.125000 ;
        RECT 5.950000 0.475000 6.340000 1.415000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  0.645000 0.910000 0.895000 ;
      RECT 0.085000  0.895000 0.315000 1.785000 ;
      RECT 0.085000  1.785000 3.780000 1.955000 ;
      RECT 0.085000  1.955000 2.280000 1.965000 ;
      RECT 0.085000  1.965000 0.400000 2.465000 ;
      RECT 0.105000  0.255000 1.380000 0.475000 ;
      RECT 0.620000  2.135000 0.870000 2.635000 ;
      RECT 1.090000  1.965000 1.340000 2.465000 ;
      RECT 1.130000  0.475000 1.380000 0.725000 ;
      RECT 1.130000  0.725000 2.320000 0.905000 ;
      RECT 1.560000  2.135000 1.810000 2.635000 ;
      RECT 1.600000  0.085000 1.770000 0.555000 ;
      RECT 1.940000  0.255000 2.320000 0.725000 ;
      RECT 2.030000  1.965000 2.280000 2.465000 ;
      RECT 2.590000  2.125000 2.840000 2.465000 ;
      RECT 2.630000  0.085000 2.800000 0.905000 ;
      RECT 2.970000  0.255000 3.350000 0.725000 ;
      RECT 2.970000  0.725000 5.755000 0.905000 ;
      RECT 3.060000  2.135000 3.310000 2.635000 ;
      RECT 3.530000  2.125000 3.855000 2.295000 ;
      RECT 3.530000  2.295000 4.755000 2.465000 ;
      RECT 3.570000  0.085000 3.740000 0.555000 ;
      RECT 3.610000  1.455000 5.205000 1.625000 ;
      RECT 3.610000  1.625000 3.780000 1.785000 ;
      RECT 3.910000  0.255000 4.325000 0.725000 ;
      RECT 4.505000  2.135000 4.755000 2.295000 ;
      RECT 4.545000  0.085000 4.715000 0.555000 ;
      RECT 5.025000  2.135000 5.275000 2.635000 ;
      RECT 5.035000  1.075000 5.745000 1.245000 ;
      RECT 5.035000  1.245000 5.205000 1.455000 ;
      RECT 5.405000  0.645000 5.755000 0.725000 ;
      RECT 5.965000  1.795000 6.340000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.665000  2.125000 2.835000 2.295000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.685000  2.125000 3.855000 2.295000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 2.605000 2.095000 2.895000 2.140000 ;
      RECT 2.605000 2.140000 3.915000 2.280000 ;
      RECT 2.605000 2.280000 2.895000 2.325000 ;
      RECT 3.625000 2.095000 3.915000 2.140000 ;
      RECT 3.625000 2.280000 3.915000 2.325000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor2_2


MACRO sky130_fd_sc_hdll__xnor2_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.04000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 1.075000 5.930000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 1.075000 2.005000 1.275000 ;
        RECT 1.835000 1.275000 2.005000 1.445000 ;
        RECT 1.835000 1.445000 6.270000 1.615000 ;
        RECT 6.100000 1.075000 8.170000 1.275000 ;
        RECT 6.100000 1.275000 6.270000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.858500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  6.750000 1.785000  9.060000 2.045000 ;
        RECT  8.730000 1.445000 10.940000 1.665000 ;
        RECT  8.730000 1.665000  9.060000 1.785000 ;
        RECT  8.730000 2.045000  9.060000 2.465000 ;
        RECT  9.150000 0.655000 10.940000 0.905000 ;
        RECT  9.710000 1.665000  9.960000 2.465000 ;
        RECT 10.610000 1.665000 10.940000 2.465000 ;
        RECT 10.705000 0.905000 10.940000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.085000  0.645000  1.910000 0.905000 ;
      RECT  0.085000  0.905000  0.320000 1.445000 ;
      RECT  0.085000  1.445000  1.400000 1.615000 ;
      RECT  0.085000  1.615000  0.460000 2.465000 ;
      RECT  0.170000  0.255000  2.380000 0.475000 ;
      RECT  0.680000  1.835000  0.930000 2.635000 ;
      RECT  1.150000  1.615000  1.400000 1.785000 ;
      RECT  1.150000  1.785000  4.220000 2.005000 ;
      RECT  1.150000  2.005000  1.400000 2.465000 ;
      RECT  1.620000  2.175000  1.870000 2.635000 ;
      RECT  2.090000  2.005000  2.340000 2.465000 ;
      RECT  2.130000  0.475000  2.380000 0.725000 ;
      RECT  2.130000  0.725000  4.260000 0.905000 ;
      RECT  2.560000  2.175000  2.810000 2.635000 ;
      RECT  2.600000  0.085000  2.770000 0.555000 ;
      RECT  2.940000  0.255000  3.320000 0.725000 ;
      RECT  3.030000  2.005000  3.280000 2.465000 ;
      RECT  3.500000  2.175000  3.750000 2.635000 ;
      RECT  3.540000  0.085000  3.710000 0.555000 ;
      RECT  3.880000  0.255000  4.260000 0.725000 ;
      RECT  3.970000  2.005000  4.220000 2.465000 ;
      RECT  4.425000  1.785000  6.580000 2.005000 ;
      RECT  4.425000  2.005000  4.740000 2.465000 ;
      RECT  4.430000  0.085000  4.700000 0.905000 ;
      RECT  4.870000  0.255000  5.250000 0.725000 ;
      RECT  4.870000  0.725000  8.170000 0.735000 ;
      RECT  4.870000  0.735000  8.980000 0.905000 ;
      RECT  4.960000  2.175000  5.210000 2.635000 ;
      RECT  5.430000  2.005000  5.680000 2.465000 ;
      RECT  5.470000  0.085000  5.640000 0.555000 ;
      RECT  5.810000  0.255000  6.190000 0.725000 ;
      RECT  5.900000  2.175000  6.150000 2.635000 ;
      RECT  6.370000  2.005000  6.580000 2.215000 ;
      RECT  6.370000  2.215000  8.540000 2.465000 ;
      RECT  6.410000  0.085000  6.580000 0.555000 ;
      RECT  6.490000  1.445000  8.560000 1.615000 ;
      RECT  6.750000  0.255000  7.130000 0.725000 ;
      RECT  7.350000  0.085000  7.520000 0.555000 ;
      RECT  7.690000  0.255000  8.070000 0.725000 ;
      RECT  8.290000  0.085000  8.460000 0.555000 ;
      RECT  8.390000  1.075000 10.535000 1.275000 ;
      RECT  8.390000  1.275000  8.560000 1.445000 ;
      RECT  8.730000  0.305000 10.940000 0.475000 ;
      RECT  8.730000  0.475000  8.980000 0.735000 ;
      RECT  9.240000  1.835000  9.490000 2.635000 ;
      RECT 10.180000  1.835000 10.430000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.165000  1.445000  1.335000 1.615000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.725000  1.445000  6.895000 1.615000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 1.055000 1.415000 1.395000 1.460000 ;
      RECT 1.055000 1.460000 7.005000 1.600000 ;
      RECT 1.055000 1.600000 1.395000 1.645000 ;
      RECT 6.655000 1.415000 7.005000 1.460000 ;
      RECT 6.655000 1.600000 7.005000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor2_4


MACRO sky130_fd_sc_hdll__o21a_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.275000 0.995000 3.535000 1.450000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.320000 1.025000 3.075000 1.400000 ;
        RECT 2.800000 1.400000 3.075000 1.985000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.010000 1.955000 1.615000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.506200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 0.255000 0.825000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  1.635000 0.345000 2.635000 ;
      RECT 0.105000  0.085000 0.345000 0.885000 ;
      RECT 0.995000  0.085000 1.375000 0.465000 ;
      RECT 0.995000  0.635000 1.895000 0.840000 ;
      RECT 0.995000  0.840000 1.355000 1.330000 ;
      RECT 0.995000  2.185000 1.895000 2.635000 ;
      RECT 1.185000  1.330000 1.355000 1.785000 ;
      RECT 1.185000  1.785000 2.375000 2.005000 ;
      RECT 1.565000  0.255000 1.895000 0.635000 ;
      RECT 2.115000  0.465000 2.325000 0.635000 ;
      RECT 2.115000  0.635000 3.530000 0.825000 ;
      RECT 2.115000  2.005000 2.375000 2.465000 ;
      RECT 2.495000  0.085000 3.035000 0.465000 ;
      RECT 3.245000  1.650000 3.530000 2.635000 ;
      RECT 3.255000  0.495000 3.530000 0.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21a_2


MACRO sky130_fd_sc_hdll__o21a_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.760000 0.990000 4.115000 1.495000 ;
        RECT 3.760000 1.495000 5.880000 1.705000 ;
        RECT 5.410000 0.995000 5.880000 1.495000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.420000 0.995000 5.070000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.075000 3.485000 1.615000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.029000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.635000 1.865000 0.805000 ;
        RECT 0.090000 0.805000 0.350000 1.530000 ;
        RECT 0.090000 1.530000 2.155000 1.700000 ;
        RECT 0.645000 0.615000 1.865000 0.635000 ;
        RECT 1.015000 1.700000 1.205000 2.465000 ;
        RECT 1.975000 1.700000 2.155000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.415000  1.870000 0.795000 2.635000 ;
      RECT 0.520000  0.995000 2.565000 1.335000 ;
      RECT 1.055000  0.085000 1.385000 0.445000 ;
      RECT 1.375000  1.870000 1.755000 2.635000 ;
      RECT 2.015000  0.085000 2.345000 0.465000 ;
      RECT 2.315000  0.655000 3.385000 0.870000 ;
      RECT 2.315000  0.870000 2.565000 0.995000 ;
      RECT 2.325000  1.335000 2.565000 1.830000 ;
      RECT 2.325000  1.830000 3.195000 1.875000 ;
      RECT 2.325000  1.875000 4.875000 2.085000 ;
      RECT 2.335000  2.255000 2.735000 2.635000 ;
      RECT 2.585000  0.255000 3.885000 0.485000 ;
      RECT 2.955000  2.085000 4.875000 2.105000 ;
      RECT 2.955000  2.105000 3.195000 2.465000 ;
      RECT 3.515000  2.275000 3.845000 2.635000 ;
      RECT 3.555000  0.485000 3.885000 0.615000 ;
      RECT 3.555000  0.615000 5.835000 0.785000 ;
      RECT 4.055000  0.085000 4.395000 0.445000 ;
      RECT 4.495000  2.105000 4.875000 2.445000 ;
      RECT 4.975000  0.085000 5.355000 0.445000 ;
      RECT 5.455000  1.935000 5.865000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21a_4


MACRO sky130_fd_sc_hdll__o21a_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 1.075000 2.675000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.725000 1.075000 2.155000 1.275000 ;
        RECT 1.985000 1.275000 2.155000 2.390000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 1.075000 1.555000 1.305000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.472000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 1.030000 ;
        RECT 0.085000 1.030000 0.365000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.535000  1.860000 1.265000 2.635000 ;
      RECT 0.600000  0.715000 1.385000 0.905000 ;
      RECT 0.600000  0.905000 0.885000 1.475000 ;
      RECT 0.600000  1.475000 1.810000 1.690000 ;
      RECT 0.615000  0.085000 0.785000 0.545000 ;
      RECT 1.025000  0.255000 1.385000 0.715000 ;
      RECT 1.480000  1.690000 1.810000 2.465000 ;
      RECT 1.555000  0.555000 1.765000 0.715000 ;
      RECT 1.555000  0.715000 2.710000 0.905000 ;
      RECT 1.980000  0.085000 2.150000 0.545000 ;
      RECT 2.380000  0.255000 2.710000 0.715000 ;
      RECT 2.380000  1.915000 3.100000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21a_1


MACRO sky130_fd_sc_hdll__nor2_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  1.840000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.075000 1.395000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.435000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.495000 0.775000 1.665000 ;
        RECT 0.095000 1.665000 0.425000 2.450000 ;
        RECT 0.515000 0.255000 0.895000 0.895000 ;
        RECT 0.605000 0.895000 0.775000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.105000  0.085000 0.345000 0.895000 ;
      RECT 1.065000  0.085000 1.575000 0.895000 ;
      RECT 1.115000  1.495000 1.625000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2_1


MACRO sky130_fd_sc_hdll__nor2_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.280000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.075000 3.930000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.200000 1.075000 7.290000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.889000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 8.025000 0.905000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 2.415000 0.255000 2.795000 0.725000 ;
        RECT 3.355000 0.255000 3.735000 0.725000 ;
        RECT 4.295000 0.255000 4.675000 0.725000 ;
        RECT 4.385000 1.445000 8.025000 1.615000 ;
        RECT 4.385000 1.615000 4.635000 2.125000 ;
        RECT 5.235000 0.255000 5.615000 0.725000 ;
        RECT 5.325000 1.615000 5.575000 2.125000 ;
        RECT 6.175000 0.255000 6.555000 0.725000 ;
        RECT 6.265000 1.615000 6.515000 2.125000 ;
        RECT 7.115000 0.255000 7.495000 0.725000 ;
        RECT 7.205000 1.615000 7.455000 2.125000 ;
        RECT 7.460000 0.905000 8.025000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 4.165000 1.665000 ;
      RECT 0.090000  1.665000 0.405000 2.465000 ;
      RECT 0.625000  1.835000 0.875000 2.635000 ;
      RECT 1.095000  1.665000 1.345000 2.465000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 1.565000  1.835000 1.815000 2.635000 ;
      RECT 2.035000  1.665000 2.285000 2.465000 ;
      RECT 2.075000  0.085000 2.245000 0.555000 ;
      RECT 2.505000  1.835000 2.755000 2.635000 ;
      RECT 2.975000  1.665000 3.225000 2.465000 ;
      RECT 3.015000  0.085000 3.185000 0.555000 ;
      RECT 3.445000  1.835000 3.695000 2.635000 ;
      RECT 3.915000  1.665000 4.165000 2.295000 ;
      RECT 3.915000  2.295000 7.925000 2.465000 ;
      RECT 3.955000  0.085000 4.125000 0.555000 ;
      RECT 4.855000  1.785000 5.105000 2.295000 ;
      RECT 4.895000  0.085000 5.065000 0.555000 ;
      RECT 5.795000  1.785000 6.045000 2.295000 ;
      RECT 5.835000  0.085000 6.005000 0.555000 ;
      RECT 6.735000  1.785000 6.985000 2.295000 ;
      RECT 6.775000  0.085000 6.945000 0.555000 ;
      RECT 7.675000  1.785000 7.925000 2.295000 ;
      RECT 7.715000  0.085000 8.005000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2_8


MACRO sky130_fd_sc_hdll__nor2_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.860000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 1.075000 1.900000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.771000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 1.855000 0.735000 ;
        RECT 0.535000 0.735000 2.310000 0.905000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 1.475000 1.445000 2.310000 1.665000 ;
        RECT 1.475000 1.665000 1.855000 2.125000 ;
        RECT 2.095000 0.905000 2.310000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 1.305000 1.665000 ;
      RECT 0.090000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.915000 2.635000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 1.135000  1.665000 1.305000 2.295000 ;
      RECT 1.135000  2.295000 2.375000 2.465000 ;
      RECT 2.075000  1.835000 2.375000 2.295000 ;
      RECT 2.140000  0.085000 2.480000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2_2


MACRO sky130_fd_sc_hdll__nor2_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.950000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.320000 1.075000 3.835000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.477000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 4.490000 0.905000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 2.415000 0.255000 2.795000 0.725000 ;
        RECT 2.545000 1.445000 4.490000 1.745000 ;
        RECT 2.545000 1.745000 2.715000 2.125000 ;
        RECT 3.355000 0.255000 3.735000 0.725000 ;
        RECT 3.485000 1.745000 3.655000 2.125000 ;
        RECT 4.095000 0.905000 4.490000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 2.325000 1.665000 ;
      RECT 0.090000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.915000 2.635000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 1.135000  1.665000 1.305000 2.465000 ;
      RECT 1.475000  1.835000 1.775000 2.635000 ;
      RECT 1.945000  1.665000 2.325000 2.295000 ;
      RECT 1.945000  2.295000 4.290000 2.465000 ;
      RECT 2.075000  0.085000 2.245000 0.555000 ;
      RECT 2.885000  1.935000 3.265000 2.295000 ;
      RECT 3.015000  0.085000 3.185000 0.555000 ;
      RECT 3.825000  1.915000 4.290000 2.295000 ;
      RECT 3.955000  0.085000 4.240000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2_4


MACRO sky130_fd_sc_hdll__tap_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE WELLTAP ;
  SYMMETRY X Y R90 ;
  SIZE  0.460000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__tap_1


MACRO sky130_fd_sc_hdll__ebufn_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.765000 0.775000 1.675000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.516600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.765000 1.300000 1.275000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.445000 4.460000 1.625000 ;
        RECT 1.985000 1.625000 3.995000 1.765000 ;
        RECT 3.545000 0.635000 4.460000 0.855000 ;
        RECT 3.595000 1.765000 3.995000 2.125000 ;
        RECT 4.230000 0.855000 4.460000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.280000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.900000 0.595000 ;
      RECT 0.515000  1.845000 1.000000 2.635000 ;
      RECT 1.070000  0.255000 1.830000 0.595000 ;
      RECT 1.220000  1.445000 1.815000 1.765000 ;
      RECT 1.220000  1.765000 1.510000 2.465000 ;
      RECT 1.550000  0.595000 1.830000 1.025000 ;
      RECT 1.550000  1.025000 3.215000 1.275000 ;
      RECT 1.550000  1.275000 1.815000 1.445000 ;
      RECT 1.700000  1.935000 3.375000 2.105000 ;
      RECT 1.700000  2.105000 1.910000 2.465000 ;
      RECT 2.000000  0.255000 2.320000 0.655000 ;
      RECT 2.000000  0.655000 3.375000 0.855000 ;
      RECT 2.080000  2.275000 2.460000 2.635000 ;
      RECT 2.490000  0.085000 2.870000 0.485000 ;
      RECT 2.680000  2.105000 3.375000 2.295000 ;
      RECT 2.680000  2.295000 4.425000 2.465000 ;
      RECT 3.090000  0.275000 4.400000 0.465000 ;
      RECT 3.090000  0.465000 3.375000 0.655000 ;
      RECT 3.495000  1.025000 3.955000 1.275000 ;
      RECT 4.165000  1.795000 4.425000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.150000  1.060000 0.320000 1.230000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.680000  1.060000 3.850000 1.230000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
    LAYER met1 ;
      RECT 0.085000 1.030000 0.380000 1.120000 ;
      RECT 0.085000 1.120000 3.910000 1.260000 ;
      RECT 3.570000 1.030000 3.910000 1.120000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__ebufn_2


MACRO sky130_fd_sc_hdll__ebufn_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.04000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.430000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.631100 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 0.620000 1.405000 0.995000 ;
        RECT 1.020000 0.995000 1.530000 1.325000 ;
        RECT 1.020000 1.325000 1.405000 1.695000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  2.145000 1.445000 10.925000 1.725000 ;
        RECT  7.225000 0.615000 10.925000 0.855000 ;
        RECT 10.675000 0.855000 10.925000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 11.040000 0.085000 ;
      RECT 0.000000  2.635000 11.040000 2.805000 ;
      RECT 0.085000  0.085000  0.445000 0.825000 ;
      RECT 0.085000  1.785000  0.445000 2.635000 ;
      RECT 0.650000  0.280000  0.850000 1.615000 ;
      RECT 0.665000  1.615000  0.850000 2.465000 ;
      RECT 1.020000  0.085000  1.405000 0.445000 ;
      RECT 1.020000  1.865000  1.405000 2.635000 ;
      RECT 1.575000  0.255000  2.135000 0.825000 ;
      RECT 1.575000  1.495000  1.975000 2.465000 ;
      RECT 1.750000  0.825000  2.135000 1.025000 ;
      RECT 1.750000  1.025000  6.875000 1.275000 ;
      RECT 1.750000  1.275000  1.975000 1.495000 ;
      RECT 2.145000  1.895000 10.925000 2.065000 ;
      RECT 2.145000  2.065000  2.395000 2.465000 ;
      RECT 2.305000  0.255000  2.685000 0.655000 ;
      RECT 2.305000  0.655000  7.055000 0.855000 ;
      RECT 2.565000  2.235000  2.995000 2.635000 ;
      RECT 2.855000  0.085000  3.285000 0.485000 ;
      RECT 3.215000  2.065000  3.385000 2.465000 ;
      RECT 3.505000  0.275000  3.725000 0.655000 ;
      RECT 3.605000  2.235000  4.035000 2.635000 ;
      RECT 3.895000  0.085000  4.325000 0.485000 ;
      RECT 4.255000  2.065000  4.425000 2.465000 ;
      RECT 4.545000  0.255000  4.765000 0.655000 ;
      RECT 4.645000  2.235000  5.075000 2.635000 ;
      RECT 4.935000  0.085000  5.365000 0.485000 ;
      RECT 5.295000  2.065000  5.465000 2.465000 ;
      RECT 5.585000  0.275000  5.805000 0.655000 ;
      RECT 5.685000  2.235000  6.115000 2.635000 ;
      RECT 5.975000  0.085000  6.405000 0.485000 ;
      RECT 6.335000  2.065000 10.925000 2.465000 ;
      RECT 6.625000  0.255000 10.925000 0.445000 ;
      RECT 6.625000  0.445000  7.055000 0.655000 ;
      RECT 7.125000  1.025000 10.455000 1.275000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.655000  1.060000  0.825000 1.230000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.630000  1.060000  7.800000 1.230000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.545000 1.030000 0.885000 1.120000 ;
      RECT 0.545000 1.120000 7.860000 1.260000 ;
      RECT 7.520000 1.030000 7.860000 1.120000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__ebufn_8


MACRO sky130_fd_sc_hdll__ebufn_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.355000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.358200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 1.075000 1.290000 1.630000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.700500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.125000 1.495000 3.585000 2.465000 ;
        RECT 3.255000 0.255000 3.585000 0.825000 ;
        RECT 3.315000 0.825000 3.585000 1.495000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT -0.005000  2.635000 3.680000 2.805000 ;
      RECT  0.000000 -0.085000 3.680000 0.085000 ;
      RECT  0.085000  0.280000 0.345000 0.615000 ;
      RECT  0.085000  0.615000 1.235000 0.825000 ;
      RECT  0.085000  1.785000 0.790000 2.005000 ;
      RECT  0.085000  2.005000 0.345000 2.465000 ;
      RECT  0.515000  0.085000 0.895000 0.445000 ;
      RECT  0.515000  2.175000 0.890000 2.635000 ;
      RECT  0.525000  0.825000 0.790000 1.785000 ;
      RECT  1.065000  0.255000 2.175000 0.465000 ;
      RECT  1.065000  0.465000 1.235000 0.615000 ;
      RECT  1.115000  1.800000 1.905000 2.005000 ;
      RECT  1.115000  2.005000 1.370000 2.460000 ;
      RECT  1.460000  0.635000 1.790000 1.075000 ;
      RECT  1.460000  1.075000 2.745000 1.325000 ;
      RECT  1.460000  1.325000 1.905000 1.800000 ;
      RECT  1.540000  2.175000 1.900000 2.635000 ;
      RECT  1.960000  0.465000 2.175000 0.735000 ;
      RECT  1.960000  0.735000 3.085000 0.905000 ;
      RECT  2.345000  0.085000 3.085000 0.565000 ;
      RECT  2.915000  0.905000 3.085000 0.995000 ;
      RECT  2.915000  0.995000 3.145000 1.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__ebufn_1


MACRO sky130_fd_sc_hdll__ebufn_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 0.765000 0.830000 1.675000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.954300 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.765000 1.380000 1.425000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.445000 6.335000 1.725000 ;
        RECT 4.495000 0.615000 6.335000 0.855000 ;
        RECT 6.105000 0.855000 6.335000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  0.280000 0.345000 0.665000 ;
      RECT 0.085000  0.665000 0.320000 1.765000 ;
      RECT 0.085000  1.765000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.980000 0.595000 ;
      RECT 0.515000  1.845000 0.980000 2.635000 ;
      RECT 1.200000  0.255000 1.825000 0.595000 ;
      RECT 1.200000  1.595000 1.825000 1.765000 ;
      RECT 1.200000  1.765000 1.455000 2.465000 ;
      RECT 1.550000  0.595000 1.825000 1.025000 ;
      RECT 1.550000  1.025000 4.160000 1.275000 ;
      RECT 1.550000  1.275000 1.825000 1.595000 ;
      RECT 1.665000  1.935000 6.285000 2.105000 ;
      RECT 1.665000  2.105000 1.910000 2.465000 ;
      RECT 1.995000  0.255000 2.325000 0.655000 ;
      RECT 1.995000  0.655000 4.325000 0.855000 ;
      RECT 1.995000  1.895000 6.285000 1.935000 ;
      RECT 2.080000  2.275000 2.460000 2.635000 ;
      RECT 2.495000  0.085000 2.875000 0.485000 ;
      RECT 2.680000  2.105000 2.850000 2.465000 ;
      RECT 3.070000  2.275000 3.400000 2.635000 ;
      RECT 3.095000  0.275000 3.265000 0.655000 ;
      RECT 3.435000  0.085000 3.815000 0.485000 ;
      RECT 3.620000  2.105000 6.285000 2.465000 ;
      RECT 4.035000  0.255000 6.285000 0.445000 ;
      RECT 4.035000  0.445000 4.325000 0.655000 ;
      RECT 4.330000  1.025000 5.935000 1.275000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.150000  1.105000 0.320000 1.275000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.710000  1.105000 4.880000 1.275000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.085000 1.075000 0.380000 1.165000 ;
      RECT 0.085000 1.165000 4.940000 1.305000 ;
      RECT 4.650000 1.075000 4.940000 1.165000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__ebufn_4


MACRO sky130_fd_sc_hdll__o22ai_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.280000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 1.565000 1.275000 ;
        RECT 1.250000 1.275000 1.565000 1.445000 ;
        RECT 1.250000 1.445000 4.030000 1.615000 ;
        RECT 3.625000 1.075000 4.030000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.835000 1.075000 3.445000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.745000 0.995000 5.490000 1.445000 ;
        RECT 4.745000 1.445000 7.735000 1.615000 ;
        RECT 7.465000 0.995000 7.735000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.660000 1.075000 7.160000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.959500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 1.785000 4.370000 1.955000 ;
        RECT 1.955000 1.955000 2.295000 2.125000 ;
        RECT 2.985000 1.955000 3.235000 2.125000 ;
        RECT 4.200000 1.445000 4.575000 1.615000 ;
        RECT 4.200000 1.615000 4.370000 1.785000 ;
        RECT 4.355000 0.645000 8.170000 0.820000 ;
        RECT 4.355000 0.820000 4.575000 1.445000 ;
        RECT 5.855000 1.785000 8.170000 1.955000 ;
        RECT 5.855000 1.955000 6.105000 2.125000 ;
        RECT 6.795000 1.955000 7.045000 2.125000 ;
        RECT 7.905000 0.820000 8.170000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.125000  0.255000 0.455000 0.725000 ;
      RECT 0.125000  0.725000 1.395000 0.735000 ;
      RECT 0.125000  0.735000 4.185000 0.905000 ;
      RECT 0.165000  1.445000 0.415000 2.635000 ;
      RECT 0.635000  1.445000 0.885000 1.785000 ;
      RECT 0.635000  1.785000 1.785000 1.955000 ;
      RECT 0.635000  1.955000 0.885000 2.465000 ;
      RECT 0.675000  0.085000 0.845000 0.555000 ;
      RECT 1.015000  0.255000 1.395000 0.725000 ;
      RECT 1.105000  2.125000 1.355000 2.635000 ;
      RECT 1.575000  1.955000 1.785000 2.295000 ;
      RECT 1.575000  2.295000 3.745000 2.465000 ;
      RECT 1.615000  0.085000 1.785000 0.555000 ;
      RECT 1.955000  0.255000 2.335000 0.725000 ;
      RECT 1.955000  0.725000 3.275000 0.735000 ;
      RECT 2.515000  2.125000 2.765000 2.295000 ;
      RECT 2.555000  0.085000 2.725000 0.555000 ;
      RECT 2.895000  0.255000 3.275000 0.725000 ;
      RECT 3.455000  2.125000 3.745000 2.295000 ;
      RECT 3.495000  0.085000 3.665000 0.555000 ;
      RECT 3.835000  0.255000 8.045000 0.475000 ;
      RECT 3.835000  0.475000 4.185000 0.735000 ;
      RECT 3.965000  2.125000 4.185000 2.635000 ;
      RECT 4.355000  2.125000 4.710000 2.465000 ;
      RECT 4.540000  1.785000 5.635000 1.955000 ;
      RECT 4.540000  1.955000 4.710000 2.125000 ;
      RECT 4.925000  2.125000 5.165000 2.635000 ;
      RECT 5.385000  1.955000 5.635000 2.295000 ;
      RECT 5.385000  2.295000 7.515000 2.465000 ;
      RECT 6.325000  2.125000 6.575000 2.295000 ;
      RECT 7.265000  2.135000 7.515000 2.295000 ;
      RECT 7.735000  2.125000 8.015000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22ai_4


MACRO sky130_fd_sc_hdll__o22ai_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 1.075000 4.565000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.835000 1.075000 3.555000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.200000 1.075000 1.115000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.325000 1.075000 2.125000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.061000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.645000 2.645000 0.905000 ;
        RECT 1.565000 1.445000 3.315000 1.625000 ;
        RECT 1.565000 1.625000 1.815000 2.125000 ;
        RECT 2.405000 0.905000 2.645000 1.445000 ;
        RECT 3.065000 1.625000 3.315000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.090000  0.305000 2.985000 0.475000 ;
      RECT 0.090000  0.475000 0.365000 0.905000 ;
      RECT 0.150000  1.455000 1.345000 1.625000 ;
      RECT 0.150000  1.625000 0.405000 2.465000 ;
      RECT 0.625000  1.795000 0.875000 2.635000 ;
      RECT 1.095000  1.625000 1.345000 2.295000 ;
      RECT 1.095000  2.295000 2.285000 2.465000 ;
      RECT 2.035000  1.795000 2.285000 2.295000 ;
      RECT 2.595000  1.795000 2.845000 2.295000 ;
      RECT 2.595000  2.295000 3.785000 2.465000 ;
      RECT 2.815000  0.475000 2.985000 0.725000 ;
      RECT 2.815000  0.725000 4.765000 0.905000 ;
      RECT 3.155000  0.085000 3.325000 0.555000 ;
      RECT 3.495000  0.255000 3.825000 0.725000 ;
      RECT 3.535000  1.455000 4.730000 1.625000 ;
      RECT 3.535000  1.625000 3.785000 2.295000 ;
      RECT 4.005000  1.795000 4.255000 2.635000 ;
      RECT 4.045000  0.085000 4.215000 0.555000 ;
      RECT 4.385000  0.255000 4.765000 0.725000 ;
      RECT 4.475000  1.625000 4.730000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22ai_2


MACRO sky130_fd_sc_hdll__o22ai_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.150000 1.075000 2.660000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.075000 1.980000 1.245000 ;
        RECT 1.750000 1.245000 1.980000 1.445000 ;
        RECT 1.750000 1.445000 2.170000 1.615000 ;
        RECT 1.920000 1.615000 2.170000 2.405000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.665000 0.325000 1.990000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.995000 1.350000 1.665000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.816800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495000 0.645000 0.895000 0.825000 ;
        RECT 0.495000 0.825000 0.790000 1.835000 ;
        RECT 0.495000 1.835000 1.680000 2.045000 ;
        RECT 1.130000 2.045000 1.680000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.295000 1.620000 0.475000 ;
      RECT 0.135000  2.175000 0.345000 2.635000 ;
      RECT 1.290000  0.475000 1.620000 0.695000 ;
      RECT 1.290000  0.695000 2.660000 0.825000 ;
      RECT 1.460000  0.825000 2.660000 0.865000 ;
      RECT 1.890000  0.085000 2.060000 0.525000 ;
      RECT 2.270000  0.280000 2.660000 0.695000 ;
      RECT 2.340000  1.455000 2.660000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o22ai_1


MACRO sky130_fd_sc_hdll__o211a_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.165000 0.995000 2.675000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 0.995000 1.945000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.930000 0.995000 1.310000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.360000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.534000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945000 0.255000 3.325000 0.615000 ;
        RECT 2.945000 0.615000 4.035000 0.785000 ;
        RECT 3.085000 1.905000 4.035000 2.075000 ;
        RECT 3.085000 2.075000 3.275000 2.465000 ;
        RECT 3.765000 0.785000 4.035000 1.905000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  1.510000 3.025000 1.735000 ;
      RECT 0.090000  1.735000 1.820000 1.765000 ;
      RECT 0.090000  1.765000 0.355000 2.465000 ;
      RECT 0.095000  0.255000 0.430000 0.425000 ;
      RECT 0.095000  0.425000 0.760000 0.825000 ;
      RECT 0.525000  1.935000 0.905000 2.635000 ;
      RECT 0.530000  0.825000 0.760000 1.510000 ;
      RECT 0.930000  0.635000 2.375000 0.825000 ;
      RECT 1.125000  1.765000 1.820000 2.465000 ;
      RECT 1.535000  0.085000 1.870000 0.465000 ;
      RECT 2.375000  1.935000 2.855000 2.635000 ;
      RECT 2.540000  0.085000 2.775000 0.525000 ;
      RECT 2.855000  0.995000 3.565000 1.325000 ;
      RECT 2.855000  1.325000 3.025000 1.510000 ;
      RECT 3.445000  2.255000 3.825000 2.635000 ;
      RECT 3.545000  0.085000 3.875000 0.445000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211a_2


MACRO sky130_fd_sc_hdll__o211a_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.900000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.825000 1.035000 5.155000 1.495000 ;
        RECT 4.825000 1.495000 6.815000 1.685000 ;
        RECT 6.300000 1.035000 6.815000 1.495000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.340000 1.035000 6.115000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 0.995000 3.085000 1.445000 ;
        RECT 2.790000 1.445000 4.600000 1.685000 ;
        RECT 4.270000 1.035000 4.600000 1.445000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.255000 1.035000 4.090000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.016000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.635000 1.755000 0.805000 ;
        RECT 0.085000 0.805000 0.365000 1.435000 ;
        RECT 0.085000 1.435000 2.230000 1.700000 ;
        RECT 0.645000 0.255000 0.815000 0.615000 ;
        RECT 0.645000 0.615000 1.755000 0.635000 ;
        RECT 1.080000 1.700000 1.260000 2.465000 ;
        RECT 1.585000 0.255000 1.755000 0.615000 ;
        RECT 2.040000 1.700000 2.230000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.480000  1.870000 0.860000 2.635000 ;
      RECT 0.535000  1.065000 2.620000 1.265000 ;
      RECT 1.035000  0.085000 1.365000 0.445000 ;
      RECT 1.440000  1.870000 1.820000 2.635000 ;
      RECT 1.925000  0.085000 2.340000 0.465000 ;
      RECT 2.400000  0.635000 3.820000 0.815000 ;
      RECT 2.400000  0.815000 2.620000 1.065000 ;
      RECT 2.400000  1.265000 2.620000 1.855000 ;
      RECT 2.400000  1.855000 5.845000 2.025000 ;
      RECT 2.400000  2.200000 2.780000 2.635000 ;
      RECT 2.580000  0.255000 4.805000 0.465000 ;
      RECT 3.000000  2.025000 3.360000 2.465000 ;
      RECT 3.535000  2.195000 3.915000 2.635000 ;
      RECT 4.085000  2.025000 4.415000 2.465000 ;
      RECT 4.475000  0.465000 4.805000 0.695000 ;
      RECT 4.475000  0.695000 6.805000 0.865000 ;
      RECT 4.595000  2.195000 4.860000 2.635000 ;
      RECT 4.980000  0.085000 5.295000 0.525000 ;
      RECT 5.465000  0.255000 5.845000 0.695000 ;
      RECT 5.465000  2.025000 5.845000 2.465000 ;
      RECT 6.065000  0.085000 6.255000 0.525000 ;
      RECT 6.425000  0.255000 6.805000 0.695000 ;
      RECT 6.425000  1.915000 6.805000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211a_4


MACRO sky130_fd_sc_hdll__o211a_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.350000 1.075000 1.815000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.075000 2.370000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.540000 1.075000 3.080000 1.275000 ;
        RECT 2.815000 0.435000 3.080000 1.075000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.640000 1.075000 4.005000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 0.885000 ;
        RECT 0.085000 0.885000 0.260000 1.495000 ;
        RECT 0.085000 1.495000 0.425000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.430000  1.075000 1.175000 1.245000 ;
      RECT 0.645000  0.085000 0.895000 0.885000 ;
      RECT 0.645000  1.495000 0.815000 2.635000 ;
      RECT 1.005000  1.245000 1.175000 1.495000 ;
      RECT 1.005000  1.495000 3.800000 1.665000 ;
      RECT 1.085000  0.255000 1.415000 0.735000 ;
      RECT 1.085000  0.735000 2.410000 0.905000 ;
      RECT 1.085000  1.835000 1.335000 2.635000 ;
      RECT 1.635000  0.085000 1.860000 0.545000 ;
      RECT 2.030000  0.255000 2.410000 0.735000 ;
      RECT 2.085000  1.665000 2.465000 2.465000 ;
      RECT 2.760000  1.835000 3.090000 2.635000 ;
      RECT 3.250000  0.255000 3.800000 0.865000 ;
      RECT 3.250000  0.865000 3.470000 1.495000 ;
      RECT 3.470000  1.665000 3.800000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211a_1


MACRO sky130_fd_sc_hdll__and4_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.765000 0.330000 1.655000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.890000 0.420000 1.345000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 0.425000 1.780000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.730000 2.275000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 0.255000 2.955000 0.640000 ;
        RECT 2.785000 0.640000 4.455000 0.810000 ;
        RECT 2.785000 1.485000 4.455000 1.655000 ;
        RECT 2.785000 1.655000 3.035000 2.465000 ;
        RECT 3.725000 0.255000 3.895000 0.640000 ;
        RECT 3.725000 1.655000 4.455000 1.745000 ;
        RECT 3.725000 1.745000 3.895000 2.465000 ;
        RECT 4.200000 0.810000 4.455000 1.485000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.105000  1.835000 0.385000 2.635000 ;
      RECT 0.175000  0.255000 0.720000 0.585000 ;
      RECT 0.500000  0.585000 0.720000 1.495000 ;
      RECT 0.500000  1.495000 2.615000 1.665000 ;
      RECT 0.605000  1.665000 0.815000 2.465000 ;
      RECT 1.055000  1.935000 1.385000 2.635000 ;
      RECT 1.605000  1.665000 1.795000 2.465000 ;
      RECT 2.225000  0.085000 2.535000 0.550000 ;
      RECT 2.225000  1.855000 2.555000 2.635000 ;
      RECT 2.445000  1.075000 3.935000 1.305000 ;
      RECT 2.445000  1.305000 2.615000 1.495000 ;
      RECT 3.125000  0.085000 3.505000 0.470000 ;
      RECT 3.255000  1.835000 3.505000 2.635000 ;
      RECT 4.065000  0.085000 4.445000 0.470000 ;
      RECT 4.065000  1.915000 4.445000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4_4


MACRO sky130_fd_sc_hdll__and4_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.325000 2.075000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 0.360000 1.235000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.405000 0.355000 1.695000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 0.715000 2.165000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.752500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.695000 0.295000 3.085000 0.805000 ;
        RECT 2.695000 2.205000 3.085000 2.465000 ;
        RECT 2.825000 0.805000 3.085000 2.205000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  2.255000 0.425000 2.635000 ;
      RECT 0.170000  0.255000 0.685000 0.585000 ;
      RECT 0.495000  0.585000 0.685000 1.495000 ;
      RECT 0.495000  1.495000 2.535000 1.665000 ;
      RECT 0.605000  1.665000 0.855000 2.465000 ;
      RECT 1.035000  1.915000 1.365000 2.635000 ;
      RECT 1.560000  1.665000 1.810000 2.465000 ;
      RECT 2.005000  1.835000 2.375000 2.635000 ;
      RECT 2.065000  0.085000 2.335000 0.545000 ;
      RECT 2.335000  0.995000 2.535000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4_1


MACRO sky130_fd_sc_hdll__and4_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.755000 0.330000 2.075000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 0.420000 1.235000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.405000 0.415000 1.705000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 0.740000 2.155000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.629500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.625000 0.295000 3.075000 0.805000 ;
        RECT 2.625000 1.835000 3.075000 2.465000 ;
        RECT 2.835000 0.805000 3.075000 1.835000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  2.255000 0.425000 2.635000 ;
      RECT 0.175000  0.255000 0.670000 0.585000 ;
      RECT 0.500000  0.585000 0.670000 1.495000 ;
      RECT 0.500000  1.495000 2.665000 1.665000 ;
      RECT 0.645000  1.665000 0.815000 2.465000 ;
      RECT 1.035000  1.915000 1.365000 2.635000 ;
      RECT 1.570000  1.665000 1.820000 2.465000 ;
      RECT 2.165000  1.835000 2.415000 2.635000 ;
      RECT 2.285000  0.085000 2.455000 0.550000 ;
      RECT 2.495000  0.995000 2.665000 1.495000 ;
      RECT 3.245000  0.085000 3.575000 0.810000 ;
      RECT 3.245000  1.835000 3.565000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4_2


MACRO sky130_fd_sc_hdll__bufinv_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.900000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.505000 1.275000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.915000 0.260000 3.295000 0.735000 ;
        RECT 2.915000 0.735000 6.805000 0.905000 ;
        RECT 2.915000 1.445000 6.805000 1.615000 ;
        RECT 2.915000 1.615000 3.295000 2.465000 ;
        RECT 3.855000 0.260000 4.235000 0.735000 ;
        RECT 3.855000 1.615000 4.235000 2.465000 ;
        RECT 4.795000 0.260000 5.175000 0.735000 ;
        RECT 4.795000 1.615000 5.175000 2.465000 ;
        RECT 5.735000 0.260000 6.115000 0.735000 ;
        RECT 5.735000 1.615000 6.115000 2.465000 ;
        RECT 6.415000 0.905000 6.805000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.175000  0.085000 0.345000 0.905000 ;
      RECT 0.175000  1.445000 0.345000 2.635000 ;
      RECT 0.515000  0.260000 0.895000 0.905000 ;
      RECT 0.515000  1.545000 0.895000 2.465000 ;
      RECT 0.725000  0.905000 0.895000 1.075000 ;
      RECT 0.725000  1.075000 2.355000 1.275000 ;
      RECT 0.725000  1.275000 0.895000 1.545000 ;
      RECT 1.085000  0.260000 1.415000 0.735000 ;
      RECT 1.085000  0.735000 2.745000 0.905000 ;
      RECT 1.085000  1.445000 2.745000 1.615000 ;
      RECT 1.085000  1.615000 1.415000 2.465000 ;
      RECT 1.635000  0.085000 1.805000 0.565000 ;
      RECT 1.635000  1.785000 1.805000 2.635000 ;
      RECT 1.975000  0.260000 2.355000 0.735000 ;
      RECT 1.975000  1.615000 2.355000 2.465000 ;
      RECT 2.575000  0.085000 2.745000 0.565000 ;
      RECT 2.575000  0.905000 2.745000 1.075000 ;
      RECT 2.575000  1.075000 6.245000 1.275000 ;
      RECT 2.575000  1.275000 2.745000 1.445000 ;
      RECT 2.575000  1.785000 2.745000 2.635000 ;
      RECT 3.515000  0.085000 3.685000 0.565000 ;
      RECT 3.515000  1.835000 3.685000 2.635000 ;
      RECT 4.455000  0.085000 4.625000 0.565000 ;
      RECT 4.455000  1.835000 4.625000 2.635000 ;
      RECT 5.395000  0.085000 5.565000 0.565000 ;
      RECT 5.395000  1.835000 5.565000 2.635000 ;
      RECT 6.335000  0.085000 6.505000 0.565000 ;
      RECT 6.335000  1.835000 6.505000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__bufinv_8


MACRO sky130_fd_sc_hdll__bufinv_16
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  12.42000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.832500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.365000 1.275000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.016500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  4.745000 0.255000  5.045000 0.260000 ;
        RECT  4.745000 0.260000  5.125000 0.735000 ;
        RECT  4.745000 0.735000 12.205000 0.905000 ;
        RECT  4.745000 1.445000 12.205000 1.615000 ;
        RECT  4.745000 1.615000  5.125000 2.465000 ;
        RECT  5.685000 0.260000  6.065000 0.735000 ;
        RECT  5.685000 1.615000  6.065000 2.465000 ;
        RECT  5.815000 0.255000  5.985000 0.260000 ;
        RECT  6.625000 0.260000  7.005000 0.735000 ;
        RECT  6.625000 1.615000  7.005000 2.465000 ;
        RECT  6.755000 0.255000  6.925000 0.260000 ;
        RECT  7.565000 0.260000  7.945000 0.735000 ;
        RECT  7.565000 1.615000  7.945000 2.465000 ;
        RECT  8.505000 0.260000  8.885000 0.735000 ;
        RECT  8.505000 1.615000  8.885000 2.465000 ;
        RECT  9.445000 0.260000  9.825000 0.735000 ;
        RECT  9.445000 1.615000  9.825000 2.465000 ;
        RECT 10.385000 0.260000 10.765000 0.735000 ;
        RECT 10.385000 1.615000 10.765000 2.465000 ;
        RECT 11.325000 0.260000 11.705000 0.735000 ;
        RECT 11.325000 1.615000 11.705000 2.465000 ;
        RECT 11.930000 0.905000 12.205000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.095000  0.260000  0.425000 0.735000 ;
      RECT  0.095000  0.735000  1.755000 0.905000 ;
      RECT  0.095000  1.445000  1.755000 1.615000 ;
      RECT  0.095000  1.615000  0.425000 2.465000 ;
      RECT  0.645000  0.085000  0.815000 0.565000 ;
      RECT  0.645000  1.785000  0.815000 2.635000 ;
      RECT  0.985000  0.260000  1.365000 0.735000 ;
      RECT  0.985000  1.615000  1.365000 2.465000 ;
      RECT  1.585000  0.085000  1.755000 0.565000 ;
      RECT  1.585000  0.905000  1.755000 1.075000 ;
      RECT  1.585000  1.075000  4.145000 1.275000 ;
      RECT  1.585000  1.275000  1.755000 1.445000 ;
      RECT  1.585000  1.785000  1.755000 2.635000 ;
      RECT  1.925000  0.260000  2.305000 0.735000 ;
      RECT  1.925000  0.735000  4.575000 0.905000 ;
      RECT  1.925000  1.445000  4.575000 1.615000 ;
      RECT  1.925000  1.615000  2.305000 2.465000 ;
      RECT  2.525000  0.085000  2.695000 0.565000 ;
      RECT  2.525000  1.835000  2.695000 2.635000 ;
      RECT  2.865000  0.260000  3.245000 0.735000 ;
      RECT  2.865000  1.615000  3.245000 2.465000 ;
      RECT  3.465000  0.085000  3.635000 0.565000 ;
      RECT  3.465000  1.835000  3.635000 2.635000 ;
      RECT  3.805000  0.260000  4.185000 0.735000 ;
      RECT  3.805000  1.615000  4.185000 2.465000 ;
      RECT  4.400000  0.905000  4.575000 1.075000 ;
      RECT  4.400000  1.075000 11.710000 1.275000 ;
      RECT  4.400000  1.275000  4.575000 1.445000 ;
      RECT  4.405000  0.085000  4.575000 0.565000 ;
      RECT  4.405000  1.835000  4.575000 2.635000 ;
      RECT  5.345000  0.085000  5.515000 0.565000 ;
      RECT  5.345000  1.835000  5.515000 2.635000 ;
      RECT  6.285000  0.085000  6.455000 0.565000 ;
      RECT  6.285000  1.835000  6.455000 2.635000 ;
      RECT  7.225000  0.085000  7.395000 0.565000 ;
      RECT  7.225000  1.835000  7.395000 2.635000 ;
      RECT  8.165000  0.085000  8.335000 0.565000 ;
      RECT  8.165000  1.835000  8.335000 2.635000 ;
      RECT  9.105000  0.085000  9.275000 0.565000 ;
      RECT  9.105000  1.835000  9.275000 2.635000 ;
      RECT 10.045000  0.085000 10.215000 0.565000 ;
      RECT 10.045000  1.835000 10.215000 2.635000 ;
      RECT 10.985000  0.085000 11.155000 0.565000 ;
      RECT 10.985000  1.835000 11.155000 2.635000 ;
      RECT 11.925000  0.085000 12.095000 0.565000 ;
      RECT 11.925000  1.835000 12.095000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__bufinv_16


MACRO sky130_fd_sc_hdll__dlygate4sd2_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.605000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.464000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.780000 0.255000 3.110000 0.825000 ;
        RECT 2.780000 1.495000 3.110000 2.465000 ;
        RECT 2.860000 0.825000 3.110000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.785000 0.945000 2.005000 ;
      RECT 0.085000  2.005000 0.380000 2.465000 ;
      RECT 0.095000  0.255000 0.380000 0.715000 ;
      RECT 0.095000  0.715000 0.945000 0.885000 ;
      RECT 0.600000  0.085000 0.815000 0.545000 ;
      RECT 0.600000  2.175000 0.815000 2.635000 ;
      RECT 0.775000  0.885000 0.945000 0.995000 ;
      RECT 0.775000  0.995000 1.080000 1.325000 ;
      RECT 0.775000  1.325000 0.945000 1.785000 ;
      RECT 0.985000  0.255000 1.420000 0.545000 ;
      RECT 0.985000  2.175000 1.420000 2.465000 ;
      RECT 1.250000  0.545000 1.420000 1.075000 ;
      RECT 1.250000  1.075000 2.095000 1.275000 ;
      RECT 1.250000  1.275000 1.420000 2.175000 ;
      RECT 1.615000  0.510000 1.840000 0.735000 ;
      RECT 1.615000  0.735000 2.610000 0.905000 ;
      RECT 1.615000  1.575000 2.610000 1.745000 ;
      RECT 1.615000  1.745000 1.840000 2.080000 ;
      RECT 2.145000  0.085000 2.555000 0.565000 ;
      RECT 2.145000  1.915000 2.515000 2.635000 ;
      RECT 2.400000  0.905000 2.610000 0.995000 ;
      RECT 2.400000  0.995000 2.690000 1.325000 ;
      RECT 2.400000  1.325000 2.610000 1.575000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlygate4sd2_1


MACRO sky130_fd_sc_hdll__sdfrtn_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  12.88000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK_N
  PIN D
    ANTENNAGATEAREA  0.160200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.120000 1.355000 3.655000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.513200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.420000 0.265000 12.785000 2.325000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.145000 0.735000  7.900000 0.780000 ;
        RECT  7.145000 0.780000 11.405000 0.920000 ;
        RECT  7.145000 0.920000  7.900000 0.965000 ;
        RECT 11.115000 0.735000 11.405000 0.780000 ;
        RECT 11.115000 0.920000 11.405000 0.965000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.172800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.610000 0.710000 4.955000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.467400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.070000 1.990000 1.335000 ;
        RECT 1.585000 1.335000 2.220000 1.745000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.880000 0.085000 ;
      RECT  0.000000  2.635000 12.880000 2.805000 ;
      RECT  0.090000  1.795000  0.915000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.885000 0.805000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.530000  2.135000  0.910000 2.635000 ;
      RECT  0.710000  0.805000  0.885000 0.995000 ;
      RECT  0.710000  0.995000  1.025000 1.325000 ;
      RECT  0.710000  1.325000  0.915000 1.795000 ;
      RECT  1.115000  0.345000  1.365000 0.675000 ;
      RECT  1.135000  1.730000  1.365000 2.465000 ;
      RECT  1.195000  0.675000  1.365000 1.730000 ;
      RECT  1.695000  0.395000  1.865000 0.730000 ;
      RECT  1.695000  0.730000  2.435000 0.900000 ;
      RECT  2.035000  0.085000  2.415000 0.560000 ;
      RECT  2.110000  1.915000  2.730000 2.085000 ;
      RECT  2.110000  2.085000  2.380000 2.400000 ;
      RECT  2.265000  0.900000  2.435000 0.995000 ;
      RECT  2.265000  0.995000  3.445000 1.165000 ;
      RECT  2.475000  1.165000  3.445000 1.185000 ;
      RECT  2.475000  1.185000  2.730000 1.915000 ;
      RECT  2.600000  2.255000  2.930000 2.635000 ;
      RECT  2.655000  0.085000  3.035000 0.825000 ;
      RECT  3.275000  0.255000  4.435000 0.425000 ;
      RECT  3.275000  0.425000  3.445000 0.995000 ;
      RECT  3.665000  0.675000  4.045000 1.075000 ;
      RECT  3.870000  1.075000  4.045000 1.935000 ;
      RECT  3.870000  1.935000  5.650000 2.105000 ;
      RECT  3.870000  2.105000  4.040000 2.465000 ;
      RECT  4.265000  0.425000  4.435000 1.685000 ;
      RECT  4.855000  2.275000  5.205000 2.635000 ;
      RECT  5.005000  0.085000  5.350000 0.540000 ;
      RECT  5.140000  0.715000  5.720000 0.895000 ;
      RECT  5.140000  0.895000  5.310000 1.935000 ;
      RECT  5.480000  1.065000  5.650000 1.395000 ;
      RECT  5.480000  2.105000  5.650000 2.185000 ;
      RECT  5.480000  2.185000  5.850000 2.435000 ;
      RECT  5.550000  0.335000  5.890000 0.505000 ;
      RECT  5.550000  0.505000  5.720000 0.715000 ;
      RECT  5.820000  1.575000  6.120000 1.955000 ;
      RECT  5.900000  0.705000  6.650000 1.035000 ;
      RECT  5.900000  1.035000  6.120000 1.575000 ;
      RECT  6.095000  2.135000  6.460000 2.465000 ;
      RECT  6.110000  0.305000  7.010000 0.475000 ;
      RECT  6.290000  1.215000  8.150000 1.385000 ;
      RECT  6.290000  1.385000  6.460000 2.135000 ;
      RECT  6.680000  1.935000  7.940000 2.105000 ;
      RECT  6.680000  2.105000  6.850000 2.375000 ;
      RECT  6.840000  0.475000  7.010000 1.215000 ;
      RECT  6.960000  1.595000  8.540000 1.765000 ;
      RECT  7.135000  2.355000  7.465000 2.635000 ;
      RECT  7.230000  0.765000  7.810000 1.045000 ;
      RECT  7.690000  0.085000  8.020000 0.545000 ;
      RECT  7.770000  2.105000  7.940000 2.375000 ;
      RECT  7.980000  1.005000  8.150000 1.215000 ;
      RECT  8.150000  2.175000  8.570000 2.635000 ;
      RECT  8.230000  0.275000  8.610000 0.445000 ;
      RECT  8.230000  0.445000  8.540000 0.835000 ;
      RECT  8.230000  1.765000  8.540000 1.835000 ;
      RECT  8.230000  1.835000  8.985000 2.005000 ;
      RECT  8.370000  0.835000  8.540000 1.595000 ;
      RECT  8.710000  0.705000  8.970000 1.495000 ;
      RECT  8.710000  1.495000  9.445000 1.660000 ;
      RECT  8.710000  1.660000  9.845000 1.665000 ;
      RECT  8.780000  0.255000  9.890000 0.535000 ;
      RECT  8.815000  2.005000  8.985000 2.465000 ;
      RECT  9.185000  1.665000  9.845000 1.955000 ;
      RECT  9.195000  2.125000 10.215000 2.465000 ;
      RECT  9.235000  0.920000  9.405000 1.325000 ;
      RECT  9.670000  0.535000  9.890000 1.315000 ;
      RECT  9.670000  1.315000 10.285000 1.485000 ;
      RECT 10.040000  1.485000 10.285000 1.575000 ;
      RECT 10.040000  1.575000 11.370000 1.745000 ;
      RECT 10.040000  1.745000 10.215000 2.125000 ;
      RECT 10.110000  0.085000 10.330000 0.525000 ;
      RECT 10.150000  0.695000 10.730000 0.865000 ;
      RECT 10.150000  0.865000 10.370000 1.145000 ;
      RECT 10.415000  2.195000 10.665000 2.635000 ;
      RECT 10.560000  0.295000 11.735000 0.465000 ;
      RECT 10.560000  0.465000 10.730000 0.695000 ;
      RECT 10.600000  1.065000 11.370000 1.275000 ;
      RECT 10.910000  1.915000 11.730000 2.085000 ;
      RECT 10.910000  2.085000 11.080000 2.375000 ;
      RECT 11.065000  0.635000 11.370000 1.065000 ;
      RECT 11.255000  2.255000 11.635000 2.635000 ;
      RECT 11.560000  0.465000 11.735000 0.995000 ;
      RECT 11.560000  0.995000 12.205000 1.325000 ;
      RECT 11.560000  1.325000 11.730000 1.915000 ;
      RECT 11.905000  0.085000 12.190000 0.710000 ;
      RECT 11.905000  1.495000 12.190000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.725000  1.785000  0.895000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.195000  1.105000  1.365000 1.275000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.480000  1.105000  5.650000 1.275000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.950000  1.785000  6.120000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.255000  0.765000  7.425000 0.935000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.615000  0.765000  7.785000 0.935000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.235000  1.105000  9.405000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.565000  1.785000  9.735000 1.955000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.175000  0.765000 11.345000 0.935000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
    LAYER met1 ;
      RECT 0.660000 1.755000 0.960000 1.800000 ;
      RECT 0.660000 1.800000 9.795000 1.940000 ;
      RECT 0.660000 1.940000 0.960000 1.985000 ;
      RECT 1.135000 1.075000 1.425000 1.120000 ;
      RECT 1.135000 1.120000 9.465000 1.260000 ;
      RECT 1.135000 1.260000 1.425000 1.305000 ;
      RECT 5.420000 1.075000 5.710000 1.120000 ;
      RECT 5.420000 1.260000 5.710000 1.305000 ;
      RECT 5.890000 1.755000 6.180000 1.800000 ;
      RECT 5.890000 1.940000 6.180000 1.985000 ;
      RECT 9.155000 1.075000 9.465000 1.120000 ;
      RECT 9.155000 1.260000 9.465000 1.305000 ;
      RECT 9.500000 1.755000 9.795000 1.800000 ;
      RECT 9.500000 1.940000 9.795000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrtn_1


MACRO sky130_fd_sc_hdll__sdfrbp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  14.72000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.160200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.120000 1.355000 3.655000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.860000 0.265000 13.260000 1.695000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.494700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.770000 1.535000 14.205000 2.080000 ;
        RECT 13.780000 0.310000 14.205000 0.825000 ;
        RECT 14.035000 0.825000 14.205000 1.535000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.145000 0.735000  7.900000 0.780000 ;
        RECT  7.145000 0.780000 11.405000 0.920000 ;
        RECT  7.145000 0.920000  7.900000 0.965000 ;
        RECT 11.115000 0.735000 11.405000 0.780000 ;
        RECT 11.115000 0.920000 11.405000 0.965000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.172800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.610000 0.710000 4.955000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.467400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.070000 1.990000 1.335000 ;
        RECT 1.585000 1.335000 2.220000 1.745000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.720000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.720000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.720000 0.085000 ;
      RECT  0.000000  2.635000 14.720000 2.805000 ;
      RECT  0.090000  1.795000  0.915000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.885000 0.805000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.530000  2.135000  0.910000 2.635000 ;
      RECT  0.710000  0.805000  0.885000 0.995000 ;
      RECT  0.710000  0.995000  1.025000 1.325000 ;
      RECT  0.710000  1.325000  0.915000 1.795000 ;
      RECT  1.115000  0.345000  1.365000 0.675000 ;
      RECT  1.135000  1.730000  1.365000 2.465000 ;
      RECT  1.195000  0.675000  1.365000 1.730000 ;
      RECT  1.695000  0.395000  1.865000 0.730000 ;
      RECT  1.695000  0.730000  2.435000 0.900000 ;
      RECT  2.035000  0.085000  2.415000 0.560000 ;
      RECT  2.110000  1.915000  2.730000 2.085000 ;
      RECT  2.110000  2.085000  2.380000 2.400000 ;
      RECT  2.265000  0.900000  2.435000 0.995000 ;
      RECT  2.265000  0.995000  3.445000 1.165000 ;
      RECT  2.475000  1.165000  3.445000 1.185000 ;
      RECT  2.475000  1.185000  2.730000 1.915000 ;
      RECT  2.600000  2.255000  2.930000 2.635000 ;
      RECT  2.655000  0.085000  3.035000 0.825000 ;
      RECT  3.275000  0.255000  4.435000 0.425000 ;
      RECT  3.275000  0.425000  3.445000 0.995000 ;
      RECT  3.665000  0.675000  4.045000 1.075000 ;
      RECT  3.870000  1.075000  4.045000 1.935000 ;
      RECT  3.870000  1.935000  5.650000 2.105000 ;
      RECT  3.870000  2.105000  4.040000 2.465000 ;
      RECT  4.265000  0.425000  4.435000 1.685000 ;
      RECT  4.855000  2.275000  5.205000 2.635000 ;
      RECT  5.005000  0.085000  5.350000 0.540000 ;
      RECT  5.140000  0.715000  5.720000 0.895000 ;
      RECT  5.140000  0.895000  5.310000 1.935000 ;
      RECT  5.480000  1.065000  5.650000 1.395000 ;
      RECT  5.480000  2.105000  5.650000 2.185000 ;
      RECT  5.480000  2.185000  5.850000 2.435000 ;
      RECT  5.550000  0.335000  5.890000 0.505000 ;
      RECT  5.550000  0.505000  5.720000 0.715000 ;
      RECT  5.820000  1.575000  6.120000 1.955000 ;
      RECT  5.900000  0.705000  6.650000 1.035000 ;
      RECT  5.900000  1.035000  6.120000 1.575000 ;
      RECT  6.095000  2.135000  6.460000 2.465000 ;
      RECT  6.110000  0.305000  7.010000 0.475000 ;
      RECT  6.290000  1.215000  8.150000 1.385000 ;
      RECT  6.290000  1.385000  6.460000 2.135000 ;
      RECT  6.680000  1.935000  7.940000 2.105000 ;
      RECT  6.680000  2.105000  6.850000 2.375000 ;
      RECT  6.840000  0.475000  7.010000 1.215000 ;
      RECT  6.960000  1.595000  8.540000 1.765000 ;
      RECT  7.135000  2.355000  7.465000 2.635000 ;
      RECT  7.230000  0.765000  7.810000 1.045000 ;
      RECT  7.690000  0.085000  8.020000 0.545000 ;
      RECT  7.770000  2.105000  7.940000 2.375000 ;
      RECT  7.980000  1.005000  8.150000 1.215000 ;
      RECT  8.150000  2.175000  8.570000 2.635000 ;
      RECT  8.230000  0.275000  8.610000 0.445000 ;
      RECT  8.230000  0.445000  8.540000 0.835000 ;
      RECT  8.230000  1.765000  8.540000 1.835000 ;
      RECT  8.230000  1.835000  8.985000 2.005000 ;
      RECT  8.370000  0.835000  8.540000 1.595000 ;
      RECT  8.710000  0.705000  8.970000 1.495000 ;
      RECT  8.710000  1.495000  9.445000 1.660000 ;
      RECT  8.710000  1.660000  9.845000 1.665000 ;
      RECT  8.780000  0.255000  9.890000 0.535000 ;
      RECT  8.815000  2.005000  8.985000 2.465000 ;
      RECT  9.185000  1.665000  9.845000 1.955000 ;
      RECT  9.195000  2.125000 10.215000 2.465000 ;
      RECT  9.235000  0.920000  9.405000 1.325000 ;
      RECT  9.670000  0.535000  9.890000 1.315000 ;
      RECT  9.670000  1.315000 10.285000 1.485000 ;
      RECT 10.040000  1.485000 10.285000 1.575000 ;
      RECT 10.040000  1.575000 11.370000 1.745000 ;
      RECT 10.040000  1.745000 10.215000 2.125000 ;
      RECT 10.110000  0.085000 10.330000 0.525000 ;
      RECT 10.150000  0.695000 10.730000 0.865000 ;
      RECT 10.150000  0.865000 10.370000 1.145000 ;
      RECT 10.415000  2.195000 10.665000 2.635000 ;
      RECT 10.560000  0.295000 11.730000 0.465000 ;
      RECT 10.560000  0.465000 10.730000 0.695000 ;
      RECT 10.600000  1.065000 11.370000 1.275000 ;
      RECT 10.910000  1.915000 11.730000 2.085000 ;
      RECT 10.910000  2.085000 11.080000 2.375000 ;
      RECT 11.065000  0.635000 11.370000 1.065000 ;
      RECT 11.255000  2.255000 11.635000 2.635000 ;
      RECT 11.560000  0.465000 11.730000 0.995000 ;
      RECT 11.560000  0.995000 12.205000 1.325000 ;
      RECT 11.560000  1.325000 11.730000 1.915000 ;
      RECT 11.900000  0.345000 12.070000 0.655000 ;
      RECT 11.900000  0.655000 12.640000 0.825000 ;
      RECT 11.900000  1.795000 12.640000 1.865000 ;
      RECT 11.900000  1.865000 13.600000 2.035000 ;
      RECT 11.900000  2.035000 12.075000 2.465000 ;
      RECT 12.255000  2.205000 12.715000 2.635000 ;
      RECT 12.325000  0.085000 12.655000 0.485000 ;
      RECT 12.465000  0.825000 12.640000 1.795000 ;
      RECT 13.270000  2.255000 13.725000 2.635000 ;
      RECT 13.430000  0.995000 13.865000 1.325000 ;
      RECT 13.430000  1.325000 13.600000 1.865000 ;
      RECT 13.440000  0.085000 13.610000 0.825000 ;
      RECT 14.375000  0.085000 14.545000 0.930000 ;
      RECT 14.375000  1.495000 14.625000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.855000  1.105000  1.025000 1.275000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.135000  1.785000  1.305000 1.955000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.480000  1.105000  5.650000 1.275000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.950000  1.785000  6.120000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.255000  0.765000  7.425000 0.935000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.615000  0.765000  7.785000 0.935000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.235000  1.105000  9.405000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.565000  1.785000  9.735000 1.955000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.175000  0.765000 11.345000 0.935000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
    LAYER met1 ;
      RECT 0.795000 1.075000 1.085000 1.120000 ;
      RECT 0.795000 1.120000 9.465000 1.260000 ;
      RECT 0.795000 1.260000 1.085000 1.305000 ;
      RECT 1.070000 1.755000 1.370000 1.800000 ;
      RECT 1.070000 1.800000 9.795000 1.940000 ;
      RECT 1.070000 1.940000 1.370000 1.985000 ;
      RECT 5.420000 1.075000 5.710000 1.120000 ;
      RECT 5.420000 1.260000 5.710000 1.305000 ;
      RECT 5.890000 1.755000 6.180000 1.800000 ;
      RECT 5.890000 1.940000 6.180000 1.985000 ;
      RECT 9.155000 1.075000 9.465000 1.120000 ;
      RECT 9.155000 1.260000 9.465000 1.305000 ;
      RECT 9.500000 1.755000 9.795000 1.800000 ;
      RECT 9.500000 1.940000 9.795000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrbp_2


MACRO sky130_fd_sc_hdll__sdfrbp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  14.26000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.160200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.120000 1.355000 3.655000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.513200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.420000 0.265000 12.770000 2.395000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.374700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.885000 0.255000 14.165000 0.870000 ;
        RECT 13.885000 1.475000 14.165000 2.465000 ;
        RECT 13.935000 0.870000 14.165000 1.475000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.145000 0.735000  7.900000 0.780000 ;
        RECT  7.145000 0.780000 11.405000 0.920000 ;
        RECT  7.145000 0.920000  7.900000 0.965000 ;
        RECT 11.115000 0.735000 11.405000 0.780000 ;
        RECT 11.115000 0.920000 11.405000 0.965000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.172800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.610000 0.710000 4.955000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.467400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.070000 1.990000 1.335000 ;
        RECT 1.585000 1.335000 2.220000 1.745000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.090000  1.795000  0.915000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.885000 0.805000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.530000  2.135000  0.910000 2.635000 ;
      RECT  0.710000  0.805000  0.885000 0.995000 ;
      RECT  0.710000  0.995000  1.025000 1.325000 ;
      RECT  0.710000  1.325000  0.915000 1.795000 ;
      RECT  1.115000  0.345000  1.365000 0.675000 ;
      RECT  1.135000  1.730000  1.365000 2.465000 ;
      RECT  1.195000  0.675000  1.365000 1.730000 ;
      RECT  1.695000  0.395000  1.865000 0.730000 ;
      RECT  1.695000  0.730000  2.435000 0.900000 ;
      RECT  2.035000  0.085000  2.415000 0.560000 ;
      RECT  2.110000  1.915000  2.730000 2.085000 ;
      RECT  2.110000  2.085000  2.380000 2.400000 ;
      RECT  2.265000  0.900000  2.435000 0.995000 ;
      RECT  2.265000  0.995000  3.445000 1.165000 ;
      RECT  2.475000  1.165000  3.445000 1.185000 ;
      RECT  2.475000  1.185000  2.730000 1.915000 ;
      RECT  2.600000  2.255000  2.930000 2.635000 ;
      RECT  2.655000  0.085000  3.035000 0.825000 ;
      RECT  3.275000  0.255000  4.435000 0.425000 ;
      RECT  3.275000  0.425000  3.445000 0.995000 ;
      RECT  3.665000  0.675000  4.045000 1.075000 ;
      RECT  3.870000  1.075000  4.045000 1.935000 ;
      RECT  3.870000  1.935000  5.650000 2.105000 ;
      RECT  3.870000  2.105000  4.040000 2.465000 ;
      RECT  4.265000  0.425000  4.435000 1.685000 ;
      RECT  4.855000  2.275000  5.205000 2.635000 ;
      RECT  5.005000  0.085000  5.350000 0.540000 ;
      RECT  5.140000  0.715000  5.720000 0.895000 ;
      RECT  5.140000  0.895000  5.310000 1.935000 ;
      RECT  5.480000  1.065000  5.650000 1.395000 ;
      RECT  5.480000  2.105000  5.650000 2.185000 ;
      RECT  5.480000  2.185000  5.850000 2.435000 ;
      RECT  5.550000  0.335000  5.890000 0.505000 ;
      RECT  5.550000  0.505000  5.720000 0.715000 ;
      RECT  5.820000  1.575000  6.120000 1.955000 ;
      RECT  5.900000  0.705000  6.650000 1.035000 ;
      RECT  5.900000  1.035000  6.120000 1.575000 ;
      RECT  6.095000  2.135000  6.460000 2.465000 ;
      RECT  6.110000  0.305000  7.010000 0.475000 ;
      RECT  6.290000  1.215000  8.150000 1.385000 ;
      RECT  6.290000  1.385000  6.460000 2.135000 ;
      RECT  6.680000  1.935000  7.940000 2.105000 ;
      RECT  6.680000  2.105000  6.850000 2.375000 ;
      RECT  6.840000  0.475000  7.010000 1.215000 ;
      RECT  6.960000  1.595000  8.540000 1.765000 ;
      RECT  7.135000  2.355000  7.465000 2.635000 ;
      RECT  7.230000  0.765000  7.810000 1.045000 ;
      RECT  7.690000  0.085000  8.020000 0.545000 ;
      RECT  7.770000  2.105000  7.940000 2.375000 ;
      RECT  7.980000  1.005000  8.150000 1.215000 ;
      RECT  8.150000  2.175000  8.570000 2.635000 ;
      RECT  8.230000  0.275000  8.610000 0.445000 ;
      RECT  8.230000  0.445000  8.540000 0.835000 ;
      RECT  8.230000  1.765000  8.540000 1.835000 ;
      RECT  8.230000  1.835000  8.985000 2.005000 ;
      RECT  8.370000  0.835000  8.540000 1.595000 ;
      RECT  8.710000  0.705000  8.970000 1.495000 ;
      RECT  8.710000  1.495000  9.445000 1.660000 ;
      RECT  8.710000  1.660000  9.845000 1.665000 ;
      RECT  8.780000  0.255000  9.890000 0.535000 ;
      RECT  8.815000  2.005000  8.985000 2.465000 ;
      RECT  9.185000  1.665000  9.845000 1.955000 ;
      RECT  9.195000  2.125000 10.215000 2.465000 ;
      RECT  9.235000  0.920000  9.405000 1.325000 ;
      RECT  9.670000  0.535000  9.890000 1.315000 ;
      RECT  9.670000  1.315000 10.285000 1.485000 ;
      RECT 10.040000  1.485000 10.285000 1.575000 ;
      RECT 10.040000  1.575000 11.370000 1.745000 ;
      RECT 10.040000  1.745000 10.215000 2.125000 ;
      RECT 10.110000  0.085000 10.330000 0.525000 ;
      RECT 10.150000  0.695000 10.730000 0.865000 ;
      RECT 10.150000  0.865000 10.370000 1.145000 ;
      RECT 10.415000  2.195000 10.665000 2.635000 ;
      RECT 10.560000  0.295000 11.735000 0.465000 ;
      RECT 10.560000  0.465000 10.730000 0.695000 ;
      RECT 10.600000  1.065000 11.370000 1.275000 ;
      RECT 10.910000  1.915000 11.730000 2.085000 ;
      RECT 10.910000  2.085000 11.080000 2.375000 ;
      RECT 11.065000  0.635000 11.370000 1.065000 ;
      RECT 11.255000  2.255000 11.635000 2.635000 ;
      RECT 11.560000  0.465000 11.735000 0.995000 ;
      RECT 11.560000  0.995000 12.205000 1.325000 ;
      RECT 11.560000  1.325000 11.730000 1.915000 ;
      RECT 11.905000  0.085000 12.190000 0.710000 ;
      RECT 11.905000  1.495000 12.190000 2.635000 ;
      RECT 12.940000  0.255000 13.110000 0.635000 ;
      RECT 12.940000  0.635000 13.605000 0.805000 ;
      RECT 12.940000  1.535000 13.605000 1.705000 ;
      RECT 12.940000  1.705000 13.110000 2.465000 ;
      RECT 13.285000  0.085000 13.695000 0.465000 ;
      RECT 13.285000  1.875000 13.695000 2.635000 ;
      RECT 13.435000  0.805000 13.605000 0.995000 ;
      RECT 13.435000  0.995000 13.765000 1.325000 ;
      RECT 13.435000  1.325000 13.605000 1.535000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.855000  1.105000  1.025000 1.275000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.135000  1.785000  1.305000 1.955000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.480000  1.105000  5.650000 1.275000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.950000  1.785000  6.120000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.255000  0.765000  7.425000 0.935000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.615000  0.765000  7.785000 0.935000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.235000  1.105000  9.405000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.565000  1.785000  9.735000 1.955000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.175000  0.765000 11.345000 0.935000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT 0.795000 1.075000 1.085000 1.120000 ;
      RECT 0.795000 1.120000 9.465000 1.260000 ;
      RECT 0.795000 1.260000 1.085000 1.305000 ;
      RECT 1.070000 1.755000 1.370000 1.800000 ;
      RECT 1.070000 1.800000 9.795000 1.940000 ;
      RECT 1.070000 1.940000 1.370000 1.985000 ;
      RECT 5.420000 1.075000 5.710000 1.120000 ;
      RECT 5.420000 1.260000 5.710000 1.305000 ;
      RECT 5.890000 1.755000 6.180000 1.800000 ;
      RECT 5.890000 1.940000 6.180000 1.985000 ;
      RECT 9.155000 1.075000 9.465000 1.120000 ;
      RECT 9.155000 1.260000 9.465000 1.305000 ;
      RECT 9.500000 1.755000 9.795000 1.800000 ;
      RECT 9.500000 1.940000 9.795000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrbp_1


MACRO sky130_fd_sc_hdll__a222oi_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.000000 3.305000 1.330000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.475000 1.000000 3.995000 1.330000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415000 1.000000 2.735000 1.330000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 1.000000 2.245000 1.330000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.000000 0.595000 1.315000 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765000 1.000000 1.235000 1.315000 ;
    END
  END C2
  PIN Y
    ANTENNADIFFAREA  0.981600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.255000 0.425000 0.645000 ;
        RECT 0.095000 0.645000 2.975000 0.815000 ;
        RECT 0.095000 1.485000 1.655000 1.795000 ;
        RECT 0.095000 1.795000 0.345000 2.295000 ;
        RECT 1.405000 0.815000 1.655000 1.485000 ;
        RECT 2.410000 0.295000 2.975000 0.645000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.565000  2.055000 0.895000 2.295000 ;
      RECT 0.565000  2.295000 2.465000 2.465000 ;
      RECT 0.925000  0.085000 1.705000 0.465000 ;
      RECT 1.825000  1.500000 4.025000 1.735000 ;
      RECT 1.825000  1.735000 2.935000 1.830000 ;
      RECT 2.170000  2.135000 2.465000 2.295000 ;
      RECT 2.685000  1.830000 2.935000 2.250000 ;
      RECT 3.155000  1.905000 3.485000 2.635000 ;
      RECT 3.555000  0.085000 3.965000 0.815000 ;
      RECT 3.765000  1.735000 4.025000 2.250000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a222oi_1


MACRO sky130_fd_sc_hdll__nand3_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.330000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.170000 1.075000 2.615000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 1.075000 4.000000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.078000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 0.895000 1.445000 ;
        RECT 0.515000 1.445000 3.295000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.465000 ;
        RECT 1.455000 1.665000 1.835000 2.465000 ;
        RECT 2.915000 1.665000 3.295000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.295000 2.305000 0.465000 ;
      RECT 0.090000  0.465000 0.345000 0.785000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 1.115000  1.835000 1.285000 2.635000 ;
      RECT 1.455000  0.635000 3.295000 0.905000 ;
      RECT 2.055000  1.835000 2.745000 2.635000 ;
      RECT 2.495000  0.085000 2.825000 0.465000 ;
      RECT 3.515000  0.085000 3.895000 0.885000 ;
      RECT 3.515000  1.445000 3.895000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3_2


MACRO sky130_fd_sc_hdll__nand3_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 0.995000 1.905000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.915000 0.765000 1.285000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.745000 0.330000 1.325000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.761500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 1.895000 0.595000 ;
        RECT 0.515000 0.595000 0.745000 1.495000 ;
        RECT 0.515000 1.495000 1.895000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.465000 ;
        RECT 1.515000 0.595000 1.895000 0.825000 ;
        RECT 1.515000 1.665000 1.895000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.575000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 1.115000  1.835000 1.345000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3_1


MACRO sky130_fd_sc_hdll__nand3_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.900000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.250000 1.075000 6.370000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275000 1.075000 4.025000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.850000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  2.156000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.445000 6.785000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.465000 ;
        RECT 1.455000 1.665000 1.835000 2.465000 ;
        RECT 2.395000 1.665000 2.775000 2.465000 ;
        RECT 3.335000 1.665000 3.715000 2.465000 ;
        RECT 4.795000 0.655000 6.785000 0.905000 ;
        RECT 4.795000 1.665000 5.175000 2.465000 ;
        RECT 5.735000 1.665000 6.115000 2.465000 ;
        RECT 6.555000 0.905000 6.785000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 4.185000 0.905000 ;
      RECT 0.090000  1.445000 0.345000 2.635000 ;
      RECT 0.645000  0.085000 0.815000 0.565000 ;
      RECT 0.985000  0.255000 1.365000 0.735000 ;
      RECT 1.115000  1.835000 1.285000 2.635000 ;
      RECT 1.585000  0.085000 1.755000 0.565000 ;
      RECT 1.925000  0.655000 2.305000 0.735000 ;
      RECT 2.055000  1.835000 2.225000 2.635000 ;
      RECT 2.395000  0.255000 6.600000 0.485000 ;
      RECT 2.865000  0.655000 3.245000 0.735000 ;
      RECT 2.995000  1.835000 3.165000 2.635000 ;
      RECT 3.805000  0.655000 4.185000 0.735000 ;
      RECT 3.935000  1.835000 4.625000 2.635000 ;
      RECT 5.395000  1.835000 5.565000 2.635000 ;
      RECT 6.335000  1.835000 6.600000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3_4


MACRO sky130_fd_sc_hdll__nand3b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.825000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 0.995000 1.795000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 0.995000 1.335000 1.325000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.775200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.180000 1.495000 2.675000 1.665000 ;
        RECT 1.180000 1.665000 1.560000 2.465000 ;
        RECT 2.130000 0.255000 2.675000 0.485000 ;
        RECT 2.130000 1.665000 2.675000 2.465000 ;
        RECT 2.410000 0.485000 2.675000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.445000 0.510000 0.655000 ;
      RECT 0.085000  0.655000 2.220000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.595000 ;
      RECT 0.085000  1.595000 0.510000 1.925000 ;
      RECT 0.760000  0.085000 1.090000 0.485000 ;
      RECT 0.760000  1.495000 1.010000 2.635000 ;
      RECT 1.790000  1.835000 1.960000 2.635000 ;
      RECT 2.000000  0.825000 2.220000 1.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3b_1


MACRO sky130_fd_sc_hdll__nand3b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.820000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.075000 0.830000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.075000 4.930000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.185000 1.075000 7.100000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  2.156000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 0.635000 3.215000 0.905000 ;
        RECT 1.505000 1.445000 7.105000 1.665000 ;
        RECT 1.505000 1.665000 1.885000 2.465000 ;
        RECT 2.445000 1.665000 3.765000 2.005000 ;
        RECT 2.445000 2.005000 2.825000 2.465000 ;
        RECT 3.045000 0.905000 3.215000 1.075000 ;
        RECT 3.045000 1.075000 3.555000 1.445000 ;
        RECT 3.385000 2.005000 3.765000 2.465000 ;
        RECT 4.325000 1.665000 4.705000 2.465000 ;
        RECT 5.785000 1.665000 6.165000 2.465000 ;
        RECT 6.725000 1.665000 7.105000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.255000 0.425000 0.715000 ;
      RECT 0.085000  0.715000 1.335000 0.905000 ;
      RECT 0.085000  0.905000 0.260000 1.445000 ;
      RECT 0.085000  1.445000 0.425000 2.465000 ;
      RECT 0.645000  0.085000 0.895000 0.545000 ;
      RECT 0.645000  1.445000 1.335000 2.635000 ;
      RECT 1.055000  0.905000 1.335000 1.075000 ;
      RECT 1.055000  1.075000 2.825000 1.275000 ;
      RECT 1.085000  0.255000 5.175000 0.465000 ;
      RECT 2.105000  1.835000 2.275000 2.635000 ;
      RECT 3.045000  2.175000 3.215000 2.635000 ;
      RECT 3.385000  0.635000 5.175000 0.715000 ;
      RECT 3.385000  0.715000 7.105000 0.905000 ;
      RECT 3.985000  1.835000 4.155000 2.635000 ;
      RECT 4.925000  1.835000 5.615000 2.635000 ;
      RECT 5.365000  0.085000 5.615000 0.545000 ;
      RECT 5.785000  0.255000 6.165000 0.715000 ;
      RECT 6.385000  0.085000 6.555000 0.545000 ;
      RECT 6.385000  1.835000 6.555000 2.635000 ;
      RECT 6.725000  0.255000 7.105000 0.715000 ;
      RECT 7.325000  0.085000 7.655000 0.905000 ;
      RECT 7.325000  1.445000 7.655000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3b_4


MACRO sky130_fd_sc_hdll__nand3b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.075000 0.830000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.150000 1.075000 3.440000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.890000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.110500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.110000 1.785000 4.490000 1.955000 ;
        RECT 1.110000 1.955000 2.430000 2.005000 ;
        RECT 1.110000 2.005000 1.490000 2.465000 ;
        RECT 2.050000 2.005000 2.430000 2.465000 ;
        RECT 3.560000 0.635000 4.490000 0.905000 ;
        RECT 3.560000 1.955000 4.490000 2.005000 ;
        RECT 3.560000 2.005000 3.860000 2.465000 ;
        RECT 4.250000 0.905000 4.490000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.255000 0.410000 0.655000 ;
      RECT 0.090000  0.655000 0.260000 1.445000 ;
      RECT 0.090000  1.445000 4.000000 1.615000 ;
      RECT 0.090000  1.615000 0.260000 2.065000 ;
      RECT 0.090000  2.065000 0.410000 2.465000 ;
      RECT 0.630000  0.085000 0.940000 0.905000 ;
      RECT 0.630000  1.835000 0.940000 2.635000 ;
      RECT 1.110000  0.255000 1.490000 0.715000 ;
      RECT 1.110000  0.715000 3.000000 0.905000 ;
      RECT 1.710000  0.085000 1.960000 0.545000 ;
      RECT 1.710000  2.175000 1.880000 2.635000 ;
      RECT 2.200000  0.255000 4.450000 0.465000 ;
      RECT 2.200000  0.635000 3.000000 0.715000 ;
      RECT 2.650000  2.175000 2.900000 2.635000 ;
      RECT 3.090000  2.175000 3.390000 2.635000 ;
      RECT 3.220000  0.465000 3.390000 0.905000 ;
      RECT 3.670000  1.075000 4.000000 1.445000 ;
      RECT 4.160000  2.175000 4.450000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3b_2


MACRO sky130_fd_sc_hdll__probe_p_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.832500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.240000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1.250000 0.560000 4.270000 2.160000 ;
      LAYER via4 ;
        RECT 1.560000 0.870000 2.360000 1.670000 ;
        RECT 3.160000 0.870000 3.960000 1.670000 ;
    END
  END X
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.615000  0.085000 0.895000 0.565000 ;
        RECT 1.505000  0.085000 1.805000 0.565000 ;
        RECT 2.475000  0.085000 2.745000 0.565000 ;
        RECT 3.415000  0.085000 3.685000 0.565000 ;
        RECT 4.355000  0.085000 4.625000 0.565000 ;
        RECT 5.295000  0.085000 5.545000 0.885000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.595000 1.835000 0.865000 2.635000 ;
        RECT 1.535000 1.835000 1.805000 2.635000 ;
        RECT 2.475000 1.835000 2.745000 2.635000 ;
        RECT 3.415000 1.835000 3.685000 2.635000 ;
        RECT 4.355000 1.835000 4.625000 2.635000 ;
        RECT 5.295000 1.485000 5.595000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 1.445000 1.595000 1.615000 ;
      RECT 0.095000 1.615000 0.425000 2.465000 ;
      RECT 0.145000 0.255000 0.445000 0.735000 ;
      RECT 0.145000 0.735000 1.595000 0.905000 ;
      RECT 1.035000 1.615000 1.365000 2.465000 ;
      RECT 1.065000 0.255000 1.335000 0.735000 ;
      RECT 1.420000 0.905000 1.595000 1.075000 ;
      RECT 1.420000 1.075000 4.045000 1.245000 ;
      RECT 1.420000 1.245000 1.595000 1.445000 ;
      RECT 1.975000 0.255000 2.305000 0.735000 ;
      RECT 1.975000 0.735000 5.125000 0.905000 ;
      RECT 1.975000 1.445000 5.125000 1.615000 ;
      RECT 1.975000 1.615000 2.305000 2.465000 ;
      RECT 2.915000 0.255000 3.245000 0.735000 ;
      RECT 2.915000 1.615000 3.245000 2.465000 ;
      RECT 3.855000 0.255000 4.185000 0.735000 ;
      RECT 3.855000 1.615000 4.185000 2.465000 ;
      RECT 4.290000 0.905000 5.125000 1.445000 ;
      RECT 4.795000 0.255000 5.125000 0.735000 ;
      RECT 4.795000 1.615000 5.125000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.560000  1.105000 4.730000 1.275000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 4.920000  1.105000 5.090000 1.275000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 3.465000 1.060000 4.105000 1.320000 ;
      RECT 4.105000 1.075000 5.150000 1.305000 ;
    LAYER met2 ;
      RECT 3.445000 1.005000 4.125000 1.375000 ;
      RECT 3.465000 1.060000 4.105000 1.320000 ;
    LAYER met3 ;
      RECT 3.395000 1.025000 3.420000 1.355000 ;
      RECT 3.395000 1.030000 4.175000 1.350000 ;
      RECT 3.420000 1.025000 4.150000 1.355000 ;
      RECT 4.150000 1.025000 4.175000 1.355000 ;
    LAYER met4 ;
      RECT 1.370000 0.680000 4.150000 1.860000 ;
      RECT 3.420000 1.025000 4.150000 1.355000 ;
    LAYER via ;
      RECT 3.550000 1.115000 3.700000 1.265000 ;
      RECT 3.870000 1.115000 4.020000 1.265000 ;
    LAYER via2 ;
      RECT 3.485000 1.090000 3.685000 1.290000 ;
      RECT 3.885000 1.090000 4.085000 1.290000 ;
    LAYER via3 ;
      RECT 3.485000 1.090000 3.685000 1.290000 ;
      RECT 3.885000 1.090000 4.085000 1.290000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__probe_p_8


MACRO sky130_fd_sc_hdll__a31o_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385000 0.415000 2.615000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.905000 0.400000 2.155000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 0.760000 1.370000 0.995000 ;
        RECT 1.030000 0.995000 1.545000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.195000 0.755000 3.535000 1.325000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.715000 0.815000 0.885000 ;
        RECT 0.090000 0.885000 0.345000 1.835000 ;
        RECT 0.090000 1.835000 0.815000 2.005000 ;
        RECT 0.645000 0.255000 0.815000 0.715000 ;
        RECT 0.645000 2.005000 0.815000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.465000 ;
      RECT 0.135000  2.175000 0.385000 2.635000 ;
      RECT 0.515000  1.075000 0.845000 1.245000 ;
      RECT 0.515000  1.245000 0.685000 1.495000 ;
      RECT 0.515000  1.495000 3.345000 1.665000 ;
      RECT 0.985000  1.835000 1.285000 2.635000 ;
      RECT 1.005000  0.085000 1.385000 0.465000 ;
      RECT 1.455000  1.835000 2.895000 2.005000 ;
      RECT 1.455000  2.005000 1.755000 2.425000 ;
      RECT 2.015000  2.175000 2.345000 2.635000 ;
      RECT 2.585000  2.005000 2.895000 2.425000 ;
      RECT 2.785000  0.255000 2.955000 1.495000 ;
      RECT 3.175000  0.085000 3.465000 0.565000 ;
      RECT 3.175000  1.665000 3.345000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31o_2


MACRO sky130_fd_sc_hdll__a31o_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.995000 2.275000 1.655000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 0.995000 1.815000 1.655000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 0.995000 1.340000 1.325000 ;
        RECT 1.075000 1.325000 1.340000 1.655000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.995000 2.745000 1.655000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.447300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.300000 0.425000 0.810000 ;
        RECT 0.095000 0.810000 0.285000 1.575000 ;
        RECT 0.095000 1.575000 0.425000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.455000  0.995000 0.815000 1.325000 ;
      RECT 0.605000  0.085000 0.935000 0.485000 ;
      RECT 0.645000  0.655000 3.085000 0.825000 ;
      RECT 0.645000  0.825000 0.815000 0.995000 ;
      RECT 0.645000  1.495000 0.895000 2.635000 ;
      RECT 1.085000  1.825000 2.525000 1.995000 ;
      RECT 1.085000  1.995000 1.385000 2.415000 ;
      RECT 1.665000  2.165000 1.995000 2.635000 ;
      RECT 2.125000  0.315000 2.505000 0.655000 ;
      RECT 2.275000  1.995000 2.525000 2.415000 ;
      RECT 2.725000  0.085000 3.055000 0.485000 ;
      RECT 2.755000  1.825000 3.085000 2.425000 ;
      RECT 2.915000  0.825000 3.085000 1.825000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31o_1


MACRO sky130_fd_sc_hdll__a31o_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.900000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 1.075000 1.855000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.775000 0.735000 2.370000 0.905000 ;
        RECT 0.775000 0.905000 1.255000 1.275000 ;
        RECT 2.185000 0.905000 2.370000 1.075000 ;
        RECT 2.185000 1.075000 2.565000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.075000 0.525000 1.445000 ;
        RECT 0.145000 1.445000 3.155000 1.615000 ;
        RECT 2.775000 1.075000 3.155000 1.445000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.925000 1.075000 4.455000 1.285000 ;
        RECT 4.215000 0.745000 4.455000 1.075000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.905000 0.655000 6.780000 0.825000 ;
        RECT 4.935000 1.785000 6.780000 1.955000 ;
        RECT 5.045000 1.955000 5.215000 2.465000 ;
        RECT 5.985000 1.955000 6.155000 2.465000 ;
        RECT 6.585000 0.825000 6.780000 1.785000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.175000  0.085000 0.345000 0.905000 ;
      RECT 0.175000  1.785000 3.285000 1.955000 ;
      RECT 0.175000  1.955000 0.345000 2.465000 ;
      RECT 0.515000  2.125000 0.895000 2.635000 ;
      RECT 1.115000  1.955000 1.285000 2.465000 ;
      RECT 1.455000  0.395000 2.770000 0.565000 ;
      RECT 1.455000  2.125000 1.835000 2.635000 ;
      RECT 2.055000  1.955000 2.225000 2.465000 ;
      RECT 2.395000  2.125000 2.775000 2.635000 ;
      RECT 2.600000  0.565000 2.770000 0.700000 ;
      RECT 2.600000  0.700000 3.835000 0.805000 ;
      RECT 2.600000  0.805000 3.695000 0.870000 ;
      RECT 2.950000  0.085000 3.285000 0.530000 ;
      RECT 3.115000  1.955000 3.285000 2.295000 ;
      RECT 3.115000  2.295000 4.225000 2.465000 ;
      RECT 3.455000  0.295000 3.835000 0.700000 ;
      RECT 3.455000  0.870000 3.695000 1.455000 ;
      RECT 3.455000  1.455000 4.820000 1.625000 ;
      RECT 3.455000  1.625000 3.835000 2.115000 ;
      RECT 4.055000  1.795000 4.225000 2.295000 ;
      RECT 4.135000  0.085000 4.665000 0.565000 ;
      RECT 4.495000  2.125000 4.825000 2.635000 ;
      RECT 4.650000  0.995000 6.355000 1.325000 ;
      RECT 4.650000  1.325000 4.820000 1.455000 ;
      RECT 5.385000  0.085000 5.765000 0.485000 ;
      RECT 5.385000  2.125000 5.765000 2.635000 ;
      RECT 6.325000  0.085000 6.705000 0.485000 ;
      RECT 6.325000  2.125000 6.705000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31o_4


MACRO sky130_fd_sc_hdll__sdlclkp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.820000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.950000 1.075000 5.240000 1.120000 ;
        RECT 4.950000 1.120000 6.230000 1.260000 ;
        RECT 4.950000 1.260000 5.240000 1.305000 ;
        RECT 5.940000 1.075000 6.230000 1.120000 ;
        RECT 5.940000 1.260000 6.230000 1.305000 ;
    END
  END CLK
  PIN GATE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.890000 0.955000 1.295000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.840000 0.255000 7.170000 0.445000 ;
        RECT 6.970000 0.445000 7.170000 0.715000 ;
        RECT 6.970000 0.715000 7.675000 0.885000 ;
        RECT 6.970000 1.485000 7.675000 1.655000 ;
        RECT 6.970000 1.655000 7.220000 2.465000 ;
        RECT 7.490000 0.885000 7.675000 1.485000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.330000 1.665000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.295000 0.785000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  0.085000 0.895000 0.445000 ;
      RECT 0.515000  0.785000 0.720000 2.125000 ;
      RECT 0.515000  2.125000 1.280000 2.465000 ;
      RECT 1.115000  0.255000 1.295000 0.615000 ;
      RECT 1.465000  0.255000 2.645000 0.535000 ;
      RECT 1.465000  0.705000 1.800000 1.205000 ;
      RECT 1.465000  1.205000 1.960000 1.955000 ;
      RECT 1.610000  2.125000 2.300000 2.465000 ;
      RECT 1.970000  0.705000 2.305000 1.035000 ;
      RECT 2.130000  1.205000 3.205000 1.375000 ;
      RECT 2.130000  1.375000 2.300000 2.125000 ;
      RECT 2.470000  1.575000 2.665000 1.635000 ;
      RECT 2.470000  1.635000 3.545000 1.905000 ;
      RECT 2.475000  0.535000 2.645000 0.995000 ;
      RECT 2.475000  0.995000 3.205000 1.205000 ;
      RECT 2.520000  2.075000 3.105000 2.635000 ;
      RECT 2.910000  0.085000 3.080000 0.825000 ;
      RECT 3.325000  1.905000 3.545000 1.915000 ;
      RECT 3.325000  1.915000 5.755000 2.085000 ;
      RECT 3.325000  2.085000 3.545000 2.465000 ;
      RECT 3.375000  0.255000 3.545000 1.635000 ;
      RECT 3.735000  0.255000 4.065000 0.765000 ;
      RECT 3.735000  0.765000 4.160000 0.935000 ;
      RECT 3.735000  0.935000 3.905000 1.575000 ;
      RECT 3.735000  1.575000 4.145000 1.745000 ;
      RECT 3.885000  2.255000 5.755000 2.635000 ;
      RECT 4.075000  1.105000 4.670000 1.275000 ;
      RECT 4.285000  0.085000 4.615000 0.445000 ;
      RECT 4.365000  1.275000 4.670000 1.495000 ;
      RECT 4.365000  1.495000 5.215000 1.745000 ;
      RECT 4.380000  0.615000 5.085000 0.785000 ;
      RECT 4.380000  0.785000 4.670000 1.105000 ;
      RECT 4.835000  0.255000 5.085000 0.615000 ;
      RECT 4.965000  0.995000 5.185000 1.325000 ;
      RECT 5.405000  0.995000 5.755000 1.915000 ;
      RECT 5.505000  0.255000 5.675000 0.615000 ;
      RECT 5.505000  0.615000 6.750000 0.785000 ;
      RECT 5.975000  0.995000 6.405000 1.325000 ;
      RECT 5.975000  1.495000 6.750000 2.085000 ;
      RECT 5.975000  2.085000 6.145000 2.465000 ;
      RECT 6.335000  0.085000 6.670000 0.445000 ;
      RECT 6.395000  2.255000 6.725000 2.635000 ;
      RECT 6.580000  0.785000 6.750000 1.055000 ;
      RECT 6.580000  1.055000 7.270000 1.315000 ;
      RECT 6.580000  1.315000 6.750000 1.495000 ;
      RECT 7.390000  0.085000 7.560000 0.545000 ;
      RECT 7.440000  1.825000 7.690000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.625000  1.445000 1.795000 1.615000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.135000  0.765000 2.305000 0.935000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 3.990000  0.765000 4.160000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.500000  1.445000 4.670000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.010000  1.105000 5.180000 1.275000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.000000  1.105000 6.170000 1.275000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 1.565000 1.415000 1.855000 1.460000 ;
      RECT 1.565000 1.460000 4.730000 1.600000 ;
      RECT 1.565000 1.600000 1.855000 1.645000 ;
      RECT 2.075000 0.735000 2.365000 0.780000 ;
      RECT 2.075000 0.780000 4.220000 0.920000 ;
      RECT 2.075000 0.920000 2.365000 0.965000 ;
      RECT 3.930000 0.735000 4.220000 0.780000 ;
      RECT 3.930000 0.920000 4.220000 0.965000 ;
      RECT 4.440000 1.415000 4.730000 1.460000 ;
      RECT 4.440000 1.600000 4.730000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdlclkp_2


MACRO sky130_fd_sc_hdll__sdlclkp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.360000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.745000 1.075000 5.035000 1.120000 ;
        RECT 4.745000 1.120000 6.230000 1.260000 ;
        RECT 4.745000 1.260000 5.035000 1.305000 ;
        RECT 5.940000 1.075000 6.230000 1.120000 ;
        RECT 5.940000 1.260000 6.230000 1.305000 ;
    END
  END CLK
  PIN GATE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 0.955000 1.235000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.480200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.985000 0.255000 7.235000 2.465000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.330000 1.665000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.295000 0.785000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  0.085000 0.895000 0.445000 ;
      RECT 0.515000  0.785000 0.685000 2.125000 ;
      RECT 0.515000  2.125000 1.280000 2.465000 ;
      RECT 1.115000  0.255000 1.295000 0.615000 ;
      RECT 1.465000  0.255000 2.645000 0.535000 ;
      RECT 1.465000  0.705000 1.800000 1.205000 ;
      RECT 1.465000  1.205000 1.960000 1.955000 ;
      RECT 1.610000  2.125000 2.300000 2.465000 ;
      RECT 1.970000  0.705000 2.305000 1.035000 ;
      RECT 2.130000  1.205000 3.205000 1.375000 ;
      RECT 2.130000  1.375000 2.300000 2.125000 ;
      RECT 2.470000  1.575000 2.665000 1.635000 ;
      RECT 2.470000  1.635000 3.545000 1.905000 ;
      RECT 2.475000  0.535000 2.645000 0.995000 ;
      RECT 2.475000  0.995000 3.205000 1.205000 ;
      RECT 2.520000  2.075000 3.105000 2.635000 ;
      RECT 2.910000  0.085000 3.080000 0.825000 ;
      RECT 3.325000  1.905000 3.545000 1.915000 ;
      RECT 3.325000  1.915000 5.735000 2.085000 ;
      RECT 3.325000  2.085000 3.545000 2.465000 ;
      RECT 3.375000  0.255000 3.545000 1.635000 ;
      RECT 3.735000  0.255000 4.065000 0.935000 ;
      RECT 3.735000  0.935000 3.905000 1.575000 ;
      RECT 3.735000  1.575000 4.145000 1.745000 ;
      RECT 3.885000  2.255000 5.735000 2.635000 ;
      RECT 4.075000  1.105000 4.550000 1.275000 ;
      RECT 4.285000  0.085000 4.615000 0.445000 ;
      RECT 4.365000  1.275000 4.550000 1.495000 ;
      RECT 4.365000  1.495000 5.215000 1.745000 ;
      RECT 4.380000  0.615000 5.215000 0.785000 ;
      RECT 4.380000  0.785000 4.550000 1.105000 ;
      RECT 4.745000  0.995000 5.060000 1.325000 ;
      RECT 4.965000  0.255000 5.215000 0.615000 ;
      RECT 5.385000  0.995000 5.735000 1.915000 ;
      RECT 5.535000  0.255000 5.705000 0.615000 ;
      RECT 5.535000  0.615000 6.815000 0.785000 ;
      RECT 5.955000  0.995000 6.395000 1.325000 ;
      RECT 5.955000  1.495000 6.815000 2.085000 ;
      RECT 5.955000  2.085000 6.125000 2.465000 ;
      RECT 6.325000  0.085000 6.685000 0.445000 ;
      RECT 6.385000  2.255000 6.715000 2.635000 ;
      RECT 6.645000  0.785000 6.815000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.625000  1.445000 1.795000 1.615000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.135000  0.765000 2.305000 0.935000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.800000  0.765000 3.970000 0.935000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.365000  1.445000 4.535000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 4.805000  1.105000 4.975000 1.275000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.000000  1.105000 6.170000 1.275000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 1.565000 1.415000 1.855000 1.460000 ;
      RECT 1.565000 1.460000 4.595000 1.600000 ;
      RECT 1.565000 1.600000 1.855000 1.645000 ;
      RECT 2.075000 0.735000 2.365000 0.780000 ;
      RECT 2.075000 0.780000 4.030000 0.920000 ;
      RECT 2.075000 0.920000 2.365000 0.965000 ;
      RECT 3.740000 0.735000 4.030000 0.780000 ;
      RECT 3.740000 0.920000 4.030000 0.965000 ;
      RECT 4.305000 1.415000 4.595000 1.460000 ;
      RECT 4.305000 1.600000 4.595000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdlclkp_1


MACRO sky130_fd_sc_hdll__sdlclkp_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.200000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.055000 1.075000 5.345000 1.120000 ;
        RECT 5.055000 1.120000 6.390000 1.260000 ;
        RECT 5.055000 1.260000 5.345000 1.305000 ;
        RECT 6.100000 1.075000 6.390000 1.120000 ;
        RECT 6.100000 1.260000 6.390000 1.305000 ;
    END
  END CLK
  PIN GATE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.905000 0.955000 1.295000 1.445000 ;
        RECT 0.905000 1.445000 1.340000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.251200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.000000 0.255000 7.380000 0.445000 ;
        RECT 7.130000 0.445000 7.380000 0.715000 ;
        RECT 7.130000 0.715000 7.820000 0.885000 ;
        RECT 7.130000 1.485000 7.820000 1.655000 ;
        RECT 7.130000 1.655000 7.380000 2.465000 ;
        RECT 7.650000 0.885000 7.820000 1.055000 ;
        RECT 7.650000 1.055000 9.055000 1.315000 ;
        RECT 7.650000 1.315000 7.820000 1.485000 ;
        RECT 8.205000 0.255000 8.595000 1.055000 ;
        RECT 8.205000 1.315000 8.595000 2.465000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.345000 1.665000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.295000 0.785000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  0.085000 0.895000 0.445000 ;
      RECT 0.515000  0.785000 0.735000 2.125000 ;
      RECT 0.515000  2.125000 1.360000 2.465000 ;
      RECT 1.115000  0.255000 1.295000 0.615000 ;
      RECT 1.465000  0.255000 2.700000 0.535000 ;
      RECT 1.465000  0.705000 1.855000 1.205000 ;
      RECT 1.465000  1.205000 2.015000 1.325000 ;
      RECT 1.510000  1.325000 2.015000 1.955000 ;
      RECT 1.530000  2.125000 2.405000 2.465000 ;
      RECT 2.025000  0.705000 2.360000 1.035000 ;
      RECT 2.235000  1.205000 3.265000 1.375000 ;
      RECT 2.235000  1.375000 2.405000 2.125000 ;
      RECT 2.530000  0.535000 2.700000 0.995000 ;
      RECT 2.530000  0.995000 3.265000 1.205000 ;
      RECT 2.575000  1.575000 2.795000 1.635000 ;
      RECT 2.575000  1.635000 3.705000 1.905000 ;
      RECT 2.575000  2.075000 3.265000 2.635000 ;
      RECT 2.920000  0.085000 3.265000 0.825000 ;
      RECT 3.485000  0.255000 3.705000 1.635000 ;
      RECT 3.485000  1.905000 3.705000 1.915000 ;
      RECT 3.485000  1.915000 5.915000 2.085000 ;
      RECT 3.485000  2.085000 3.705000 2.465000 ;
      RECT 3.895000  0.255000 4.225000 0.765000 ;
      RECT 3.895000  0.765000 4.320000 0.935000 ;
      RECT 3.895000  0.935000 4.065000 1.575000 ;
      RECT 3.895000  1.575000 4.305000 1.745000 ;
      RECT 3.895000  2.255000 5.915000 2.635000 ;
      RECT 4.235000  1.105000 4.830000 1.275000 ;
      RECT 4.395000  0.085000 4.775000 0.445000 ;
      RECT 4.525000  1.275000 4.830000 1.495000 ;
      RECT 4.525000  1.495000 5.375000 1.745000 ;
      RECT 4.540000  0.615000 5.245000 0.785000 ;
      RECT 4.540000  0.785000 4.830000 1.105000 ;
      RECT 4.995000  0.255000 5.245000 0.615000 ;
      RECT 5.055000  0.995000 5.345000 1.325000 ;
      RECT 5.415000  0.255000 5.835000 0.615000 ;
      RECT 5.415000  0.615000 6.910000 0.785000 ;
      RECT 5.565000  0.995000 5.915000 1.915000 ;
      RECT 6.005000  0.085000 6.830000 0.445000 ;
      RECT 6.135000  0.995000 6.565000 1.325000 ;
      RECT 6.135000  1.495000 6.910000 2.085000 ;
      RECT 6.135000  2.085000 6.305000 2.465000 ;
      RECT 6.555000  2.255000 6.885000 2.635000 ;
      RECT 6.740000  0.785000 6.910000 1.055000 ;
      RECT 6.740000  1.055000 7.430000 1.315000 ;
      RECT 6.740000  1.315000 6.910000 1.495000 ;
      RECT 7.600000  0.085000 7.850000 0.545000 ;
      RECT 7.600000  1.825000 7.850000 2.635000 ;
      RECT 8.765000  0.085000 9.035000 0.885000 ;
      RECT 8.765000  1.485000 9.035000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.680000  1.445000 1.850000 1.615000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.190000  0.765000 2.360000 0.935000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.150000  0.765000 4.320000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.660000  1.445000 4.830000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.115000  1.105000 5.285000 1.275000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.160000  1.105000 6.330000 1.275000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 1.620000 1.415000 1.910000 1.460000 ;
      RECT 1.620000 1.460000 4.890000 1.600000 ;
      RECT 1.620000 1.600000 1.910000 1.645000 ;
      RECT 2.130000 0.735000 2.420000 0.780000 ;
      RECT 2.130000 0.780000 4.380000 0.920000 ;
      RECT 2.130000 0.920000 2.420000 0.965000 ;
      RECT 4.090000 0.735000 4.380000 0.780000 ;
      RECT 4.090000 0.920000 4.380000 0.965000 ;
      RECT 4.600000 1.415000 4.890000 1.460000 ;
      RECT 4.600000 1.600000 4.890000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdlclkp_4


MACRO sky130_fd_sc_hdll__sdfxbp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  13.34000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.755000 1.355000 3.125000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.210000 0.255000 10.490000 2.455000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.515000 0.265000 12.785000 2.325000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 1.055000 4.345000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.860000 0.615000 3.535000 0.785000 ;
        RECT 1.860000 0.785000 2.030000 1.685000 ;
        RECT 3.315000 0.785000 3.535000 1.115000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.340000 0.085000 ;
      RECT  0.000000  2.635000 13.340000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.860000 0.805000 ;
      RECT  0.175000  1.795000  0.895000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.515000  2.135000  0.895000 2.635000 ;
      RECT  0.665000  0.805000  0.860000 0.970000 ;
      RECT  0.665000  0.970000  0.895000 1.795000 ;
      RECT  1.115000  0.345000  1.285000 2.465000 ;
      RECT  1.520000  0.255000  1.905000 0.445000 ;
      RECT  1.520000  0.445000  1.690000 1.860000 ;
      RECT  1.520000  1.860000  3.530000 2.075000 ;
      RECT  1.520000  2.075000  1.805000 2.445000 ;
      RECT  1.975000  2.245000  2.355000 2.635000 ;
      RECT  2.145000  0.085000  2.475000 0.445000 ;
      RECT  2.250000  0.955000  2.695000 1.125000 ;
      RECT  2.250000  1.125000  2.420000 1.860000 ;
      RECT  2.875000  2.245000  3.870000 2.415000 ;
      RECT  3.050000  0.275000  3.875000 0.445000 ;
      RECT  3.335000  1.355000  3.555000 1.685000 ;
      RECT  3.335000  1.685000  3.530000 1.860000 ;
      RECT  3.700000  1.825000  4.685000 1.995000 ;
      RECT  3.700000  1.995000  3.870000 2.245000 ;
      RECT  3.705000  0.445000  3.875000 0.715000 ;
      RECT  3.705000  0.715000  4.685000 0.885000 ;
      RECT  4.090000  2.165000  4.260000 2.635000 ;
      RECT  4.095000  0.085000  4.295000 0.545000 ;
      RECT  4.515000  0.365000  4.865000 0.535000 ;
      RECT  4.515000  0.535000  4.685000 0.715000 ;
      RECT  4.515000  0.885000  4.685000 1.825000 ;
      RECT  4.515000  1.995000  4.685000 2.070000 ;
      RECT  4.515000  2.070000  4.800000 2.440000 ;
      RECT  4.855000  0.705000  5.485000 1.035000 ;
      RECT  4.855000  1.035000  5.145000 1.905000 ;
      RECT  4.995000  2.190000  6.215000 2.360000 ;
      RECT  5.085000  0.365000  5.875000 0.535000 ;
      RECT  5.335000  1.655000  5.825000 2.010000 ;
      RECT  5.705000  0.535000  5.875000 1.315000 ;
      RECT  5.705000  1.315000  6.555000 1.485000 ;
      RECT  5.995000  1.485000  6.555000 1.575000 ;
      RECT  5.995000  1.575000  6.215000 2.190000 ;
      RECT  6.095000  0.765000  6.945000 1.065000 ;
      RECT  6.095000  1.065000  6.265000 1.095000 ;
      RECT  6.175000  0.085000  6.545000 0.585000 ;
      RECT  6.385000  1.245000  6.555000 1.315000 ;
      RECT  6.385000  1.835000  6.555000 2.635000 ;
      RECT  6.725000  0.365000  7.235000 0.535000 ;
      RECT  6.725000  0.535000  6.945000 0.765000 ;
      RECT  6.725000  1.065000  6.945000 2.135000 ;
      RECT  6.725000  2.135000  7.025000 2.465000 ;
      RECT  7.115000  0.705000  7.715000 1.035000 ;
      RECT  7.115000  1.245000  7.355000 1.965000 ;
      RECT  7.250000  2.165000  8.285000 2.335000 ;
      RECT  7.515000  0.365000  8.155000 0.535000 ;
      RECT  7.525000  1.035000  7.715000 1.575000 ;
      RECT  7.525000  1.575000  7.895000 1.905000 ;
      RECT  7.935000  0.535000  8.155000 0.995000 ;
      RECT  7.935000  0.995000  9.045000 1.325000 ;
      RECT  7.935000  1.325000  8.285000 1.405000 ;
      RECT  8.115000  1.405000  8.285000 2.165000 ;
      RECT  8.380000  0.085000  8.800000 0.615000 ;
      RECT  8.485000  1.575000  9.400000 1.905000 ;
      RECT  8.515000  2.135000  8.820000 2.635000 ;
      RECT  9.035000  0.300000  9.400000 0.825000 ;
      RECT  9.070000  1.905000  9.400000 2.455000 ;
      RECT  9.215000  0.825000  9.400000 0.995000 ;
      RECT  9.215000  0.995000 10.000000 1.325000 ;
      RECT  9.215000  1.325000  9.400000 1.575000 ;
      RECT  9.570000  0.085000  9.990000 0.695000 ;
      RECT  9.570000  1.625000  9.990000 2.635000 ;
      RECT 10.680000  0.085000 10.910000 0.690000 ;
      RECT 10.690000  1.615000 10.860000 2.635000 ;
      RECT 11.130000  0.345000 11.380000 0.995000 ;
      RECT 11.130000  0.995000 12.340000 1.325000 ;
      RECT 11.130000  1.325000 11.460000 2.425000 ;
      RECT 11.665000  0.085000 12.295000 0.805000 ;
      RECT 11.690000  1.495000 12.295000 2.635000 ;
      RECT 12.985000  0.085000 13.155000 0.955000 ;
      RECT 12.985000  1.395000 13.155000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.695000  1.785000  0.865000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.115000  0.425000  1.285000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.145000  0.765000  5.315000 0.935000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.615000  1.785000  5.785000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.175000  1.785000  7.345000 1.955000 ;
      RECT  7.185000  0.765000  7.355000 0.935000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
    LAYER met1 ;
      RECT 0.635000 1.755000 0.925000 1.800000 ;
      RECT 0.635000 1.800000 7.405000 1.940000 ;
      RECT 0.635000 1.940000 0.925000 1.985000 ;
      RECT 1.005000 0.395000 1.345000 0.440000 ;
      RECT 1.005000 0.440000 5.225000 0.580000 ;
      RECT 1.005000 0.580000 1.345000 0.625000 ;
      RECT 5.085000 0.580000 5.225000 0.735000 ;
      RECT 5.085000 0.735000 5.375000 0.780000 ;
      RECT 5.085000 0.780000 7.415000 0.920000 ;
      RECT 5.085000 0.920000 5.375000 0.965000 ;
      RECT 5.555000 1.755000 5.845000 1.800000 ;
      RECT 5.555000 1.940000 5.845000 1.985000 ;
      RECT 7.115000 1.755000 7.405000 1.800000 ;
      RECT 7.115000 1.940000 7.405000 1.985000 ;
      RECT 7.125000 0.735000 7.415000 0.780000 ;
      RECT 7.125000 0.920000 7.415000 0.965000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfxbp_2


MACRO sky130_fd_sc_hdll__sdfxbp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.96000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.755000 1.355000 3.125000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.960000 0.305000 10.440000 0.825000 ;
        RECT  9.980000 1.505000 10.440000 2.465000 ;
        RECT 10.220000 0.825000 10.440000 1.505000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.615000 0.265000 11.870000 2.325000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 1.055000 4.345000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.860000 0.615000 3.535000 0.785000 ;
        RECT 1.860000 0.785000 2.030000 1.685000 ;
        RECT 3.315000 0.785000 3.535000 1.115000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.860000 0.805000 ;
      RECT  0.175000  1.795000  0.895000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.515000  2.135000  0.895000 2.635000 ;
      RECT  0.665000  0.805000  0.860000 0.970000 ;
      RECT  0.665000  0.970000  0.895000 1.795000 ;
      RECT  1.115000  0.345000  1.285000 2.465000 ;
      RECT  1.520000  0.255000  1.905000 0.445000 ;
      RECT  1.520000  0.445000  1.690000 1.860000 ;
      RECT  1.520000  1.860000  3.530000 2.075000 ;
      RECT  1.520000  2.075000  1.805000 2.445000 ;
      RECT  1.975000  2.245000  2.355000 2.635000 ;
      RECT  2.145000  0.085000  2.475000 0.445000 ;
      RECT  2.250000  0.955000  2.695000 1.125000 ;
      RECT  2.250000  1.125000  2.420000 1.860000 ;
      RECT  2.875000  2.245000  3.870000 2.415000 ;
      RECT  3.050000  0.275000  3.875000 0.445000 ;
      RECT  3.335000  1.355000  3.555000 1.685000 ;
      RECT  3.335000  1.685000  3.530000 1.860000 ;
      RECT  3.700000  1.825000  4.685000 1.995000 ;
      RECT  3.700000  1.995000  3.870000 2.245000 ;
      RECT  3.705000  0.445000  3.875000 0.715000 ;
      RECT  3.705000  0.715000  4.685000 0.885000 ;
      RECT  4.090000  2.165000  4.260000 2.635000 ;
      RECT  4.095000  0.085000  4.295000 0.545000 ;
      RECT  4.515000  0.365000  4.865000 0.535000 ;
      RECT  4.515000  0.535000  4.685000 0.715000 ;
      RECT  4.515000  0.885000  4.685000 1.825000 ;
      RECT  4.515000  1.995000  4.685000 2.070000 ;
      RECT  4.515000  2.070000  4.800000 2.440000 ;
      RECT  4.855000  0.705000  5.485000 1.035000 ;
      RECT  4.855000  1.035000  5.145000 1.905000 ;
      RECT  4.995000  2.190000  6.215000 2.360000 ;
      RECT  5.085000  0.365000  5.875000 0.535000 ;
      RECT  5.335000  1.655000  5.825000 2.010000 ;
      RECT  5.705000  0.535000  5.875000 1.315000 ;
      RECT  5.705000  1.315000  6.555000 1.485000 ;
      RECT  5.995000  1.485000  6.555000 1.575000 ;
      RECT  5.995000  1.575000  6.215000 2.190000 ;
      RECT  6.095000  0.765000  6.945000 1.065000 ;
      RECT  6.095000  1.065000  6.265000 1.095000 ;
      RECT  6.175000  0.085000  6.545000 0.585000 ;
      RECT  6.385000  1.245000  6.555000 1.315000 ;
      RECT  6.385000  1.835000  6.555000 2.635000 ;
      RECT  6.725000  0.365000  7.235000 0.535000 ;
      RECT  6.725000  0.535000  6.945000 0.765000 ;
      RECT  6.725000  1.065000  6.945000 2.135000 ;
      RECT  6.725000  2.135000  7.025000 2.465000 ;
      RECT  7.115000  0.705000  7.715000 1.035000 ;
      RECT  7.115000  1.245000  7.355000 1.965000 ;
      RECT  7.250000  2.165000  8.285000 2.335000 ;
      RECT  7.515000  0.365000  8.155000 0.535000 ;
      RECT  7.525000  1.035000  7.715000 1.575000 ;
      RECT  7.525000  1.575000  7.895000 1.905000 ;
      RECT  7.935000  0.535000  8.155000 0.995000 ;
      RECT  7.935000  0.995000  9.045000 1.325000 ;
      RECT  7.935000  1.325000  8.285000 1.405000 ;
      RECT  8.115000  1.405000  8.285000 2.165000 ;
      RECT  8.380000  0.085000  8.800000 0.615000 ;
      RECT  8.485000  1.575000  9.400000 1.905000 ;
      RECT  8.515000  2.135000  8.820000 2.635000 ;
      RECT  9.070000  0.300000  9.400000 0.825000 ;
      RECT  9.110000  1.905000  9.400000 2.455000 ;
      RECT  9.215000  0.825000  9.400000 0.995000 ;
      RECT  9.215000  0.995000 10.050000 1.325000 ;
      RECT  9.215000  1.325000  9.400000 1.575000 ;
      RECT  9.620000  0.085000  9.790000 0.695000 ;
      RECT  9.620000  1.625000  9.790000 2.635000 ;
      RECT 10.610000  0.345000 10.860000 0.995000 ;
      RECT 10.610000  0.995000 11.440000 1.325000 ;
      RECT 10.610000  1.325000 10.860000 2.425000 ;
      RECT 11.065000  0.085000 11.395000 0.805000 ;
      RECT 11.090000  1.495000 11.395000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.695000  1.785000  0.865000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.115000  0.425000  1.285000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  0.765000  5.375000 0.935000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.615000  1.785000  5.785000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.175000  1.785000  7.345000 1.955000 ;
      RECT  7.185000  0.765000  7.355000 0.935000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.635000 1.755000 0.925000 1.800000 ;
      RECT 0.635000 1.800000 7.405000 1.940000 ;
      RECT 0.635000 1.940000 0.925000 1.985000 ;
      RECT 1.005000 0.395000 1.345000 0.440000 ;
      RECT 1.005000 0.440000 5.285000 0.580000 ;
      RECT 1.005000 0.580000 1.345000 0.625000 ;
      RECT 5.145000 0.580000 5.285000 0.735000 ;
      RECT 5.145000 0.735000 5.435000 0.780000 ;
      RECT 5.145000 0.780000 7.415000 0.920000 ;
      RECT 5.145000 0.920000 5.435000 0.965000 ;
      RECT 5.555000 1.755000 5.845000 1.800000 ;
      RECT 5.555000 1.940000 5.845000 1.985000 ;
      RECT 7.115000 1.755000 7.405000 1.800000 ;
      RECT 7.115000 1.940000 7.405000 1.985000 ;
      RECT 7.125000 0.735000 7.415000 0.780000 ;
      RECT 7.125000 0.920000 7.415000 0.965000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfxbp_1


MACRO sky130_fd_sc_hdll__bufbuf_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.360000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.480000 0.260000 3.860000 0.735000 ;
        RECT 3.480000 0.735000 7.240000 0.905000 ;
        RECT 3.480000 1.445000 7.240000 1.615000 ;
        RECT 3.480000 1.615000 3.860000 2.465000 ;
        RECT 4.420000 0.260000 4.800000 0.735000 ;
        RECT 4.420000 1.615000 4.800000 2.465000 ;
        RECT 5.360000 0.260000 5.740000 0.735000 ;
        RECT 5.360000 1.615000 5.740000 2.465000 ;
        RECT 6.300000 0.260000 6.680000 0.735000 ;
        RECT 6.300000 1.615000 6.680000 2.465000 ;
        RECT 6.860000 0.905000 7.240000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.095000  0.260000 0.425000 0.735000 ;
      RECT 0.095000  0.735000 0.830000 0.905000 ;
      RECT 0.095000  1.445000 0.830000 1.615000 ;
      RECT 0.095000  1.615000 0.425000 2.160000 ;
      RECT 0.645000  0.085000 0.815000 0.565000 ;
      RECT 0.645000  1.785000 0.815000 2.635000 ;
      RECT 0.660000  0.905000 0.830000 0.995000 ;
      RECT 0.660000  0.995000 1.140000 1.325000 ;
      RECT 0.660000  1.325000 0.830000 1.445000 ;
      RECT 1.050000  0.260000 1.480000 0.825000 ;
      RECT 1.050000  1.545000 1.480000 2.465000 ;
      RECT 1.310000  0.825000 1.480000 1.075000 ;
      RECT 1.310000  1.075000 2.920000 1.275000 ;
      RECT 1.310000  1.275000 1.480000 1.545000 ;
      RECT 1.650000  0.260000 1.980000 0.735000 ;
      RECT 1.650000  0.735000 3.310000 0.905000 ;
      RECT 1.650000  1.445000 3.310000 1.615000 ;
      RECT 1.650000  1.615000 1.980000 2.465000 ;
      RECT 2.200000  0.085000 2.370000 0.565000 ;
      RECT 2.200000  1.785000 2.370000 2.635000 ;
      RECT 2.540000  0.260000 2.920000 0.735000 ;
      RECT 2.540000  1.615000 2.920000 2.465000 ;
      RECT 3.140000  0.085000 3.310000 0.565000 ;
      RECT 3.140000  0.905000 3.310000 1.075000 ;
      RECT 3.140000  1.075000 5.910000 1.275000 ;
      RECT 3.140000  1.275000 3.310000 1.445000 ;
      RECT 3.140000  1.785000 3.310000 2.635000 ;
      RECT 4.080000  0.085000 4.250000 0.565000 ;
      RECT 4.080000  1.835000 4.250000 2.635000 ;
      RECT 5.020000  0.085000 5.190000 0.565000 ;
      RECT 5.020000  1.835000 5.190000 2.635000 ;
      RECT 5.960000  0.085000 6.130000 0.565000 ;
      RECT 5.960000  1.835000 6.130000 2.635000 ;
      RECT 6.900000  0.085000 7.070000 0.565000 ;
      RECT 6.900000  1.835000 7.070000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__bufbuf_8


MACRO sky130_fd_sc_hdll__bufbuf_16
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  13.34000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  4.016500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  5.735000 0.255000  6.035000 0.260000 ;
        RECT  5.735000 0.260000  6.115000 0.735000 ;
        RECT  5.735000 0.735000 13.220000 0.905000 ;
        RECT  5.735000 1.445000 13.220000 1.615000 ;
        RECT  5.735000 1.615000  6.115000 2.465000 ;
        RECT  6.675000 0.260000  7.055000 0.735000 ;
        RECT  6.675000 1.615000  7.055000 2.465000 ;
        RECT  6.805000 0.255000  6.975000 0.260000 ;
        RECT  7.615000 0.260000  7.995000 0.735000 ;
        RECT  7.615000 1.615000  7.995000 2.465000 ;
        RECT  7.745000 0.255000  7.915000 0.260000 ;
        RECT  8.555000 0.260000  8.935000 0.735000 ;
        RECT  8.555000 1.615000  8.935000 2.465000 ;
        RECT  9.495000 0.260000  9.875000 0.735000 ;
        RECT  9.495000 1.615000  9.875000 2.465000 ;
        RECT 10.435000 0.260000 10.815000 0.735000 ;
        RECT 10.435000 1.615000 10.815000 2.465000 ;
        RECT 11.375000 0.260000 11.755000 0.735000 ;
        RECT 11.375000 1.615000 11.755000 2.465000 ;
        RECT 12.315000 0.260000 12.695000 0.735000 ;
        RECT 12.315000 1.615000 12.695000 2.465000 ;
        RECT 12.920000 0.905000 13.220000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.340000 0.085000 ;
      RECT  0.000000  2.635000 13.340000 2.805000 ;
      RECT  0.175000  0.085000  0.345000 0.905000 ;
      RECT  0.175000  1.445000  0.345000 2.635000 ;
      RECT  0.515000  0.260000  0.895000 0.905000 ;
      RECT  0.515000  1.445000  0.895000 2.465000 ;
      RECT  0.660000  0.905000  0.895000 1.075000 ;
      RECT  0.660000  1.075000  2.355000 1.275000 ;
      RECT  0.660000  1.275000  0.895000 1.445000 ;
      RECT  1.085000  0.260000  1.415000 0.735000 ;
      RECT  1.085000  0.735000  2.745000 0.905000 ;
      RECT  1.085000  1.445000  2.745000 1.615000 ;
      RECT  1.085000  1.615000  1.415000 2.465000 ;
      RECT  1.635000  0.085000  1.805000 0.565000 ;
      RECT  1.635000  1.785000  1.805000 2.635000 ;
      RECT  1.975000  0.260000  2.355000 0.735000 ;
      RECT  1.975000  1.615000  2.355000 2.465000 ;
      RECT  2.575000  0.085000  2.745000 0.565000 ;
      RECT  2.575000  0.905000  2.745000 1.075000 ;
      RECT  2.575000  1.075000  5.135000 1.275000 ;
      RECT  2.575000  1.275000  2.745000 1.445000 ;
      RECT  2.575000  1.785000  2.745000 2.635000 ;
      RECT  2.915000  0.260000  3.295000 0.735000 ;
      RECT  2.915000  0.735000  5.565000 0.905000 ;
      RECT  2.915000  1.445000  5.565000 1.615000 ;
      RECT  2.915000  1.615000  3.295000 2.465000 ;
      RECT  3.515000  0.085000  3.685000 0.565000 ;
      RECT  3.515000  1.835000  3.685000 2.635000 ;
      RECT  3.855000  0.260000  4.235000 0.735000 ;
      RECT  3.855000  1.615000  4.235000 2.465000 ;
      RECT  4.455000  0.085000  4.625000 0.565000 ;
      RECT  4.455000  1.835000  4.625000 2.635000 ;
      RECT  4.795000  0.260000  5.175000 0.735000 ;
      RECT  4.795000  1.615000  5.175000 2.465000 ;
      RECT  5.390000  0.905000  5.565000 1.075000 ;
      RECT  5.390000  1.075000 12.700000 1.275000 ;
      RECT  5.390000  1.275000  5.565000 1.445000 ;
      RECT  5.395000  0.085000  5.565000 0.565000 ;
      RECT  5.395000  1.835000  5.565000 2.635000 ;
      RECT  6.335000  0.085000  6.505000 0.565000 ;
      RECT  6.335000  1.835000  6.505000 2.635000 ;
      RECT  7.275000  0.085000  7.445000 0.565000 ;
      RECT  7.275000  1.835000  7.445000 2.635000 ;
      RECT  8.215000  0.085000  8.385000 0.565000 ;
      RECT  8.215000  1.835000  8.385000 2.635000 ;
      RECT  9.155000  0.085000  9.325000 0.565000 ;
      RECT  9.155000  1.835000  9.325000 2.635000 ;
      RECT 10.095000  0.085000 10.265000 0.565000 ;
      RECT 10.095000  1.835000 10.265000 2.635000 ;
      RECT 11.035000  0.085000 11.205000 0.565000 ;
      RECT 11.035000  1.835000 11.205000 2.635000 ;
      RECT 11.975000  0.085000 12.145000 0.565000 ;
      RECT 11.975000  1.835000 12.145000 2.635000 ;
      RECT 12.915000  0.085000 13.085000 0.565000 ;
      RECT 12.915000  1.835000 13.085000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__bufbuf_16


MACRO sky130_fd_sc_hdll__probec_p_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.832500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.240000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -0.715000 1.030000 0.065000 1.350000 ;
      LAYER via3 ;
        RECT -0.625000 1.090000 -0.425000 1.290000 ;
        RECT -0.225000 1.090000 -0.025000 1.290000 ;
    END
  END X
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.615000  0.085000 0.895000 0.565000 ;
        RECT 1.505000  0.085000 1.805000 0.565000 ;
        RECT 2.475000  0.085000 2.745000 0.565000 ;
        RECT 3.415000  0.085000 3.685000 0.565000 ;
        RECT 4.355000  0.085000 4.625000 0.565000 ;
        RECT 5.295000  0.085000 5.545000 0.885000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
      LAYER via ;
        RECT 5.285000 -0.075000 5.435000 0.075000 ;
        RECT 5.605000 -0.075000 5.755000 0.075000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.595000 1.835000 0.865000 2.635000 ;
        RECT 1.535000 1.835000 1.805000 2.635000 ;
        RECT 2.475000 1.835000 2.745000 2.635000 ;
        RECT 3.415000 1.835000 3.685000 2.635000 ;
        RECT 4.355000 1.835000 4.625000 2.635000 ;
        RECT 5.295000 1.485000 5.595000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
      LAYER via ;
        RECT 5.285000 2.645000 5.435000 2.795000 ;
        RECT 5.605000 2.645000 5.755000 2.795000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 1.445000 1.595000 1.615000 ;
      RECT 0.095000 1.615000 0.425000 2.465000 ;
      RECT 0.145000 0.255000 0.445000 0.735000 ;
      RECT 0.145000 0.735000 1.595000 0.905000 ;
      RECT 1.035000 1.615000 1.365000 2.465000 ;
      RECT 1.065000 0.255000 1.335000 0.735000 ;
      RECT 1.420000 0.905000 1.595000 1.075000 ;
      RECT 1.420000 1.075000 4.045000 1.245000 ;
      RECT 1.420000 1.245000 1.595000 1.445000 ;
      RECT 1.975000 0.255000 2.305000 0.735000 ;
      RECT 1.975000 0.735000 5.125000 0.905000 ;
      RECT 1.975000 1.445000 5.125000 1.615000 ;
      RECT 1.975000 1.615000 2.305000 2.465000 ;
      RECT 2.915000 0.255000 3.245000 0.735000 ;
      RECT 2.915000 1.615000 3.245000 2.465000 ;
      RECT 3.855000 0.255000 4.185000 0.735000 ;
      RECT 3.855000 1.615000 4.185000 2.465000 ;
      RECT 4.290000 0.905000 5.125000 1.445000 ;
      RECT 4.795000 0.255000 5.125000 0.735000 ;
      RECT 4.795000 1.615000 5.125000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.305000  1.105000 4.475000 1.275000 ;
      RECT 4.665000  1.105000 4.835000 1.275000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 2.020000 1.060000 2.660000 1.120000 ;
      RECT 2.020000 1.120000 4.895000 1.260000 ;
      RECT 2.020000 1.260000 2.660000 1.320000 ;
      RECT 4.245000 1.075000 4.895000 1.120000 ;
      RECT 4.245000 1.260000 4.895000 1.305000 ;
    LAYER met2 ;
      RECT 1.890000  1.050000 2.660000 1.330000 ;
      RECT 5.135000 -0.140000 5.905000 0.140000 ;
      RECT 5.135000  2.580000 5.905000 2.860000 ;
    LAYER met3 ;
      RECT 1.885000  1.025000 2.665000 1.355000 ;
      RECT 5.130000 -0.165000 5.910000 0.165000 ;
      RECT 5.130000  2.555000 5.910000 2.885000 ;
    LAYER met4 ;
      RECT -1.140000  0.770000 0.040000 1.950000 ;
      RECT  1.460000  0.770000 2.640000 1.950000 ;
      RECT  4.930000 -0.895000 6.110000 0.285000 ;
      RECT  4.930000  2.435000 6.110000 3.615000 ;
    LAYER met5 ;
      RECT -1.260000  0.560000 2.760000 2.160000 ;
      RECT  1.160000 -1.105000 2.760000 0.560000 ;
      RECT  1.160000  2.160000 2.760000 3.825000 ;
      RECT  4.360000 -1.170000 6.675000 0.560000 ;
      RECT  4.360000  2.160000 6.675000 3.890000 ;
    LAYER via ;
      RECT 2.105000 1.115000 2.255000 1.265000 ;
      RECT 2.425000 1.115000 2.575000 1.265000 ;
    LAYER via2 ;
      RECT 1.975000  1.090000 2.175000 1.290000 ;
      RECT 2.375000  1.090000 2.575000 1.290000 ;
      RECT 5.220000 -0.100000 5.420000 0.100000 ;
      RECT 5.220000  2.620000 5.420000 2.820000 ;
      RECT 5.620000 -0.100000 5.820000 0.100000 ;
      RECT 5.620000  2.620000 5.820000 2.820000 ;
    LAYER via3 ;
      RECT 1.975000  1.090000 2.175000 1.290000 ;
      RECT 2.375000  1.090000 2.575000 1.290000 ;
      RECT 5.220000 -0.100000 5.420000 0.100000 ;
      RECT 5.220000  2.620000 5.420000 2.820000 ;
      RECT 5.620000 -0.100000 5.820000 0.100000 ;
      RECT 5.620000  2.620000 5.820000 2.820000 ;
    LAYER via4 ;
      RECT -0.950000  0.960000 -0.150000 1.760000 ;
      RECT  1.650000  0.960000  2.450000 1.760000 ;
      RECT  5.120000 -0.705000  5.920000 0.095000 ;
      RECT  5.120000  2.625000  5.920000 3.425000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__probec_p_8


MACRO sky130_fd_sc_hdll__a32oi_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 1.075000 3.255000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.720000 1.075000 4.575000 1.625000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.075000 6.320000 1.625000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.795000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.075000 0.875000 1.285000 ;
        RECT 0.145000 1.285000 0.325000 1.625000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.455000 2.195000 1.625000 ;
        RECT 0.565000 1.625000 0.895000 2.125000 ;
        RECT 1.455000 0.655000 3.245000 0.825000 ;
        RECT 1.585000 1.625000 1.755000 2.125000 ;
        RECT 1.965000 0.825000 2.195000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.095000  0.295000 0.425000 0.715000 ;
      RECT 0.095000  0.715000 1.285000 0.885000 ;
      RECT 0.175000  1.795000 0.345000 2.295000 ;
      RECT 0.175000  2.295000 2.225000 2.465000 ;
      RECT 0.645000  0.085000 0.815000 0.545000 ;
      RECT 1.035000  0.295000 2.305000 0.465000 ;
      RECT 1.035000  0.465000 1.285000 0.715000 ;
      RECT 1.115000  1.795000 1.285000 2.295000 ;
      RECT 2.055000  1.795000 6.265000 1.965000 ;
      RECT 2.055000  1.965000 2.225000 2.295000 ;
      RECT 2.445000  2.255000 3.165000 2.635000 ;
      RECT 2.495000  0.295000 4.605000 0.465000 ;
      RECT 3.415000  1.965000 3.585000 2.465000 ;
      RECT 3.755000  0.635000 5.800000 0.805000 ;
      RECT 3.770000  2.255000 4.525000 2.635000 ;
      RECT 4.695000  1.965000 4.865000 2.465000 ;
      RECT 4.865000  0.085000 5.250000 0.465000 ;
      RECT 5.125000  2.255000 5.845000 2.635000 ;
      RECT 5.420000  0.275000 5.800000 0.635000 ;
      RECT 6.095000  0.085000 6.265000 0.885000 ;
      RECT 6.095000  1.965000 6.265000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32oi_2


MACRO sky130_fd_sc_hdll__a32oi_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.50000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 1.075000 6.065000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.745000 1.075000 8.545000 1.300000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.145000 1.075000 11.035000 1.280000 ;
        RECT 10.755000 0.755000 11.035000 1.075000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.835000 0.995000 3.955000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.900000 1.305000 ;
        RECT 0.110000 1.305000 0.330000 1.965000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.575000 3.715000 1.745000 ;
        RECT 0.515000 1.745000 0.895000 2.085000 ;
        RECT 1.455000 1.745000 1.835000 2.085000 ;
        RECT 2.175000 0.990000 2.615000 1.575000 ;
        RECT 2.175000 1.745000 2.775000 2.085000 ;
        RECT 2.395000 0.635000 6.165000 0.805000 ;
        RECT 2.395000 0.805000 2.615000 0.990000 ;
        RECT 3.335000 1.745000 3.715000 2.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.500000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.500000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.500000 0.085000 ;
      RECT  0.000000  2.635000 11.500000 2.805000 ;
      RECT  0.095000  2.255000  4.105000 2.425000 ;
      RECT  0.175000  0.255000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  2.225000 0.805000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  1.115000  0.255000  1.285000 0.635000 ;
      RECT  1.455000  0.085000  1.835000 0.465000 ;
      RECT  2.055000  0.295000  4.185000 0.465000 ;
      RECT  2.055000  0.465000  2.225000 0.635000 ;
      RECT  3.935000  1.575000 10.975000 1.745000 ;
      RECT  3.935000  1.745000  4.105000 2.255000 ;
      RECT  4.295000  1.915000  4.675000 2.635000 ;
      RECT  4.425000  0.295000  8.655000 0.465000 ;
      RECT  4.895000  1.745000  5.065000 2.465000 ;
      RECT  5.320000  1.915000  6.040000 2.635000 ;
      RECT  6.290000  1.745000  6.460000 2.465000 ;
      RECT  6.865000  0.635000 10.505000 0.805000 ;
      RECT  6.865000  1.915000  7.245000 2.635000 ;
      RECT  7.465000  1.745000  7.635000 2.465000 ;
      RECT  7.805000  1.915000  8.185000 2.635000 ;
      RECT  8.405000  1.745000  8.575000 2.465000 ;
      RECT  8.845000  0.085000  9.175000 0.465000 ;
      RECT  9.265000  1.915000  9.645000 2.635000 ;
      RECT  9.395000  0.255000  9.565000 0.635000 ;
      RECT  9.735000  0.085000 10.115000 0.465000 ;
      RECT  9.865000  1.745000 10.035000 2.465000 ;
      RECT 10.205000  1.915000 10.585000 2.635000 ;
      RECT 10.335000  0.255000 10.505000 0.635000 ;
      RECT 10.685000  0.085000 11.075000 0.465000 ;
      RECT 10.805000  1.745000 10.975000 2.465000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32oi_4


MACRO sky130_fd_sc_hdll__a32oi_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 0.345000 1.695000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.415000 2.185000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.390000 1.015000 2.855000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.995000 1.235000 1.615000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.345000 1.325000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.634500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 1.265000 0.805000 ;
        RECT 0.515000 0.805000 0.775000 1.785000 ;
        RECT 0.515000 1.785000 0.915000 2.085000 ;
        RECT 0.965000 0.295000 1.265000 0.635000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.235000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.835000 0.345000 2.255000 ;
      RECT 0.085000  2.255000 1.445000 2.465000 ;
      RECT 0.110000  0.085000 0.440000 0.465000 ;
      RECT 1.195000  1.785000 2.385000 1.955000 ;
      RECT 1.195000  1.955000 1.445000 2.255000 ;
      RECT 1.705000  2.135000 1.955000 2.635000 ;
      RECT 2.215000  1.745000 2.385000 1.785000 ;
      RECT 2.215000  1.955000 2.385000 2.465000 ;
      RECT 2.555000  1.495000 2.945000 2.635000 ;
      RECT 2.570000  0.085000 2.960000 0.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32oi_1


MACRO sky130_fd_sc_hdll__o221a_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.820000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.305000 1.075000 3.955000 1.445000 ;
        RECT 3.305000 1.445000 5.225000 1.615000 ;
        RECT 4.975000 1.075000 5.535000 1.275000 ;
        RECT 4.975000 1.275000 5.225000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.125000 1.075000 4.755000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.730000 1.445000 ;
        RECT 1.065000 1.445000 3.045000 1.615000 ;
        RECT 2.665000 1.075000 3.045000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.950000 1.075000 2.495000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.440000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.735000 0.255000 6.115000 0.725000 ;
        RECT 5.735000 0.725000 7.055000 0.735000 ;
        RECT 5.735000 0.735000 7.710000 0.905000 ;
        RECT 5.865000 1.785000 6.500000 1.955000 ;
        RECT 5.865000 1.955000 6.075000 2.465000 ;
        RECT 6.330000 1.445000 7.710000 1.615000 ;
        RECT 6.330000 1.615000 6.500000 1.785000 ;
        RECT 6.675000 0.255000 7.055000 0.725000 ;
        RECT 6.765000 1.615000 7.015000 2.465000 ;
        RECT 7.365000 0.905000 7.710000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.255000 3.255000 0.475000 ;
      RECT 0.085000  0.475000 0.345000 0.895000 ;
      RECT 0.145000  1.455000 0.395000 2.635000 ;
      RECT 0.515000  0.645000 0.895000 0.865000 ;
      RECT 0.615000  0.865000 0.895000 1.785000 ;
      RECT 0.615000  1.785000 5.645000 1.955000 ;
      RECT 0.615000  1.955000 0.865000 2.465000 ;
      RECT 1.085000  2.125000 1.335000 2.635000 ;
      RECT 1.115000  0.475000 1.285000 0.905000 ;
      RECT 1.455000  0.645000 4.235000 0.725000 ;
      RECT 1.455000  0.725000 5.175000 0.905000 ;
      RECT 1.555000  2.125000 1.805000 2.295000 ;
      RECT 1.555000  2.295000 2.745000 2.465000 ;
      RECT 2.495000  2.125000 2.745000 2.295000 ;
      RECT 2.965000  2.125000 3.725000 2.635000 ;
      RECT 3.435000  0.085000 3.765000 0.465000 ;
      RECT 3.945000  2.125000 4.195000 2.295000 ;
      RECT 3.945000  2.295000 5.135000 2.465000 ;
      RECT 3.985000  0.255000 4.235000 0.645000 ;
      RECT 4.455000  0.085000 4.625000 0.555000 ;
      RECT 4.795000  0.255000 5.175000 0.725000 ;
      RECT 4.885000  2.125000 5.135000 2.295000 ;
      RECT 5.355000  2.125000 5.605000 2.635000 ;
      RECT 5.395000  0.085000 5.565000 0.905000 ;
      RECT 5.475000  1.445000 5.925000 1.615000 ;
      RECT 5.475000  1.615000 5.645000 1.785000 ;
      RECT 5.705000  1.075000 7.055000 1.275000 ;
      RECT 5.705000  1.275000 5.925000 1.445000 ;
      RECT 6.295000  2.125000 6.545000 2.635000 ;
      RECT 6.335000  0.085000 6.505000 0.555000 ;
      RECT 7.235000  1.795000 7.485000 2.635000 ;
      RECT 7.275000  0.085000 7.530000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221a_4


MACRO sky130_fd_sc_hdll__o221a_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815000 1.075000 3.145000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.980000 0.985000 2.615000 1.255000 ;
        RECT 1.980000 1.255000 2.315000 1.705000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.925000 0.985000 1.235000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.405000 0.985000 1.790000 1.705000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.415000 1.285000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.504500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.445000 0.265000 4.030000 0.825000 ;
        RECT 3.465000 1.875000 4.030000 2.465000 ;
        RECT 3.715000 0.825000 4.030000 1.875000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  1.455000 0.755000 1.495000 ;
      RECT 0.085000  1.495000 1.235000 1.720000 ;
      RECT 0.085000  1.720000 0.365000 2.465000 ;
      RECT 0.170000  0.255000 0.500000 0.645000 ;
      RECT 0.170000  0.645000 0.755000 0.825000 ;
      RECT 0.560000  2.085000 0.860000 2.635000 ;
      RECT 0.585000  0.825000 0.755000 1.455000 ;
      RECT 0.700000  0.305000 1.905000 0.475000 ;
      RECT 1.030000  1.720000 1.235000 1.875000 ;
      RECT 1.030000  1.875000 2.745000 2.045000 ;
      RECT 1.035000  0.645000 2.935000 0.815000 ;
      RECT 1.500000  2.045000 2.355000 2.465000 ;
      RECT 2.085000  0.085000 2.425000 0.475000 ;
      RECT 2.575000  1.455000 3.545000 1.625000 ;
      RECT 2.575000  1.625000 2.745000 1.875000 ;
      RECT 2.605000  0.270000 2.935000 0.645000 ;
      RECT 2.915000  1.795000 3.295000 2.635000 ;
      RECT 3.105000  0.085000 3.275000 0.640000 ;
      RECT 3.375000  0.995000 3.545000 1.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221a_1


MACRO sky130_fd_sc_hdll__o221a_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.835000 1.075000 3.325000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.235000 1.075000 2.615000 1.705000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 1.075000 1.330000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 1.075000 1.905000 1.705000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.345000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.545000 0.265000 3.925000 0.735000 ;
        RECT 3.545000 0.735000 4.490000 0.905000 ;
        RECT 3.545000 1.875000 4.490000 2.045000 ;
        RECT 3.545000 2.045000 3.845000 2.465000 ;
        RECT 4.180000 0.905000 4.490000 1.875000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.170000  0.255000 0.500000 0.635000 ;
      RECT 0.170000  0.635000 0.765000 0.805000 ;
      RECT 0.250000  1.495000 1.350000 1.670000 ;
      RECT 0.250000  1.670000 0.580000 2.465000 ;
      RECT 0.545000  0.805000 0.765000 1.445000 ;
      RECT 0.545000  1.445000 1.350000 1.495000 ;
      RECT 0.670000  0.295000 2.005000 0.465000 ;
      RECT 0.800000  1.850000 1.010000 2.635000 ;
      RECT 1.135000  0.645000 1.570000 0.735000 ;
      RECT 1.135000  0.735000 2.985000 0.905000 ;
      RECT 1.180000  1.670000 1.350000 1.875000 ;
      RECT 1.180000  1.875000 2.965000 2.045000 ;
      RECT 1.700000  2.045000 2.455000 2.465000 ;
      RECT 2.265000  0.085000 2.435000 0.555000 ;
      RECT 2.605000  0.270000 2.985000 0.735000 ;
      RECT 2.795000  1.455000 3.715000 1.625000 ;
      RECT 2.795000  1.625000 2.965000 1.875000 ;
      RECT 3.145000  1.795000 3.375000 2.635000 ;
      RECT 3.205000  0.085000 3.375000 0.905000 ;
      RECT 3.495000  1.075000 3.875000 1.285000 ;
      RECT 3.495000  1.285000 3.715000 1.455000 ;
      RECT 4.015000  2.215000 4.405000 2.635000 ;
      RECT 4.145000  0.085000 4.315000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221a_2


MACRO sky130_fd_sc_hdll__inputiso1n_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 2.085000 1.895000 2.415000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.325000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.472000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675000 0.415000 3.080000 0.760000 ;
        RECT 2.675000 1.495000 3.080000 2.465000 ;
        RECT 2.910000 0.760000 3.080000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.110000  0.265000 0.420000 0.735000 ;
      RECT 0.110000  0.735000 0.895000 0.905000 ;
      RECT 0.640000  0.085000 1.375000 0.565000 ;
      RECT 0.645000  0.905000 0.895000 0.995000 ;
      RECT 0.645000  0.995000 1.385000 1.325000 ;
      RECT 0.645000  1.325000 0.815000 1.885000 ;
      RECT 1.040000  1.495000 2.505000 1.665000 ;
      RECT 1.040000  1.665000 1.460000 1.915000 ;
      RECT 1.655000  0.305000 1.825000 0.655000 ;
      RECT 1.655000  0.655000 2.505000 0.825000 ;
      RECT 1.995000  0.085000 2.425000 0.485000 ;
      RECT 2.125000  1.835000 2.405000 2.635000 ;
      RECT 2.335000  0.825000 2.505000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inputiso1n_1


MACRO sky130_fd_sc_hdll__einvp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385000 0.975000 2.625000 1.955000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.236100 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.595000 1.725000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.488000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.980000 0.255000 2.625000 0.805000 ;
        RECT 1.980000 0.805000 2.155000 2.125000 ;
        RECT 1.980000 2.125000 2.625000 2.465000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 1.690000 0.825000 ;
      RECT 0.085000  1.895000 1.690000 2.065000 ;
      RECT 0.085000  2.065000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 1.500000 0.485000 ;
      RECT 0.515000  2.235000 1.740000 2.635000 ;
      RECT 0.765000  0.825000 1.690000 1.895000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvp_1


MACRO sky130_fd_sc_hdll__einvp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.245000 0.765000 3.535000 1.615000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.373200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.330000 1.615000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.645000 0.595000 3.075000 2.125000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.925000 0.825000 ;
      RECT 0.085000  1.785000 0.925000 1.955000 ;
      RECT 0.085000  1.955000 0.345000 2.465000 ;
      RECT 0.500000  0.825000 0.925000 0.995000 ;
      RECT 0.500000  0.995000 2.105000 1.325000 ;
      RECT 0.500000  1.325000 0.925000 1.785000 ;
      RECT 0.515000  0.085000 0.925000 0.485000 ;
      RECT 0.515000  2.125000 0.925000 2.635000 ;
      RECT 1.145000  0.255000 1.340000 0.655000 ;
      RECT 1.145000  0.655000 2.475000 0.825000 ;
      RECT 1.145000  1.555000 2.355000 1.725000 ;
      RECT 1.145000  1.725000 1.385000 2.465000 ;
      RECT 1.510000  0.085000 1.880000 0.485000 ;
      RECT 1.605000  1.895000 1.935000 2.635000 ;
      RECT 2.140000  0.255000 3.530000 0.425000 ;
      RECT 2.140000  0.425000 2.475000 0.655000 ;
      RECT 2.185000  1.725000 2.355000 2.295000 ;
      RECT 2.185000  2.295000 3.530000 2.465000 ;
      RECT 3.245000  0.425000 3.530000 0.595000 ;
      RECT 3.245000  1.785000 3.530000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvp_2


MACRO sky130_fd_sc_hdll__einvp_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.200000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.020000 1.020000 9.050000 1.275000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  1.057500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.330000 1.615000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.370000 0.635000 9.095000 0.850000 ;
        RECT 5.370000 0.850000 5.800000 1.445000 ;
        RECT 5.370000 1.445000 8.570000 1.615000 ;
        RECT 5.370000 1.615000 5.750000 2.125000 ;
        RECT 6.310000 1.615000 6.690000 2.125000 ;
        RECT 7.250000 1.615000 7.630000 2.125000 ;
        RECT 8.190000 1.615000 8.570000 2.125000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.745000 0.825000 ;
      RECT 0.085000  1.785000 0.925000 1.955000 ;
      RECT 0.085000  1.955000 0.345000 2.465000 ;
      RECT 0.500000  0.825000 0.745000 0.995000 ;
      RECT 0.500000  0.995000 5.200000 1.325000 ;
      RECT 0.500000  1.325000 0.925000 1.785000 ;
      RECT 0.515000  0.085000 0.895000 0.485000 ;
      RECT 0.515000  2.125000 0.925000 2.635000 ;
      RECT 1.135000  0.255000 1.305000 0.655000 ;
      RECT 1.135000  0.655000 5.200000 0.825000 ;
      RECT 1.175000  1.555000 5.200000 1.725000 ;
      RECT 1.175000  1.725000 1.385000 2.465000 ;
      RECT 1.475000  0.085000 1.855000 0.485000 ;
      RECT 1.605000  1.895000 1.935000 2.635000 ;
      RECT 2.075000  0.255000 2.245000 0.655000 ;
      RECT 2.155000  1.725000 2.325000 2.465000 ;
      RECT 2.415000  0.085000 2.795000 0.485000 ;
      RECT 2.545000  1.895000 2.875000 2.635000 ;
      RECT 3.015000  0.255000 3.185000 0.655000 ;
      RECT 3.095000  1.725000 3.265000 2.465000 ;
      RECT 3.355000  0.085000 3.735000 0.485000 ;
      RECT 3.485000  1.895000 3.815000 2.635000 ;
      RECT 3.955000  0.255000 4.125000 0.655000 ;
      RECT 4.035000  1.725000 4.205000 2.465000 ;
      RECT 4.295000  0.085000 4.685000 0.485000 ;
      RECT 4.425000  1.895000 4.755000 2.635000 ;
      RECT 4.855000  0.255000 9.095000 0.465000 ;
      RECT 4.855000  0.465000 5.200000 0.655000 ;
      RECT 4.975000  1.725000 5.200000 2.295000 ;
      RECT 4.975000  2.295000 9.095000 2.465000 ;
      RECT 5.970000  1.785000 6.140000 2.295000 ;
      RECT 6.910000  1.785000 7.080000 2.295000 ;
      RECT 7.850000  1.785000 8.020000 2.295000 ;
      RECT 8.790000  1.445000 9.095000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvp_8


MACRO sky130_fd_sc_hdll__einvp_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.520000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.210000 1.020000 5.410000 1.275000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.667500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.330000 1.615000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.490000 0.635000 5.410000 0.850000 ;
        RECT 3.490000 0.850000 4.030000 1.445000 ;
        RECT 3.490000 1.445000 4.810000 1.615000 ;
        RECT 3.490000 1.615000 3.870000 2.125000 ;
        RECT 4.430000 1.615000 4.810000 2.125000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.745000 0.825000 ;
      RECT 0.085000  1.785000 0.925000 1.955000 ;
      RECT 0.085000  1.955000 0.345000 2.465000 ;
      RECT 0.500000  0.825000 0.745000 0.995000 ;
      RECT 0.500000  0.995000 3.320000 1.325000 ;
      RECT 0.500000  1.325000 0.925000 1.785000 ;
      RECT 0.515000  0.085000 0.895000 0.485000 ;
      RECT 0.515000  2.125000 0.925000 2.635000 ;
      RECT 1.135000  0.255000 1.305000 0.655000 ;
      RECT 1.135000  0.655000 3.320000 0.825000 ;
      RECT 1.175000  1.555000 3.295000 1.725000 ;
      RECT 1.175000  1.725000 1.385000 2.465000 ;
      RECT 1.475000  0.085000 1.855000 0.485000 ;
      RECT 1.605000  1.895000 1.935000 2.635000 ;
      RECT 2.075000  0.255000 2.245000 0.655000 ;
      RECT 2.155000  1.725000 2.325000 2.465000 ;
      RECT 2.415000  0.085000 2.805000 0.485000 ;
      RECT 2.545000  1.895000 2.905000 2.635000 ;
      RECT 2.985000  0.255000 5.410000 0.465000 ;
      RECT 2.985000  0.465000 3.320000 0.655000 ;
      RECT 3.125000  1.725000 3.295000 2.295000 ;
      RECT 3.125000  2.295000 5.410000 2.465000 ;
      RECT 4.090000  1.785000 4.260000 2.295000 ;
      RECT 5.030000  1.445000 5.410000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvp_4


MACRO sky130_fd_sc_hdll__dlrtn_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.820000 BY  2.720000 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.955000 1.765000 1.300000 ;
    END
  END D
  PIN GATE_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.435000 1.625000 ;
    END
  END GATE_N
  PIN Q
    ANTENNADIFFAREA  0.931000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.815000 0.255000 6.195000 0.735000 ;
        RECT 5.815000 0.735000 7.085000 0.905000 ;
        RECT 5.815000 2.255000 6.145000 2.465000 ;
        RECT 5.845000 1.875000 6.145000 2.255000 ;
        RECT 5.895000 1.495000 7.085000 1.665000 ;
        RECT 5.895000 1.665000 6.145000 1.875000 ;
        RECT 6.405000 0.905000 7.085000 1.055000 ;
        RECT 6.405000 1.055000 7.265000 1.325000 ;
        RECT 6.405000 1.325000 7.085000 1.495000 ;
        RECT 6.755000 0.255000 7.085000 0.735000 ;
        RECT 6.755000 1.665000 7.085000 2.465000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.890000 0.995000 5.385000 1.325000 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  1.795000 0.895000 1.965000 ;
      RECT 0.085000  1.965000 0.395000 2.465000 ;
      RECT 0.225000  0.280000 0.395000 0.635000 ;
      RECT 0.225000  0.635000 0.775000 0.805000 ;
      RECT 0.565000  0.085000 0.895000 0.465000 ;
      RECT 0.565000  2.135000 0.895000 2.635000 ;
      RECT 0.605000  0.805000 0.775000 1.070000 ;
      RECT 0.605000  1.070000 0.895000 1.795000 ;
      RECT 1.065000  0.280000 1.235000 1.445000 ;
      RECT 1.065000  1.445000 1.335000 2.465000 ;
      RECT 1.555000  1.495000 2.115000 1.665000 ;
      RECT 1.555000  1.665000 1.885000 2.465000 ;
      RECT 1.660000  0.345000 1.855000 0.615000 ;
      RECT 1.660000  0.615000 2.115000 0.765000 ;
      RECT 1.660000  0.765000 2.535000 0.785000 ;
      RECT 1.945000  0.785000 2.535000 1.095000 ;
      RECT 1.945000  1.095000 2.115000 1.495000 ;
      RECT 2.025000  0.085000 2.355000 0.445000 ;
      RECT 2.055000  1.835000 2.325000 2.635000 ;
      RECT 2.445000  1.265000 2.955000 1.685000 ;
      RECT 2.780000  0.735000 3.295000 1.095000 ;
      RECT 3.020000  2.165000 3.850000 2.385000 ;
      RECT 3.040000  0.280000 3.660000 0.565000 ;
      RECT 3.125000  1.095000 3.295000 1.575000 ;
      RECT 3.125000  1.575000 3.510000 1.995000 ;
      RECT 3.490000  0.565000 3.660000 0.995000 ;
      RECT 3.490000  0.995000 4.380000 1.165000 ;
      RECT 3.680000  1.165000 4.380000 1.325000 ;
      RECT 3.680000  1.325000 3.850000 2.165000 ;
      RECT 3.870000  0.085000 4.200000 0.610000 ;
      RECT 4.020000  1.535000 5.725000 1.705000 ;
      RECT 4.020000  1.705000 5.175000 1.865000 ;
      RECT 4.020000  2.135000 4.705000 2.635000 ;
      RECT 4.455000  0.255000 4.785000 0.825000 ;
      RECT 4.550000  0.825000 4.720000 1.535000 ;
      RECT 4.875000  1.865000 5.175000 2.435000 ;
      RECT 5.315000  0.085000 5.645000 0.825000 ;
      RECT 5.345000  1.875000 5.675000 2.150000 ;
      RECT 5.345000  2.150000 5.645000 2.635000 ;
      RECT 5.555000  1.075000 6.235000 1.325000 ;
      RECT 5.555000  1.325000 5.725000 1.535000 ;
      RECT 6.315000  1.835000 6.585000 2.635000 ;
      RECT 6.375000  0.085000 6.585000 0.565000 ;
      RECT 7.255000  0.085000 7.465000 0.885000 ;
      RECT 7.255000  1.495000 7.510000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.635000  1.785000 0.805000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.095000  1.445000 1.265000 1.615000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.725000  1.445000 2.895000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.280000  1.785000 3.450000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 0.575000 1.755000 0.865000 1.800000 ;
      RECT 0.575000 1.800000 3.510000 1.940000 ;
      RECT 0.575000 1.940000 0.865000 1.985000 ;
      RECT 1.035000 1.415000 1.325000 1.460000 ;
      RECT 1.035000 1.460000 2.955000 1.600000 ;
      RECT 1.035000 1.600000 1.325000 1.645000 ;
      RECT 2.665000 1.415000 2.955000 1.460000 ;
      RECT 2.665000 1.600000 2.955000 1.645000 ;
      RECT 3.220000 1.755000 3.510000 1.800000 ;
      RECT 3.220000 1.940000 3.510000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtn_4


MACRO sky130_fd_sc_hdll__dlrtn_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.955000 1.765000 1.300000 ;
    END
  END D
  PIN GATE_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.435000 1.625000 ;
    END
  END GATE_N
  PIN Q
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.765000 0.255000 6.295000 0.495000 ;
        RECT 5.815000 2.255000 6.295000 2.465000 ;
        RECT 5.820000 0.495000 6.295000 0.885000 ;
        RECT 5.895000 1.495000 6.295000 2.255000 ;
        RECT 6.065000 0.885000 6.295000 1.495000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.890000 0.995000 5.385000 1.325000 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  1.795000 0.895000 1.965000 ;
      RECT 0.085000  1.965000 0.395000 2.465000 ;
      RECT 0.225000  0.280000 0.395000 0.635000 ;
      RECT 0.225000  0.635000 0.775000 0.805000 ;
      RECT 0.565000  0.085000 0.895000 0.465000 ;
      RECT 0.565000  2.135000 0.895000 2.635000 ;
      RECT 0.605000  0.805000 0.775000 1.070000 ;
      RECT 0.605000  1.070000 0.895000 1.795000 ;
      RECT 1.065000  0.280000 1.235000 1.445000 ;
      RECT 1.065000  1.445000 1.335000 2.465000 ;
      RECT 1.555000  1.495000 2.115000 1.665000 ;
      RECT 1.555000  1.665000 1.885000 2.465000 ;
      RECT 1.660000  0.345000 1.855000 0.615000 ;
      RECT 1.660000  0.615000 2.115000 0.765000 ;
      RECT 1.660000  0.765000 2.535000 0.785000 ;
      RECT 1.945000  0.785000 2.535000 1.095000 ;
      RECT 1.945000  1.095000 2.115000 1.495000 ;
      RECT 2.025000  0.085000 2.355000 0.445000 ;
      RECT 2.055000  1.835000 2.325000 2.635000 ;
      RECT 2.445000  1.265000 2.955000 1.685000 ;
      RECT 2.780000  0.735000 3.295000 1.095000 ;
      RECT 3.020000  2.165000 3.850000 2.385000 ;
      RECT 3.040000  0.280000 3.660000 0.565000 ;
      RECT 3.125000  1.095000 3.295000 1.575000 ;
      RECT 3.125000  1.575000 3.510000 1.995000 ;
      RECT 3.490000  0.565000 3.660000 0.995000 ;
      RECT 3.490000  0.995000 4.380000 1.165000 ;
      RECT 3.680000  1.165000 4.380000 1.325000 ;
      RECT 3.680000  1.325000 3.850000 2.165000 ;
      RECT 3.870000  0.085000 4.200000 0.610000 ;
      RECT 4.020000  1.535000 5.725000 1.705000 ;
      RECT 4.020000  1.705000 5.170000 1.865000 ;
      RECT 4.050000  2.135000 4.635000 2.635000 ;
      RECT 4.455000  0.255000 4.785000 0.825000 ;
      RECT 4.550000  0.825000 4.720000 1.535000 ;
      RECT 4.885000  1.865000 5.170000 2.465000 ;
      RECT 5.320000  0.085000 5.595000 0.625000 ;
      RECT 5.320000  0.625000 5.650000 0.825000 ;
      RECT 5.345000  1.885000 5.675000 2.150000 ;
      RECT 5.345000  2.150000 5.645000 2.635000 ;
      RECT 5.555000  1.055000 5.895000 1.325000 ;
      RECT 5.555000  1.325000 5.725000 1.535000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.635000  1.785000 0.805000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.095000  1.445000 1.265000 1.615000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.725000  1.445000 2.895000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.280000  1.785000 3.450000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.575000 1.755000 0.865000 1.800000 ;
      RECT 0.575000 1.800000 3.510000 1.940000 ;
      RECT 0.575000 1.940000 0.865000 1.985000 ;
      RECT 1.035000 1.415000 1.325000 1.460000 ;
      RECT 1.035000 1.460000 2.955000 1.600000 ;
      RECT 1.035000 1.600000 1.325000 1.645000 ;
      RECT 2.665000 1.415000 2.955000 1.460000 ;
      RECT 2.665000 1.600000 2.955000 1.645000 ;
      RECT 3.220000 1.755000 3.510000 1.800000 ;
      RECT 3.220000 1.940000 3.510000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtn_1


MACRO sky130_fd_sc_hdll__dlrtn_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.900000 BY  2.720000 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.955000 1.765000 1.300000 ;
    END
  END D
  PIN GATE_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.435000 1.625000 ;
    END
  END GATE_N
  PIN Q
    ANTENNADIFFAREA  0.465500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.815000 0.255000 6.205000 0.825000 ;
        RECT 5.815000 2.255000 6.205000 2.455000 ;
        RECT 5.895000 1.495000 6.205000 2.255000 ;
        RECT 6.035000 0.825000 6.205000 1.055000 ;
        RECT 6.035000 1.055000 6.435000 1.325000 ;
        RECT 6.035000 1.325000 6.205000 1.495000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.890000 0.995000 5.385000 1.325000 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.085000  1.795000 0.895000 1.965000 ;
      RECT 0.085000  1.965000 0.395000 2.465000 ;
      RECT 0.225000  0.280000 0.395000 0.635000 ;
      RECT 0.225000  0.635000 0.775000 0.805000 ;
      RECT 0.565000  0.085000 0.895000 0.465000 ;
      RECT 0.565000  2.135000 0.895000 2.635000 ;
      RECT 0.605000  0.805000 0.775000 1.070000 ;
      RECT 0.605000  1.070000 0.895000 1.795000 ;
      RECT 1.065000  0.280000 1.235000 1.445000 ;
      RECT 1.065000  1.445000 1.335000 2.465000 ;
      RECT 1.555000  1.495000 2.115000 1.665000 ;
      RECT 1.555000  1.665000 1.885000 2.465000 ;
      RECT 1.660000  0.345000 1.855000 0.615000 ;
      RECT 1.660000  0.615000 2.115000 0.765000 ;
      RECT 1.660000  0.765000 2.535000 0.785000 ;
      RECT 1.945000  0.785000 2.535000 1.095000 ;
      RECT 1.945000  1.095000 2.115000 1.495000 ;
      RECT 2.025000  0.085000 2.355000 0.445000 ;
      RECT 2.055000  1.835000 2.325000 2.635000 ;
      RECT 2.445000  1.265000 2.955000 1.685000 ;
      RECT 2.780000  0.735000 3.295000 1.095000 ;
      RECT 3.020000  2.165000 3.850000 2.385000 ;
      RECT 3.040000  0.280000 3.660000 0.565000 ;
      RECT 3.125000  1.095000 3.295000 1.575000 ;
      RECT 3.125000  1.575000 3.510000 1.995000 ;
      RECT 3.490000  0.565000 3.660000 0.995000 ;
      RECT 3.490000  0.995000 4.380000 1.165000 ;
      RECT 3.680000  1.165000 4.380000 1.325000 ;
      RECT 3.680000  1.325000 3.850000 2.165000 ;
      RECT 3.870000  0.085000 4.200000 0.610000 ;
      RECT 4.020000  1.535000 5.725000 1.705000 ;
      RECT 4.020000  1.705000 5.170000 1.865000 ;
      RECT 4.050000  2.135000 4.635000 2.635000 ;
      RECT 4.455000  0.255000 4.785000 0.825000 ;
      RECT 4.550000  0.825000 4.720000 1.535000 ;
      RECT 4.885000  1.865000 5.170000 2.465000 ;
      RECT 5.315000  0.085000 5.645000 0.825000 ;
      RECT 5.345000  1.885000 5.675000 2.150000 ;
      RECT 5.345000  2.150000 5.645000 2.635000 ;
      RECT 5.555000  0.995000 5.865000 1.325000 ;
      RECT 5.555000  1.325000 5.725000 1.535000 ;
      RECT 6.375000  0.085000 6.585000 0.885000 ;
      RECT 6.375000  1.495000 6.580000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.635000  1.785000 0.805000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.095000  1.445000 1.265000 1.615000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.725000  1.445000 2.895000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.280000  1.785000 3.450000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
    LAYER met1 ;
      RECT 0.575000 1.755000 0.865000 1.800000 ;
      RECT 0.575000 1.800000 3.510000 1.940000 ;
      RECT 0.575000 1.940000 0.865000 1.985000 ;
      RECT 1.035000 1.415000 1.325000 1.460000 ;
      RECT 1.035000 1.460000 2.955000 1.600000 ;
      RECT 1.035000 1.600000 1.325000 1.645000 ;
      RECT 2.665000 1.415000 2.955000 1.460000 ;
      RECT 2.665000 1.600000 2.955000 1.645000 ;
      RECT 3.220000 1.755000 3.510000 1.800000 ;
      RECT 3.220000 1.940000 3.510000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlrtn_2


MACRO sky130_fd_sc_hdll__o221ai_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.730000 1.075000 4.110000 1.445000 ;
        RECT 3.730000 1.445000 5.265000 1.615000 ;
        RECT 5.095000 1.075000 5.835000 1.275000 ;
        RECT 5.095000 1.275000 5.265000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.280000 1.075000 4.875000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.120000 1.075000 2.185000 1.445000 ;
        RECT 1.120000 1.445000 3.560000 1.615000 ;
        RECT 3.180000 1.075000 3.560000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.355000 1.075000 3.010000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.435000 1.275000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.078000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.520000 0.645000 0.900000 0.865000 ;
        RECT 0.610000 1.445000 0.900000 1.785000 ;
        RECT 0.610000 1.785000 4.750000 1.955000 ;
        RECT 0.610000 1.955000 0.860000 2.465000 ;
        RECT 0.655000 0.865000 0.900000 1.445000 ;
        RECT 2.540000 1.955000 2.790000 2.125000 ;
        RECT 4.500000 1.955000 4.750000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.100000  0.255000 1.370000 0.475000 ;
      RECT 0.100000  0.475000 0.350000 0.895000 ;
      RECT 0.140000  1.455000 0.390000 2.635000 ;
      RECT 1.080000  2.125000 1.850000 2.635000 ;
      RECT 1.120000  0.475000 1.370000 0.645000 ;
      RECT 1.120000  0.645000 3.300000 0.905000 ;
      RECT 1.560000  0.255000 3.850000 0.475000 ;
      RECT 2.070000  2.125000 2.320000 2.295000 ;
      RECT 2.070000  2.295000 3.260000 2.465000 ;
      RECT 3.010000  2.125000 3.260000 2.295000 ;
      RECT 3.480000  2.125000 3.810000 2.635000 ;
      RECT 3.520000  0.475000 3.850000 0.735000 ;
      RECT 3.520000  0.735000 5.730000 0.905000 ;
      RECT 4.030000  2.125000 4.280000 2.295000 ;
      RECT 4.030000  2.295000 5.220000 2.465000 ;
      RECT 4.070000  0.085000 4.240000 0.555000 ;
      RECT 4.410000  0.255000 4.790000 0.725000 ;
      RECT 4.410000  0.725000 5.730000 0.735000 ;
      RECT 4.970000  1.785000 5.220000 2.295000 ;
      RECT 5.010000  0.085000 5.180000 0.555000 ;
      RECT 5.350000  0.255000 5.730000 0.725000 ;
      RECT 5.485000  1.455000 5.690000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221ai_2


MACRO sky130_fd_sc_hdll__o221ai_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.065000 1.075000 3.575000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.075000 2.895000 1.245000 ;
        RECT 2.635000 1.245000 2.895000 1.445000 ;
        RECT 2.635000 1.445000 3.125000 1.615000 ;
        RECT 2.855000 1.615000 3.125000 2.405000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 0.995000 1.595000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.815000 0.995000 2.325000 1.325000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.465000 1.325000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.974500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.365000 0.345000 0.645000 ;
        RECT 0.085000 0.645000 0.845000 0.825000 ;
        RECT 0.085000 1.495000 2.465000 1.705000 ;
        RECT 0.085000 1.705000 0.365000 2.465000 ;
        RECT 0.675000 0.825000 0.845000 1.495000 ;
        RECT 1.900000 1.705000 2.465000 2.180000 ;
        RECT 1.900000 2.180000 2.505000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.515000  0.305000 2.065000 0.475000 ;
      RECT 0.600000  1.875000 1.580000 2.635000 ;
      RECT 1.250000  0.645000 2.560000 0.695000 ;
      RECT 1.250000  0.695000 3.575000 0.825000 ;
      RECT 2.285000  0.280000 2.560000 0.645000 ;
      RECT 2.445000  0.825000 3.575000 0.865000 ;
      RECT 2.845000  0.085000 3.015000 0.525000 ;
      RECT 3.185000  0.280000 3.575000 0.695000 ;
      RECT 3.315000  1.455000 3.575000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221ai_1


MACRO sky130_fd_sc_hdll__o221ai_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.58000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.565000 1.075000  6.945000 1.445000 ;
        RECT 6.565000 1.445000  9.320000 1.615000 ;
        RECT 9.005000 1.075000 10.135000 1.275000 ;
        RECT 9.005000 1.275000  9.320000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.125000 1.075000 8.735000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.560000 1.075000 4.925000 1.275000 ;
        RECT 4.735000 1.275000 4.925000 1.445000 ;
        RECT 4.735000 1.445000 6.395000 1.615000 ;
        RECT 6.015000 1.075000 6.395000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.095000 0.995000 5.835000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.900000 1.275000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.156000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.645000 2.325000 0.865000 ;
        RECT 0.625000 1.445000 4.565000 1.615000 ;
        RECT 0.625000 1.615000 0.875000 2.465000 ;
        RECT 1.565000 1.615000 2.325000 1.955000 ;
        RECT 1.565000 1.955000 1.815000 2.465000 ;
        RECT 2.120000 0.865000 2.325000 1.445000 ;
        RECT 4.345000 1.615000 4.565000 1.785000 ;
        RECT 4.345000 1.785000 8.565000 2.005000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.115000  0.255000  6.135000 0.475000 ;
      RECT  0.115000  0.475000  0.365000 0.895000 ;
      RECT  0.155000  1.485000  0.405000 2.635000 ;
      RECT  1.095000  1.825000  1.345000 2.635000 ;
      RECT  2.035000  2.125000  2.805000 2.635000 ;
      RECT  2.515000  0.645000  6.685000 0.735000 ;
      RECT  2.515000  0.735000 10.445000 0.820000 ;
      RECT  3.025000  1.785000  4.175000 1.955000 ;
      RECT  3.025000  1.955000  3.275000 2.465000 ;
      RECT  3.495000  2.125000  3.745000 2.635000 ;
      RECT  3.965000  1.955000  4.175000 2.265000 ;
      RECT  3.965000  2.265000  6.135000 2.465000 ;
      RECT  6.015000  0.820000 10.445000 0.905000 ;
      RECT  6.355000  0.255000  6.685000 0.645000 ;
      RECT  6.355000  2.175000  6.605000 2.635000 ;
      RECT  6.775000  2.265000  8.995000 2.465000 ;
      RECT  6.905000  0.085000  7.075000 0.555000 ;
      RECT  7.245000  0.255000  7.625000 0.725000 ;
      RECT  7.245000  0.725000  8.565000 0.735000 ;
      RECT  7.845000  0.085000  8.015000 0.555000 ;
      RECT  8.185000  0.255000  8.565000 0.725000 ;
      RECT  8.785000  0.085000  8.955000 0.555000 ;
      RECT  8.785000  1.785000  9.935000 1.955000 ;
      RECT  8.785000  1.955000  8.995000 2.265000 ;
      RECT  9.125000  0.255000  9.505000 0.725000 ;
      RECT  9.125000  0.725000 10.445000 0.735000 ;
      RECT  9.215000  2.125000  9.465000 2.635000 ;
      RECT  9.685000  1.445000  9.935000 1.785000 ;
      RECT  9.685000  1.955000  9.935000 2.465000 ;
      RECT  9.725000  0.085000  9.895000 0.555000 ;
      RECT 10.065000  0.255000 10.445000 0.725000 ;
      RECT 10.155000  1.445000 10.405000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221ai_4


MACRO sky130_fd_sc_hdll__and2_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 0.665000 1.325000 ;
        RECT 0.100000 1.325000 0.455000 1.685000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885000 1.075000 1.235000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.757200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.255000 2.155000 0.545000 ;
        RECT 1.730000 1.915000 2.155000 2.465000 ;
        RECT 1.860000 0.545000 2.155000 1.915000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.125000  0.355000 0.455000 0.715000 ;
      RECT 0.125000  0.715000 1.575000 0.905000 ;
      RECT 0.125000  1.965000 0.405000 2.635000 ;
      RECT 0.625000  1.575000 1.575000 1.745000 ;
      RECT 0.625000  1.745000 0.925000 2.295000 ;
      RECT 1.095000  1.915000 1.425000 2.635000 ;
      RECT 1.105000  0.085000 1.355000 0.545000 ;
      RECT 1.405000  0.905000 1.575000 0.995000 ;
      RECT 1.405000  0.995000 1.660000 1.325000 ;
      RECT 1.405000  1.325000 1.575000 1.575000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2_1


MACRO sky130_fd_sc_hdll__and2_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 0.995000 1.535000 1.295000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.615000 1.325000 ;
        RECT 0.435000 1.325000 0.615000 1.465000 ;
        RECT 0.435000 1.465000 1.885000 1.635000 ;
        RECT 1.705000 0.995000 1.965000 1.325000 ;
        RECT 1.705000 1.325000 1.885000 1.465000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.862000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.475000 0.255000 2.745000 0.715000 ;
        RECT 2.475000 0.715000 5.915000 0.885000 ;
        RECT 2.475000 1.445000 5.915000 1.615000 ;
        RECT 2.475000 1.615000 2.745000 2.465000 ;
        RECT 3.415000 0.255000 3.685000 0.715000 ;
        RECT 3.415000 1.615000 3.685000 2.465000 ;
        RECT 4.355000 0.255000 4.625000 0.715000 ;
        RECT 4.355000 1.615000 4.625000 2.465000 ;
        RECT 5.295000 0.255000 5.565000 0.715000 ;
        RECT 5.295000 1.615000 5.565000 2.465000 ;
        RECT 5.495000 0.885000 5.915000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.825000 ;
      RECT 0.095000  1.805000 0.395000 2.635000 ;
      RECT 0.565000  1.805000 2.305000 1.975000 ;
      RECT 0.565000  1.975000 0.865000 2.465000 ;
      RECT 1.015000  0.255000 1.345000 0.655000 ;
      RECT 1.015000  0.655000 2.305000 0.825000 ;
      RECT 1.035000  2.145000 1.365000 2.635000 ;
      RECT 1.535000  1.975000 1.805000 2.465000 ;
      RECT 1.940000  0.085000 2.270000 0.485000 ;
      RECT 1.975000  2.160000 2.305000 2.635000 ;
      RECT 2.135000  0.825000 2.305000 1.055000 ;
      RECT 2.135000  1.055000 5.325000 1.265000 ;
      RECT 2.135000  1.265000 2.305000 1.805000 ;
      RECT 2.915000  0.085000 3.245000 0.545000 ;
      RECT 2.915000  1.785000 3.245000 2.635000 ;
      RECT 3.855000  0.085000 4.185000 0.545000 ;
      RECT 3.855000  1.785000 4.185000 2.635000 ;
      RECT 4.795000  0.085000 5.125000 0.545000 ;
      RECT 4.795000  1.785000 5.125000 2.635000 ;
      RECT 5.735000  0.085000 6.065000 0.545000 ;
      RECT 5.735000  1.785000 6.065000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2_8


MACRO sky130_fd_sc_hdll__and2_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.075000 0.715000 1.325000 ;
        RECT 0.095000 1.325000 0.350000 1.765000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885000 1.075000 1.265000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.728500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595000 0.255000 2.205000 0.545000 ;
        RECT 1.745000 1.915000 2.205000 2.465000 ;
        RECT 1.935000 0.545000 2.205000 1.915000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.115000  0.355000 0.445000 0.715000 ;
      RECT 0.115000  0.715000 1.605000 0.905000 ;
      RECT 0.115000  1.965000 0.395000 2.635000 ;
      RECT 0.615000  1.575000 1.605000 1.745000 ;
      RECT 0.615000  1.745000 0.915000 2.295000 ;
      RECT 1.165000  1.915000 1.505000 2.635000 ;
      RECT 1.175000  0.085000 1.425000 0.545000 ;
      RECT 1.435000  0.905000 1.605000 0.995000 ;
      RECT 1.435000  0.995000 1.765000 1.325000 ;
      RECT 1.435000  1.325000 1.605000 1.575000 ;
      RECT 2.375000  0.085000 2.665000 0.885000 ;
      RECT 2.375000  1.495000 2.665000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2_2


MACRO sky130_fd_sc_hdll__and2_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.995000 0.435000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.995000 1.080000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.061500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.680000 0.515000 1.870000 0.615000 ;
        RECT 1.680000 0.615000 3.570000 0.845000 ;
        RECT 1.680000 1.535000 3.570000 1.760000 ;
        RECT 1.680000 1.760000 1.870000 2.465000 ;
        RECT 2.640000 0.255000 2.830000 0.615000 ;
        RECT 2.640000 1.760000 3.570000 1.765000 ;
        RECT 2.640000 1.765000 2.830000 2.465000 ;
        RECT 3.290000 0.845000 3.570000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  0.255000 0.425000 0.615000 ;
      RECT 0.095000  0.615000 1.460000 0.805000 ;
      RECT 0.095000  1.880000 0.425000 2.635000 ;
      RECT 0.655000  1.580000 1.460000 1.750000 ;
      RECT 0.655000  1.750000 0.835000 2.465000 ;
      RECT 1.055000  0.085000 1.385000 0.445000 ;
      RECT 1.090000  1.935000 1.420000 2.635000 ;
      RECT 1.250000  0.805000 1.460000 1.020000 ;
      RECT 1.250000  1.020000 2.935000 1.355000 ;
      RECT 1.250000  1.355000 1.460000 1.580000 ;
      RECT 2.040000  0.085000 2.420000 0.445000 ;
      RECT 2.040000  1.935000 2.420000 2.635000 ;
      RECT 3.000000  0.085000 3.380000 0.445000 ;
      RECT 3.000000  1.935000 3.380000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2_4


MACRO sky130_fd_sc_hdll__and2_6
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.520000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 0.995000 1.535000 1.295000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.615000 1.325000 ;
        RECT 0.435000 1.325000 0.615000 1.465000 ;
        RECT 0.435000 1.465000 1.885000 1.635000 ;
        RECT 1.705000 0.995000 1.965000 1.325000 ;
        RECT 1.705000 1.325000 1.885000 1.465000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.396500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.475000 0.255000 2.745000 0.715000 ;
        RECT 2.475000 0.715000 4.975000 0.885000 ;
        RECT 2.475000 1.445000 4.975000 1.615000 ;
        RECT 2.475000 1.615000 2.745000 2.465000 ;
        RECT 3.415000 0.255000 3.685000 0.715000 ;
        RECT 3.415000 1.615000 3.685000 2.465000 ;
        RECT 4.355000 0.255000 4.625000 0.715000 ;
        RECT 4.355000 1.615000 4.625000 2.465000 ;
        RECT 4.475000 0.885000 4.975000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.825000 ;
      RECT 0.095000  1.805000 0.395000 2.635000 ;
      RECT 0.565000  1.805000 2.305000 1.975000 ;
      RECT 0.565000  1.975000 0.865000 2.465000 ;
      RECT 1.015000  0.255000 1.345000 0.655000 ;
      RECT 1.015000  0.655000 2.305000 0.825000 ;
      RECT 1.035000  2.145000 1.365000 2.635000 ;
      RECT 1.535000  1.975000 1.805000 2.465000 ;
      RECT 1.940000  0.085000 2.270000 0.485000 ;
      RECT 1.975000  2.160000 2.305000 2.635000 ;
      RECT 2.135000  0.825000 2.305000 1.055000 ;
      RECT 2.135000  1.055000 4.305000 1.265000 ;
      RECT 2.135000  1.265000 2.305000 1.805000 ;
      RECT 2.915000  0.085000 3.245000 0.545000 ;
      RECT 2.915000  1.785000 3.245000 2.635000 ;
      RECT 3.855000  0.085000 4.185000 0.545000 ;
      RECT 3.855000  1.785000 4.185000 2.635000 ;
      RECT 4.795000  0.085000 5.125000 0.545000 ;
      RECT 4.795000  1.785000 5.125000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2_6


MACRO sky130_fd_sc_hdll__a21bo_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.885000 0.995000 3.085000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375000 0.995000 3.665000 1.615000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 0.995000 1.695000 1.325000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.547000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.715000 0.900000 0.885000 ;
        RECT 0.110000 0.885000 0.380000 1.835000 ;
        RECT 0.110000 1.835000 0.900000 2.005000 ;
        RECT 0.520000 0.315000 0.900000 0.715000 ;
        RECT 0.645000 2.005000 0.900000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.545000 ;
      RECT 0.090000  2.255000 0.425000 2.635000 ;
      RECT 0.620000  1.075000 0.950000 1.495000 ;
      RECT 0.620000  1.495000 1.385000 1.665000 ;
      RECT 1.070000  0.085000 1.400000 0.785000 ;
      RECT 1.140000  2.275000 1.470000 2.635000 ;
      RECT 1.215000  1.665000 1.385000 1.895000 ;
      RECT 1.215000  1.895000 2.375000 2.105000 ;
      RECT 1.555000  1.555000 2.035000 1.725000 ;
      RECT 1.605000  0.655000 2.035000 0.825000 ;
      RECT 1.865000  0.825000 2.035000 0.995000 ;
      RECT 1.865000  0.995000 2.325000 1.325000 ;
      RECT 1.865000  1.325000 2.035000 1.555000 ;
      RECT 2.125000  0.085000 2.455000 0.465000 ;
      RECT 2.125000  2.105000 2.375000 2.465000 ;
      RECT 2.205000  1.505000 2.715000 1.675000 ;
      RECT 2.205000  1.675000 2.375000 1.895000 ;
      RECT 2.495000  0.635000 2.940000 0.825000 ;
      RECT 2.495000  0.825000 2.715000 1.505000 ;
      RECT 2.545000  1.845000 3.875000 2.015000 ;
      RECT 2.545000  2.015000 2.925000 2.465000 ;
      RECT 3.155000  2.185000 3.325000 2.635000 ;
      RECT 3.495000  0.085000 3.875000 0.825000 ;
      RECT 3.495000  2.015000 3.875000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21bo_2


MACRO sky130_fd_sc_hdll__a21bo_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.960000 1.010000 5.375000 1.360000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.345000 1.010000 4.790000 1.275000 ;
        RECT 4.565000 1.275000 4.790000 1.595000 ;
        RECT 4.565000 1.595000 5.860000 1.765000 ;
        RECT 5.630000 1.055000 6.220000 1.290000 ;
        RECT 5.630000 1.290000 5.860000 1.595000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.470000 1.010000 0.850000 1.625000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  1.029000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.615000 2.510000 0.785000 ;
        RECT 1.050000 0.785000 1.540000 1.595000 ;
        RECT 1.050000 1.595000 2.580000 1.765000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.105000  0.255000 0.510000 0.840000 ;
      RECT 0.105000  0.840000 0.300000 1.795000 ;
      RECT 0.105000  1.795000 0.535000 1.935000 ;
      RECT 0.105000  1.935000 3.090000 2.105000 ;
      RECT 0.105000  2.105000 0.520000 2.465000 ;
      RECT 0.680000  0.085000 1.070000 0.445000 ;
      RECT 0.690000  2.275000 1.070000 2.635000 ;
      RECT 1.650000  0.085000 2.030000 0.445000 ;
      RECT 1.650000  2.275000 2.030000 2.635000 ;
      RECT 1.710000  0.995000 3.030000 1.185000 ;
      RECT 1.710000  1.185000 2.750000 1.325000 ;
      RECT 2.605000  2.275000 2.990000 2.635000 ;
      RECT 2.735000  0.085000 3.505000 0.445000 ;
      RECT 2.860000  0.615000 3.915000 0.670000 ;
      RECT 2.860000  0.670000 5.385000 0.785000 ;
      RECT 2.860000  0.785000 3.030000 0.995000 ;
      RECT 2.920000  1.355000 3.525000 1.525000 ;
      RECT 2.920000  1.525000 3.090000 1.935000 ;
      RECT 3.215000  0.995000 3.525000 1.355000 ;
      RECT 3.275000  1.695000 3.445000 2.210000 ;
      RECT 3.275000  2.210000 4.385000 2.380000 ;
      RECT 3.745000  0.255000 3.915000 0.615000 ;
      RECT 3.745000  0.785000 5.385000 0.840000 ;
      RECT 3.745000  0.840000 3.915000 1.805000 ;
      RECT 4.175000  0.085000 4.505000 0.445000 ;
      RECT 4.205000  1.445000 4.385000 1.935000 ;
      RECT 4.205000  1.935000 6.345000 2.105000 ;
      RECT 4.205000  2.105000 4.385000 2.210000 ;
      RECT 4.555000  2.275000 4.935000 2.635000 ;
      RECT 5.105000  0.405000 5.385000 0.670000 ;
      RECT 5.495000  2.275000 5.875000 2.635000 ;
      RECT 6.065000  0.085000 6.345000 0.885000 ;
      RECT 6.090000  1.460000 6.345000 1.935000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21bo_4


MACRO sky130_fd_sc_hdll__a21bo_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.900000 0.995000 2.275000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.995000 2.705000 1.615000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.325000 0.335000 1.665000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.628800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.715000 0.265000 3.995000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.105000  1.845000 0.965000 2.045000 ;
      RECT 0.105000  2.045000 0.345000 2.435000 ;
      RECT 0.515000  0.265000 0.795000 1.165000 ;
      RECT 0.515000  1.165000 0.965000 1.845000 ;
      RECT 0.515000  2.225000 0.915000 2.635000 ;
      RECT 1.045000  0.085000 1.290000 0.865000 ;
      RECT 1.135000  1.045000 1.730000 1.345000 ;
      RECT 1.135000  1.345000 1.465000 2.455000 ;
      RECT 1.460000  0.265000 1.940000 0.625000 ;
      RECT 1.460000  0.625000 3.545000 0.815000 ;
      RECT 1.460000  0.815000 1.730000 1.045000 ;
      RECT 1.685000  1.785000 2.810000 1.985000 ;
      RECT 1.685000  1.985000 1.865000 2.455000 ;
      RECT 2.035000  2.155000 2.415000 2.635000 ;
      RECT 2.620000  0.085000 3.350000 0.455000 ;
      RECT 2.640000  1.985000 2.810000 2.455000 ;
      RECT 3.075000  1.495000 3.360000 2.635000 ;
      RECT 3.285000  0.815000 3.545000 1.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21bo_1


MACRO sky130_fd_sc_hdll__nand4b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.660000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.180000 1.075000 5.040000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.240000 1.075000 7.110000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.665000 1.075000 9.505000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.736000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 0.635000 2.840000 0.905000 ;
        RECT 1.505000 1.445000 8.985000 1.665000 ;
        RECT 1.505000 1.665000 1.885000 2.465000 ;
        RECT 2.410000 0.905000 2.840000 1.445000 ;
        RECT 2.445000 1.665000 2.825000 2.465000 ;
        RECT 3.385000 1.665000 3.765000 2.465000 ;
        RECT 4.325000 1.665000 4.705000 2.465000 ;
        RECT 5.785000 1.665000 6.165000 2.465000 ;
        RECT 6.725000 1.665000 7.105000 2.465000 ;
        RECT 7.665000 1.665000 8.045000 2.465000 ;
        RECT 8.605000 1.665000 8.985000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 0.855000 0.905000 ;
      RECT 0.090000  1.495000 0.855000 1.665000 ;
      RECT 0.090000  1.665000 0.425000 2.465000 ;
      RECT 0.645000  0.085000 0.895000 0.545000 ;
      RECT 0.645000  1.835000 1.335000 2.635000 ;
      RECT 0.660000  0.905000 0.855000 1.075000 ;
      RECT 0.660000  1.075000 1.975000 1.275000 ;
      RECT 0.660000  1.275000 0.855000 1.495000 ;
      RECT 1.045000  1.495000 1.335000 1.835000 ;
      RECT 1.085000  0.255000 5.175000 0.465000 ;
      RECT 1.085000  0.465000 1.335000 0.905000 ;
      RECT 2.105000  1.835000 2.275000 2.635000 ;
      RECT 3.045000  1.835000 3.215000 2.635000 ;
      RECT 3.385000  0.635000 7.105000 0.905000 ;
      RECT 3.985000  1.835000 4.155000 2.635000 ;
      RECT 4.925000  1.835000 5.615000 2.635000 ;
      RECT 5.365000  0.255000 7.575000 0.465000 ;
      RECT 6.385000  1.835000 6.555000 2.635000 ;
      RECT 7.325000  0.465000 7.575000 0.735000 ;
      RECT 7.325000  0.735000 9.460000 0.905000 ;
      RECT 7.325000  1.835000 7.495000 2.635000 ;
      RECT 7.795000  0.085000 7.965000 0.545000 ;
      RECT 8.135000  0.255000 8.515000 0.735000 ;
      RECT 8.265000  1.835000 8.435000 2.635000 ;
      RECT 8.735000  0.085000 8.905000 0.545000 ;
      RECT 9.075000  0.255000 9.460000 0.735000 ;
      RECT 9.205000  1.445000 9.460000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4b_4


MACRO sky130_fd_sc_hdll__nand4b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.330000 1.615000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.160000 1.075000 3.350000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 1.075000 4.685000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.020000 1.075000 5.885000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.368000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 0.635000 1.885000 1.445000 ;
        RECT 1.505000 1.445000 5.265000 1.665000 ;
        RECT 1.505000 1.665000 1.885000 2.465000 ;
        RECT 2.445000 1.665000 2.825000 2.465000 ;
        RECT 3.855000 1.665000 4.235000 2.465000 ;
        RECT 4.885000 1.665000 5.265000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.090000  0.255000 0.345000 0.635000 ;
      RECT 0.090000  0.635000 0.720000 0.805000 ;
      RECT 0.090000  1.915000 0.720000 2.085000 ;
      RECT 0.090000  2.085000 0.345000 2.465000 ;
      RECT 0.500000  0.805000 0.720000 1.075000 ;
      RECT 0.500000  1.075000 1.335000 1.245000 ;
      RECT 0.500000  1.245000 0.720000 1.915000 ;
      RECT 0.515000  0.085000 0.895000 0.465000 ;
      RECT 0.515000  2.255000 1.335000 2.635000 ;
      RECT 1.085000  0.255000 2.275000 0.465000 ;
      RECT 1.085000  0.465000 1.335000 0.905000 ;
      RECT 1.085000  1.445000 1.335000 2.255000 ;
      RECT 2.105000  0.465000 2.275000 0.635000 ;
      RECT 2.105000  0.635000 3.295000 0.905000 ;
      RECT 2.105000  1.835000 2.275000 2.635000 ;
      RECT 2.445000  0.255000 4.285000 0.465000 ;
      RECT 3.045000  1.835000 3.685000 2.635000 ;
      RECT 3.485000  0.635000 4.805000 0.715000 ;
      RECT 3.485000  0.715000 5.790000 0.905000 ;
      RECT 4.455000  1.835000 4.715000 2.635000 ;
      RECT 4.505000  0.255000 4.765000 0.615000 ;
      RECT 4.505000  0.615000 4.805000 0.635000 ;
      RECT 5.065000  0.085000 5.235000 0.545000 ;
      RECT 5.455000  0.255000 5.790000 0.715000 ;
      RECT 5.485000  1.495000 5.880000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4b_2


MACRO sky130_fd_sc_hdll__nand4b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.820000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.930000 0.765000 2.225000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 0.960000 1.760000 1.325000 ;
        RECT 1.540000 0.765000 1.760000 0.960000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.995000 1.330000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.882500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.175000 1.495000 3.135000 1.665000 ;
        RECT 1.175000 1.665000 1.555000 2.465000 ;
        RECT 2.175000 1.665000 2.505000 2.465000 ;
        RECT 2.775000 0.255000 3.135000 0.835000 ;
        RECT 2.875000 0.835000 3.135000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.445000 0.470000 0.655000 ;
      RECT 0.085000  0.655000 1.370000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.595000 ;
      RECT 0.085000  1.595000 0.505000 1.925000 ;
      RECT 0.665000  0.085000 1.030000 0.485000 ;
      RECT 0.755000  1.495000 1.005000 2.635000 ;
      RECT 1.200000  0.425000 2.600000 0.595000 ;
      RECT 1.200000  0.595000 1.370000 0.655000 ;
      RECT 1.725000  1.835000 2.000000 2.635000 ;
      RECT 2.395000  0.595000 2.600000 0.995000 ;
      RECT 2.395000  0.995000 2.705000 1.325000 ;
      RECT 2.875000  1.835000 3.090000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4b_1


MACRO sky130_fd_sc_hdll__dlygate4sd3_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.605000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.190000 0.255000 3.595000 0.825000 ;
        RECT 3.190000 1.495000 3.595000 2.465000 ;
        RECT 3.325000 0.825000 3.595000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  1.785000 0.945000 2.005000 ;
      RECT 0.085000  2.005000 0.380000 2.465000 ;
      RECT 0.095000  0.255000 0.380000 0.715000 ;
      RECT 0.095000  0.715000 0.945000 0.885000 ;
      RECT 0.600000  0.085000 0.815000 0.545000 ;
      RECT 0.605000  2.175000 0.855000 2.635000 ;
      RECT 0.775000  0.885000 0.945000 0.995000 ;
      RECT 0.775000  0.995000 1.400000 1.325000 ;
      RECT 0.775000  1.325000 0.945000 1.785000 ;
      RECT 1.305000  0.255000 1.740000 0.545000 ;
      RECT 1.305000  2.175000 1.740000 2.465000 ;
      RECT 1.570000  0.545000 1.740000 1.075000 ;
      RECT 1.570000  1.075000 2.475000 1.275000 ;
      RECT 1.570000  1.275000 1.740000 2.175000 ;
      RECT 1.910000  0.510000 2.140000 0.735000 ;
      RECT 1.910000  0.735000 3.020000 0.905000 ;
      RECT 1.910000  1.575000 3.020000 1.745000 ;
      RECT 1.910000  1.745000 2.130000 2.080000 ;
      RECT 2.690000  0.085000 3.020000 0.565000 ;
      RECT 2.690000  1.915000 3.020000 2.635000 ;
      RECT 2.810000  0.905000 3.020000 0.995000 ;
      RECT 2.810000  0.995000 3.155000 1.325000 ;
      RECT 2.810000  1.325000 3.020000 1.575000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlygate4sd3_1


MACRO sky130_fd_sc_hdll__mux2_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.450000 0.995000 1.795000 1.615000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 0.995000 2.585000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.790000 1.325000 ;
        RECT 0.620000 0.635000 3.050000 0.805000 ;
        RECT 0.620000 0.805000 0.790000 0.995000 ;
        RECT 2.880000 0.805000 3.050000 0.995000 ;
        RECT 2.880000 0.995000 3.595000 1.325000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.215000 0.255000 4.385000 0.635000 ;
        RECT 4.215000 0.635000 5.880000 0.805000 ;
        RECT 4.215000 1.575000 5.880000 1.745000 ;
        RECT 4.215000 1.745000 4.385000 2.465000 ;
        RECT 5.155000 0.255000 5.325000 0.635000 ;
        RECT 5.155000 1.745000 5.325000 2.465000 ;
        RECT 5.650000 0.805000 5.880000 1.575000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.090000  0.295000 0.345000 0.625000 ;
      RECT 0.090000  0.625000 0.260000 1.495000 ;
      RECT 0.090000  1.495000 1.180000 1.665000 ;
      RECT 0.090000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.895000 0.465000 ;
      RECT 0.515000  1.835000 0.870000 2.635000 ;
      RECT 0.960000  0.995000 1.180000 1.495000 ;
      RECT 1.040000  1.935000 1.440000 2.275000 ;
      RECT 1.040000  2.275000 2.970000 2.445000 ;
      RECT 1.630000  1.935000 3.445000 2.105000 ;
      RECT 2.075000  0.295000 3.430000 0.465000 ;
      RECT 2.130000  1.595000 3.985000 1.765000 ;
      RECT 3.260000  0.465000 3.430000 0.655000 ;
      RECT 3.260000  0.655000 3.985000 0.825000 ;
      RECT 3.275000  2.105000 3.445000 2.465000 ;
      RECT 3.615000  0.085000 3.995000 0.465000 ;
      RECT 3.615000  2.255000 3.995000 2.635000 ;
      RECT 3.815000  0.825000 3.985000 1.075000 ;
      RECT 3.815000  1.075000 5.430000 1.245000 ;
      RECT 3.815000  1.245000 3.985000 1.595000 ;
      RECT 4.555000  0.085000 4.935000 0.465000 ;
      RECT 4.555000  1.915000 4.935000 2.635000 ;
      RECT 5.495000  0.085000 5.875000 0.465000 ;
      RECT 5.495000  1.915000 5.875000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_4


MACRO sky130_fd_sc_hdll__mux2_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.290000 0.255000 2.615000 1.415000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.815000 1.950000 1.615000 ;
        RECT 1.780000 1.615000 3.075000 1.785000 ;
        RECT 2.855000 0.255000 3.075000 1.615000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.277200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 0.995000 1.270000 1.325000 ;
        RECT 1.070000 1.325000 1.270000 2.295000 ;
        RECT 1.070000 2.295000 3.415000 2.465000 ;
        RECT 3.245000 1.440000 4.045000 1.630000 ;
        RECT 3.245000 1.630000 3.415000 2.295000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.255000 0.345000 1.495000 ;
        RECT 0.090000 1.495000 0.425000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.515000  0.085000 0.895000 0.485000 ;
      RECT 0.515000  0.655000 1.610000 0.825000 ;
      RECT 0.515000  0.825000 0.685000 1.325000 ;
      RECT 0.645000  1.495000 0.815000 2.635000 ;
      RECT 1.435000  0.255000 1.955000 0.620000 ;
      RECT 1.435000  0.620000 1.610000 0.655000 ;
      RECT 1.440000  0.825000 1.610000 1.955000 ;
      RECT 1.440000  1.955000 2.750000 2.125000 ;
      RECT 3.250000  0.085000 3.765000 0.620000 ;
      RECT 3.285000  0.895000 4.500000 1.065000 ;
      RECT 3.585000  1.875000 3.755000 2.635000 ;
      RECT 4.035000  0.290000 4.280000 0.895000 ;
      RECT 4.040000  1.875000 4.500000 2.285000 ;
      RECT 4.215000  1.065000 4.500000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_1


MACRO sky130_fd_sc_hdll__mux2_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.58000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.580000 0.645000 7.495000 0.815000 ;
        RECT 5.580000 0.815000 5.800000 1.325000 ;
        RECT 5.755000 0.425000 6.390000 0.645000 ;
        RECT 7.325000 0.815000 7.495000 0.995000 ;
        RECT 7.325000 0.995000 7.845000 1.165000 ;
        RECT 7.625000 1.165000 7.845000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.620000 1.075000 4.960000 1.120000 ;
        RECT 4.620000 1.120000 9.115000 1.260000 ;
        RECT 4.620000 1.260000 4.960000 1.305000 ;
        RECT 8.765000 1.075000 9.115000 1.120000 ;
        RECT 8.765000 1.260000 9.115000 1.305000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.110000 1.415000  6.400000 1.460000 ;
        RECT 6.110000 1.460000 10.035000 1.600000 ;
        RECT 6.110000 1.600000  6.400000 1.645000 ;
        RECT 9.745000 1.415000 10.035000 1.460000 ;
        RECT 9.745000 1.600000 10.035000 1.645000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.255000 0.815000 0.635000 ;
        RECT 0.605000 0.635000 3.635000 0.805000 ;
        RECT 0.605000 0.805000 0.865000 1.575000 ;
        RECT 0.605000 1.575000 3.635000 1.745000 ;
        RECT 0.605000 1.745000 0.815000 2.465000 ;
        RECT 1.585000 0.295000 1.755000 0.635000 ;
        RECT 1.585000 1.745000 1.755000 2.465000 ;
        RECT 2.525000 0.255000 2.695000 0.635000 ;
        RECT 2.525000 1.745000 2.695000 2.465000 ;
        RECT 3.465000 0.295000 3.635000 0.635000 ;
        RECT 3.465000 1.745000 3.635000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.090000  0.085000  0.425000 0.465000 ;
      RECT  0.090000  1.915000  0.425000 2.635000 ;
      RECT  0.985000  0.085000  1.365000 0.465000 ;
      RECT  0.985000  1.915000  1.365000 2.635000 ;
      RECT  1.085000  1.075000  3.975000 1.245000 ;
      RECT  1.925000  0.085000  2.305000 0.465000 ;
      RECT  1.925000  1.915000  2.305000 2.635000 ;
      RECT  2.865000  0.085000  3.245000 0.465000 ;
      RECT  2.865000  1.915000  3.245000 2.635000 ;
      RECT  3.805000  0.085000  4.185000 0.465000 ;
      RECT  3.805000  0.635000  5.340000 0.805000 ;
      RECT  3.805000  0.805000  3.975000 1.075000 ;
      RECT  3.805000  1.245000  3.975000 1.835000 ;
      RECT  3.805000  1.835000  8.975000 2.005000 ;
      RECT  3.805000  2.255000  4.185000 2.635000 ;
      RECT  4.145000  0.995000  4.365000 1.495000 ;
      RECT  4.145000  1.495000  6.585000 1.665000 ;
      RECT  4.355000  0.295000  5.525000 0.465000 ;
      RECT  4.630000  2.255000  6.405000 2.425000 ;
      RECT  4.690000  1.105000  4.925000 1.275000 ;
      RECT  4.705000  0.995000  4.925000 1.105000 ;
      RECT  4.705000  1.275000  4.925000 1.325000 ;
      RECT  5.170000  0.805000  5.340000 0.935000 ;
      RECT  6.170000  0.995000  6.585000 1.495000 ;
      RECT  6.660000  0.085000  6.990000 0.465000 ;
      RECT  6.675000  2.175000  6.845000 2.635000 ;
      RECT  6.895000  0.995000  7.115000 1.495000 ;
      RECT  6.895000  1.495000  9.635000 1.665000 ;
      RECT  7.030000  2.255000  9.445000 2.425000 ;
      RECT  7.175000  0.295000  8.565000 0.465000 ;
      RECT  7.715000  0.635000  8.370000 0.805000 ;
      RECT  8.150000  0.805000  8.370000 0.935000 ;
      RECT  8.885000  0.995000  9.170000 1.325000 ;
      RECT  9.415000  0.645000 10.385000 0.815000 ;
      RECT  9.415000  0.815000  9.635000 1.495000 ;
      RECT  9.415000  1.665000  9.635000 1.915000 ;
      RECT  9.415000  1.915000 10.385000 2.085000 ;
      RECT  9.665000  0.085000 10.045000 0.465000 ;
      RECT  9.665000  2.255000 10.045000 2.635000 ;
      RECT  9.805000  0.995000 10.235000 1.615000 ;
      RECT 10.215000  0.295000 10.385000 0.645000 ;
      RECT 10.215000  1.795000 10.385000 1.915000 ;
      RECT 10.215000  2.085000 10.385000 2.465000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.690000  1.105000  4.860000 1.275000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.170000  0.765000  5.340000 0.935000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.170000  1.445000  6.340000 1.615000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.150000  0.765000  8.320000 0.935000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  1.105000  9.055000 1.275000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  1.445000  9.975000 1.615000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 5.110000 0.735000 5.400000 0.780000 ;
      RECT 5.110000 0.780000 8.430000 0.920000 ;
      RECT 5.110000 0.920000 5.400000 0.965000 ;
      RECT 8.090000 0.735000 8.430000 0.780000 ;
      RECT 8.090000 0.920000 8.430000 0.965000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_8


MACRO sky130_fd_sc_hdll__mux2_12
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  16.56000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.105000 1.075000 9.455000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.075000 1.915000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.075000 4.275000 1.325000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  2.793000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.585000 0.255000 10.915000 0.725000 ;
        RECT 10.585000 0.725000 15.615000 0.905000 ;
        RECT 10.585000 1.495000 15.615000 1.665000 ;
        RECT 10.585000 1.665000 10.915000 2.465000 ;
        RECT 11.525000 0.255000 11.855000 0.725000 ;
        RECT 11.525000 1.665000 11.855000 2.465000 ;
        RECT 12.465000 0.255000 12.795000 0.725000 ;
        RECT 12.465000 1.665000 12.795000 2.465000 ;
        RECT 13.405000 0.255000 13.735000 0.725000 ;
        RECT 13.405000 1.665000 13.735000 2.465000 ;
        RECT 14.345000 0.255000 14.675000 0.725000 ;
        RECT 14.345000 1.665000 14.675000 2.465000 ;
        RECT 15.285000 0.255000 15.615000 0.725000 ;
        RECT 15.285000 0.905000 15.615000 1.495000 ;
        RECT 15.285000 1.665000 15.615000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 16.560000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 16.560000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.560000 0.085000 ;
      RECT  0.000000  2.635000 16.560000 2.805000 ;
      RECT  0.095000  0.255000  2.305000 0.425000 ;
      RECT  0.095000  0.425000  0.395000 2.295000 ;
      RECT  0.095000  2.295000  2.305000 2.465000 ;
      RECT  0.565000  0.595000  0.895000 0.725000 ;
      RECT  0.565000  0.725000  4.235000 0.905000 ;
      RECT  0.565000  1.495000  1.835000 1.665000 ;
      RECT  0.565000  1.665000  0.895000 2.125000 ;
      RECT  1.065000  0.425000  1.335000 0.545000 ;
      RECT  1.065000  1.835000  1.335000 2.295000 ;
      RECT  1.505000  0.595000  1.835000 0.725000 ;
      RECT  1.505000  1.665000  1.835000 2.125000 ;
      RECT  2.005000  0.425000  2.305000 0.550000 ;
      RECT  2.005000  1.495000  2.305000 2.295000 ;
      RECT  2.525000  0.085000  2.795000 0.550000 ;
      RECT  2.525000  1.495000  2.795000 2.635000 ;
      RECT  2.965000  0.255000  3.295000 0.725000 ;
      RECT  2.965000  1.495000  4.235000 1.665000 ;
      RECT  2.965000  1.665000  3.295000 2.465000 ;
      RECT  3.465000  0.085000  3.735000 0.545000 ;
      RECT  3.465000  1.835000  3.735000 2.635000 ;
      RECT  3.905000  0.255000  4.235000 0.725000 ;
      RECT  3.905000  1.665000  4.235000 2.465000 ;
      RECT  4.405000  0.085000  4.675000 0.905000 ;
      RECT  4.405000  1.495000  4.675000 2.635000 ;
      RECT  4.845000  0.255000  5.175000 1.075000 ;
      RECT  4.845000  1.075000  7.095000 1.325000 ;
      RECT  4.845000  1.325000  5.175000 2.465000 ;
      RECT  5.345000  0.085000  5.615000 0.905000 ;
      RECT  5.345000  1.495000  5.615000 2.635000 ;
      RECT  5.785000  0.255000  6.115000 0.725000 ;
      RECT  5.785000  0.725000  9.455000 0.905000 ;
      RECT  5.785000  1.495000  7.055000 1.665000 ;
      RECT  5.785000  1.665000  6.115000 2.465000 ;
      RECT  6.285000  0.085000  6.555000 0.545000 ;
      RECT  6.285000  1.835000  6.555000 2.635000 ;
      RECT  6.725000  0.255000  7.055000 0.725000 ;
      RECT  6.725000  1.665000  7.055000 2.465000 ;
      RECT  7.225000  0.085000  7.495000 0.550000 ;
      RECT  7.225000  1.495000  7.495000 2.635000 ;
      RECT  7.715000  0.255000  9.925000 0.425000 ;
      RECT  7.715000  0.425000  8.015000 0.550000 ;
      RECT  7.715000  1.495000  8.015000 2.295000 ;
      RECT  7.715000  2.295000  9.925000 2.465000 ;
      RECT  8.185000  0.595000  8.515000 0.725000 ;
      RECT  8.185000  1.495000  9.455000 1.665000 ;
      RECT  8.185000  1.665000  8.515000 2.125000 ;
      RECT  8.685000  0.425000  8.955000 0.545000 ;
      RECT  8.685000  1.835000  8.955000 2.295000 ;
      RECT  9.125000  0.595000  9.455000 0.725000 ;
      RECT  9.125000  1.665000  9.455000 2.125000 ;
      RECT  9.625000  0.425000  9.925000 1.075000 ;
      RECT  9.625000  1.075000 14.825000 1.325000 ;
      RECT  9.625000  1.325000  9.925000 2.295000 ;
      RECT 10.145000  0.085000 10.415000 0.905000 ;
      RECT 10.145000  1.495000 10.415000 2.635000 ;
      RECT 11.085000  0.085000 11.355000 0.545000 ;
      RECT 11.085000  1.835000 11.355000 2.635000 ;
      RECT 12.025000  0.085000 12.295000 0.545000 ;
      RECT 12.025000  1.835000 12.295000 2.635000 ;
      RECT 12.965000  0.085000 13.235000 0.545000 ;
      RECT 12.965000  1.835000 13.235000 2.635000 ;
      RECT 13.905000  0.085000 14.175000 0.550000 ;
      RECT 13.905000  1.835000 14.175000 2.635000 ;
      RECT 14.845000  0.085000 15.115000 0.545000 ;
      RECT 14.845000  1.835000 15.115000 2.635000 ;
      RECT 15.785000  0.085000 16.055000 0.905000 ;
      RECT 15.785000  1.495000 16.055000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.175000  0.425000  0.345000 0.595000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.645000  1.785000  0.815000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.585000  1.785000  1.755000 1.955000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.045000  2.125000  3.215000 2.295000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  3.985000  2.125000  4.155000 2.295000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.865000  1.785000  6.035000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.805000  1.785000  6.975000 1.955000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.265000  1.785000  8.435000 1.955000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.205000  1.785000  9.375000 1.955000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.675000  0.425000  9.845000 0.595000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
    LAYER met1 ;
      RECT 0.115000 0.395000 0.405000 0.440000 ;
      RECT 0.115000 0.440000 9.905000 0.580000 ;
      RECT 0.115000 0.580000 0.405000 0.625000 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 7.035000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 1.525000 1.755000 1.815000 1.800000 ;
      RECT 1.525000 1.940000 1.815000 1.985000 ;
      RECT 2.985000 2.095000 3.275000 2.140000 ;
      RECT 2.985000 2.140000 7.660000 2.280000 ;
      RECT 2.985000 2.280000 3.275000 2.325000 ;
      RECT 3.925000 2.095000 4.215000 2.140000 ;
      RECT 3.925000 2.280000 4.215000 2.325000 ;
      RECT 5.805000 1.755000 6.095000 1.800000 ;
      RECT 5.805000 1.940000 6.095000 1.985000 ;
      RECT 6.745000 1.755000 7.035000 1.800000 ;
      RECT 6.745000 1.940000 7.035000 1.985000 ;
      RECT 7.520000 1.800000 9.435000 1.940000 ;
      RECT 7.520000 1.940000 7.660000 2.140000 ;
      RECT 8.205000 1.755000 8.495000 1.800000 ;
      RECT 8.205000 1.940000 8.495000 1.985000 ;
      RECT 9.145000 1.755000 9.435000 1.800000 ;
      RECT 9.145000 1.940000 9.435000 1.985000 ;
      RECT 9.615000 0.395000 9.905000 0.440000 ;
      RECT 9.615000 0.580000 9.905000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_12


MACRO sky130_fd_sc_hdll__mux2_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.920000 0.765000 2.295000 1.280000 ;
        RECT 1.920000 1.280000 3.075000 1.325000 ;
        RECT 2.125000 1.325000 3.075000 1.410000 ;
        RECT 2.135000 1.410000 3.075000 1.625000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.530000 0.775000 3.075000 1.105000 ;
        RECT 2.870000 0.420000 3.075000 0.775000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.355000 0.755000 3.545000 1.625000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.800000 1.595000 ;
        RECT 0.515000 1.595000 0.875000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.885000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.970000  0.995000 1.265000 1.325000 ;
      RECT 0.985000  0.085000 1.365000 0.465000 ;
      RECT 1.095000  0.635000 1.705000 0.805000 ;
      RECT 1.095000  0.805000 1.265000 0.995000 ;
      RECT 1.095000  1.325000 1.265000 1.835000 ;
      RECT 1.095000  1.835000 1.625000 2.005000 ;
      RECT 1.115000  2.175000 1.285000 2.635000 ;
      RECT 1.435000  0.995000 1.655000 1.495000 ;
      RECT 1.435000  1.495000 1.965000 1.665000 ;
      RECT 1.455000  2.005000 1.625000 2.255000 ;
      RECT 1.455000  2.255000 2.860000 2.425000 ;
      RECT 1.535000  0.265000 2.250000 0.595000 ;
      RECT 1.535000  0.595000 1.705000 0.635000 ;
      RECT 1.795000  1.665000 1.965000 1.835000 ;
      RECT 1.795000  1.835000 4.235000 2.005000 ;
      RECT 3.460000  2.175000 3.680000 2.635000 ;
      RECT 3.485000  0.085000 3.685000 0.585000 ;
      RECT 3.850000  2.005000 4.235000 2.465000 ;
      RECT 3.985000  0.255000 4.235000 1.835000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_2


MACRO sky130_fd_sc_hdll__mux2_16
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  18.40000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.105000 1.075000 9.455000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.075000 1.915000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.075000 4.275000 1.325000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  3.724000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.585000 0.255000 10.915000 0.725000 ;
        RECT 10.585000 0.725000 17.495000 0.905000 ;
        RECT 10.585000 1.495000 17.495000 1.665000 ;
        RECT 10.585000 1.665000 10.915000 2.465000 ;
        RECT 11.525000 0.255000 11.855000 0.725000 ;
        RECT 11.525000 1.665000 11.855000 2.465000 ;
        RECT 12.465000 0.255000 12.795000 0.725000 ;
        RECT 12.465000 1.665000 12.795000 2.465000 ;
        RECT 13.405000 0.255000 13.735000 0.725000 ;
        RECT 13.405000 1.665000 13.735000 2.465000 ;
        RECT 14.345000 0.255000 14.675000 0.725000 ;
        RECT 14.345000 1.665000 14.675000 2.465000 ;
        RECT 15.285000 0.255000 15.615000 0.725000 ;
        RECT 15.285000 1.665000 15.615000 2.465000 ;
        RECT 16.225000 0.255000 16.555000 0.725000 ;
        RECT 16.225000 1.665000 16.555000 2.465000 ;
        RECT 17.085000 0.905000 17.495000 1.495000 ;
        RECT 17.165000 0.255000 17.495000 0.725000 ;
        RECT 17.165000 1.665000 17.495000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 18.400000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 18.400000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 18.400000 0.085000 ;
      RECT  0.000000  2.635000 18.400000 2.805000 ;
      RECT  0.095000  0.255000  2.305000 0.425000 ;
      RECT  0.095000  0.425000  0.395000 2.295000 ;
      RECT  0.095000  2.295000  2.305000 2.465000 ;
      RECT  0.565000  0.595000  0.895000 0.725000 ;
      RECT  0.565000  0.725000  4.235000 0.905000 ;
      RECT  0.565000  1.495000  1.835000 1.665000 ;
      RECT  0.565000  1.665000  0.895000 2.125000 ;
      RECT  1.065000  0.425000  1.335000 0.545000 ;
      RECT  1.065000  1.835000  1.335000 2.295000 ;
      RECT  1.505000  0.595000  1.835000 0.725000 ;
      RECT  1.505000  1.665000  1.835000 2.125000 ;
      RECT  2.005000  0.425000  2.305000 0.550000 ;
      RECT  2.005000  1.495000  2.305000 2.295000 ;
      RECT  2.525000  0.085000  2.795000 0.550000 ;
      RECT  2.525000  1.495000  2.795000 2.635000 ;
      RECT  2.965000  0.255000  3.295000 0.725000 ;
      RECT  2.965000  1.495000  4.235000 1.665000 ;
      RECT  2.965000  1.665000  3.295000 2.465000 ;
      RECT  3.465000  0.085000  3.735000 0.545000 ;
      RECT  3.465000  1.835000  3.735000 2.635000 ;
      RECT  3.905000  0.255000  4.235000 0.725000 ;
      RECT  3.905000  1.665000  4.235000 2.465000 ;
      RECT  4.405000  0.085000  4.675000 0.905000 ;
      RECT  4.405000  1.495000  4.675000 2.635000 ;
      RECT  4.845000  0.255000  5.175000 1.075000 ;
      RECT  4.845000  1.075000  7.095000 1.325000 ;
      RECT  4.845000  1.325000  5.175000 2.465000 ;
      RECT  5.345000  0.085000  5.615000 0.905000 ;
      RECT  5.345000  1.495000  5.615000 2.635000 ;
      RECT  5.785000  0.255000  6.115000 0.725000 ;
      RECT  5.785000  0.725000  9.455000 0.905000 ;
      RECT  5.785000  1.495000  7.055000 1.665000 ;
      RECT  5.785000  1.665000  6.115000 2.465000 ;
      RECT  6.285000  0.085000  6.555000 0.545000 ;
      RECT  6.285000  1.835000  6.555000 2.635000 ;
      RECT  6.725000  0.255000  7.055000 0.725000 ;
      RECT  6.725000  1.665000  7.055000 2.465000 ;
      RECT  7.225000  0.085000  7.495000 0.550000 ;
      RECT  7.225000  1.495000  7.495000 2.635000 ;
      RECT  7.715000  0.255000  9.925000 0.425000 ;
      RECT  7.715000  0.425000  8.015000 0.550000 ;
      RECT  7.715000  1.495000  8.015000 2.295000 ;
      RECT  7.715000  2.295000  9.925000 2.465000 ;
      RECT  8.185000  0.595000  8.515000 0.725000 ;
      RECT  8.185000  1.495000  9.455000 1.665000 ;
      RECT  8.185000  1.665000  8.515000 2.125000 ;
      RECT  8.685000  0.425000  8.955000 0.545000 ;
      RECT  8.685000  1.835000  8.955000 2.295000 ;
      RECT  9.125000  0.595000  9.455000 0.725000 ;
      RECT  9.125000  1.665000  9.455000 2.125000 ;
      RECT  9.625000  0.425000  9.925000 1.075000 ;
      RECT  9.625000  1.075000 16.865000 1.325000 ;
      RECT  9.625000  1.325000  9.925000 2.295000 ;
      RECT 10.145000  0.085000 10.415000 0.905000 ;
      RECT 10.145000  1.495000 10.415000 2.635000 ;
      RECT 11.085000  0.085000 11.355000 0.545000 ;
      RECT 11.085000  1.835000 11.355000 2.635000 ;
      RECT 12.025000  0.085000 12.295000 0.545000 ;
      RECT 12.025000  1.835000 12.295000 2.635000 ;
      RECT 12.965000  0.085000 13.235000 0.545000 ;
      RECT 12.965000  1.835000 13.235000 2.635000 ;
      RECT 13.905000  0.085000 14.175000 0.550000 ;
      RECT 13.905000  1.835000 14.175000 2.635000 ;
      RECT 14.845000  0.085000 15.115000 0.545000 ;
      RECT 14.845000  1.835000 15.115000 2.635000 ;
      RECT 15.785000  0.085000 16.055000 0.545000 ;
      RECT 15.785000  1.835000 16.055000 2.635000 ;
      RECT 16.725000  0.085000 16.995000 0.545000 ;
      RECT 16.725000  1.835000 16.995000 2.635000 ;
      RECT 17.665000  0.085000 17.935000 0.905000 ;
      RECT 17.665000  1.495000 17.935000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.175000  0.425000  0.345000 0.595000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.645000  1.785000  0.815000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.585000  1.785000  1.755000 1.955000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.045000  2.125000  3.215000 2.295000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  3.985000  2.125000  4.155000 2.295000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.865000  1.785000  6.035000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.805000  1.785000  6.975000 1.955000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.265000  1.785000  8.435000 1.955000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.205000  1.785000  9.375000 1.955000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.675000  0.425000  9.845000 0.595000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
      RECT 17.165000 -0.085000 17.335000 0.085000 ;
      RECT 17.165000  2.635000 17.335000 2.805000 ;
      RECT 17.625000 -0.085000 17.795000 0.085000 ;
      RECT 17.625000  2.635000 17.795000 2.805000 ;
      RECT 18.085000 -0.085000 18.255000 0.085000 ;
      RECT 18.085000  2.635000 18.255000 2.805000 ;
    LAYER met1 ;
      RECT 0.115000 0.395000 0.405000 0.440000 ;
      RECT 0.115000 0.440000 9.905000 0.580000 ;
      RECT 0.115000 0.580000 0.405000 0.625000 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 7.035000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 1.525000 1.755000 1.815000 1.800000 ;
      RECT 1.525000 1.940000 1.815000 1.985000 ;
      RECT 2.985000 2.095000 3.275000 2.140000 ;
      RECT 2.985000 2.140000 7.660000 2.280000 ;
      RECT 2.985000 2.280000 3.275000 2.325000 ;
      RECT 3.925000 2.095000 4.215000 2.140000 ;
      RECT 3.925000 2.280000 4.215000 2.325000 ;
      RECT 5.805000 1.755000 6.095000 1.800000 ;
      RECT 5.805000 1.940000 6.095000 1.985000 ;
      RECT 6.745000 1.755000 7.035000 1.800000 ;
      RECT 6.745000 1.940000 7.035000 1.985000 ;
      RECT 7.520000 1.800000 9.435000 1.940000 ;
      RECT 7.520000 1.940000 7.660000 2.140000 ;
      RECT 8.205000 1.755000 8.495000 1.800000 ;
      RECT 8.205000 1.940000 8.495000 1.985000 ;
      RECT 9.145000 1.755000 9.435000 1.800000 ;
      RECT 9.145000 1.940000 9.435000 1.985000 ;
      RECT 9.615000 0.395000 9.905000 0.440000 ;
      RECT 9.615000 0.580000 9.905000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_16


MACRO sky130_fd_sc_hdll__a2bb2o_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.820000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.615000 1.075000 4.005000 1.325000 ;
        RECT 3.775000 1.325000 4.005000 1.445000 ;
        RECT 3.775000 1.445000 5.465000 1.615000 ;
        RECT 5.085000 1.075000 5.465000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.205000 1.075000 4.915000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.625000 1.445000 ;
        RECT 0.085000 1.445000 1.835000 1.615000 ;
        RECT 1.665000 1.075000 2.095000 1.245000 ;
        RECT 1.665000 1.245000 1.835000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 1.075000 1.445000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.735000 0.275000 6.115000 0.725000 ;
        RECT 5.735000 0.725000 7.675000 0.905000 ;
        RECT 5.825000 1.785000 7.015000 1.955000 ;
        RECT 5.825000 1.955000 6.075000 2.465000 ;
        RECT 6.675000 0.275000 7.055000 0.725000 ;
        RECT 6.765000 1.415000 7.675000 1.655000 ;
        RECT 6.765000 1.655000 7.015000 1.785000 ;
        RECT 6.765000 1.955000 7.015000 2.465000 ;
        RECT 7.310000 0.905000 7.675000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.135000  1.785000 2.265000 1.955000 ;
      RECT 0.135000  1.955000 0.385000 2.465000 ;
      RECT 0.175000  0.085000 0.345000 0.895000 ;
      RECT 0.515000  0.255000 1.835000 0.475000 ;
      RECT 0.515000  0.475000 0.815000 0.905000 ;
      RECT 0.605000  2.125000 0.855000 2.635000 ;
      RECT 0.985000  0.645000 1.370000 0.735000 ;
      RECT 0.985000  0.735000 2.775000 0.905000 ;
      RECT 1.075000  1.955000 1.325000 2.465000 ;
      RECT 1.545000  2.125000 1.795000 2.635000 ;
      RECT 2.015000  1.955000 2.265000 2.295000 ;
      RECT 2.015000  2.295000 3.205000 2.465000 ;
      RECT 2.055000  0.085000 2.225000 0.555000 ;
      RECT 2.055000  1.455000 2.265000 1.785000 ;
      RECT 2.395000  0.255000 2.775000 0.735000 ;
      RECT 2.485000  0.905000 2.695000 1.415000 ;
      RECT 2.485000  1.415000 2.870000 1.965000 ;
      RECT 2.485000  1.965000 2.735000 2.125000 ;
      RECT 2.865000  1.075000 3.445000 1.245000 ;
      RECT 2.955000  2.135000 3.205000 2.295000 ;
      RECT 2.995000  0.085000 3.685000 0.555000 ;
      RECT 3.255000  0.725000 5.175000 0.905000 ;
      RECT 3.255000  0.905000 3.445000 1.075000 ;
      RECT 3.255000  1.245000 3.445000 1.495000 ;
      RECT 3.255000  1.495000 3.605000 1.665000 ;
      RECT 3.435000  1.665000 3.605000 1.785000 ;
      RECT 3.435000  1.785000 4.665000 1.965000 ;
      RECT 3.475000  2.135000 3.725000 2.635000 ;
      RECT 3.855000  0.255000 4.235000 0.725000 ;
      RECT 3.945000  2.135000 4.195000 2.295000 ;
      RECT 3.945000  2.295000 5.135000 2.465000 ;
      RECT 4.415000  1.965000 4.665000 2.125000 ;
      RECT 4.455000  0.085000 4.625000 0.555000 ;
      RECT 4.795000  0.255000 5.175000 0.725000 ;
      RECT 4.885000  1.785000 5.135000 2.295000 ;
      RECT 5.355000  1.795000 5.605000 2.635000 ;
      RECT 5.395000  0.085000 5.565000 0.895000 ;
      RECT 5.635000  1.075000 7.090000 1.245000 ;
      RECT 5.635000  1.245000 6.010000 1.615000 ;
      RECT 6.295000  2.165000 6.545000 2.635000 ;
      RECT 6.335000  0.085000 6.505000 0.555000 ;
      RECT 7.235000  1.825000 7.485000 2.635000 ;
      RECT 7.275000  0.085000 7.445000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.700000  1.445000 2.870000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.730000  1.445000 5.900000 1.615000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 2.640000 1.415000 2.980000 1.460000 ;
      RECT 2.640000 1.460000 5.960000 1.600000 ;
      RECT 2.640000 1.600000 2.980000 1.645000 ;
      RECT 5.670000 1.415000 5.960000 1.460000 ;
      RECT 5.670000 1.600000 5.960000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2o_4


MACRO sky130_fd_sc_hdll__a2bb2o_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 0.995000 1.815000 1.615000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.995000 2.335000 1.375000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.080000 0.765000 4.455000 1.655000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.300000 1.050000 3.760000 1.655000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 0.255000 0.830000 0.810000 ;
        RECT 0.525000 0.810000 0.745000 1.525000 ;
        RECT 0.525000 1.525000 0.830000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.600000 0.085000 ;
        RECT 0.185000  0.085000 0.355000 0.930000 ;
        RECT 1.000000  0.085000 1.480000 0.530000 ;
        RECT 2.155000  0.085000 2.890000 0.485000 ;
        RECT 3.905000  0.085000 4.355000 0.595000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.600000 2.805000 ;
        RECT 0.185000 1.445000 0.355000 2.635000 ;
        RECT 1.000000 2.235000 1.380000 2.635000 ;
        RECT 3.675000 2.175000 3.925000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.915000 0.995000 1.220000 1.325000 ;
      RECT 1.000000 1.325000 1.220000 1.805000 ;
      RECT 1.000000 1.805000 1.860000 1.975000 ;
      RECT 1.640000 1.975000 1.860000 2.200000 ;
      RECT 1.640000 2.200000 2.870000 2.370000 ;
      RECT 1.765000 0.255000 1.935000 0.655000 ;
      RECT 1.765000 0.655000 2.710000 0.825000 ;
      RECT 2.175000 1.545000 2.710000 1.715000 ;
      RECT 2.175000 1.715000 2.345000 1.905000 ;
      RECT 2.540000 0.825000 2.710000 1.545000 ;
      RECT 2.640000 1.895000 3.100000 2.065000 ;
      RECT 2.640000 2.065000 2.870000 2.200000 ;
      RECT 2.700000 2.370000 2.870000 2.465000 ;
      RECT 2.880000 0.700000 3.280000 0.870000 ;
      RECT 2.880000 0.870000 3.100000 1.895000 ;
      RECT 3.110000 0.255000 3.280000 0.700000 ;
      RECT 3.125000 2.255000 3.455000 2.425000 ;
      RECT 3.285000 1.835000 4.315000 2.005000 ;
      RECT 3.285000 2.005000 3.455000 2.255000 ;
      RECT 4.145000 2.005000 4.315000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2o_2


MACRO sky130_fd_sc_hdll__a2bb2o_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.995000 1.325000 1.615000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 0.995000 1.730000 1.375000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 0.765000 3.625000 1.655000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895000 1.040000 3.155000 1.655000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.345000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.140000 0.085000 ;
        RECT 0.515000  0.085000 0.995000 0.530000 ;
        RECT 1.670000  0.085000 2.390000 0.485000 ;
        RECT 3.490000  0.085000 3.940000 0.595000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.140000 2.805000 ;
        RECT 0.515000 2.235000 0.895000 2.635000 ;
        RECT 3.155000 2.175000 3.415000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515000 0.995000 0.685000 1.805000 ;
      RECT 0.515000 1.805000 1.375000 1.975000 ;
      RECT 1.155000 1.975000 1.375000 2.200000 ;
      RECT 1.155000 2.200000 2.385000 2.370000 ;
      RECT 1.265000 0.255000 1.435000 0.655000 ;
      RECT 1.265000 0.655000 2.210000 0.825000 ;
      RECT 1.690000 1.545000 2.210000 1.715000 ;
      RECT 1.690000 1.715000 1.860000 1.905000 ;
      RECT 2.040000 0.825000 2.210000 1.545000 ;
      RECT 2.130000 1.895000 2.600000 2.065000 ;
      RECT 2.130000 2.065000 2.385000 2.200000 ;
      RECT 2.130000 2.370000 2.385000 2.465000 ;
      RECT 2.380000 0.700000 2.855000 0.870000 ;
      RECT 2.380000 0.870000 2.600000 1.895000 ;
      RECT 2.605000 2.255000 2.945000 2.425000 ;
      RECT 2.685000 0.255000 2.855000 0.700000 ;
      RECT 2.775000 1.835000 3.815000 2.005000 ;
      RECT 2.775000 2.005000 2.945000 2.255000 ;
      RECT 3.635000 2.005000 3.815000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2o_1


MACRO sky130_fd_sc_hdll__and2b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.200000 0.625000 3.545000 1.745000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.995000 1.075000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.071500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.635000 1.535000 2.980000 1.745000 ;
        RECT 1.675000 0.495000 1.865000 0.615000 ;
        RECT 1.675000 0.615000 2.980000 0.825000 ;
        RECT 2.445000 0.825000 2.980000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.615000 ;
      RECT 0.090000  0.615000 1.455000 0.805000 ;
      RECT 0.090000  2.255000 0.425000 2.635000 ;
      RECT 0.165000  0.995000 0.425000 1.325000 ;
      RECT 0.165000  1.325000 0.335000 1.915000 ;
      RECT 0.165000  1.915000 3.940000 2.085000 ;
      RECT 0.515000  1.500000 1.415000 1.745000 ;
      RECT 1.055000  0.085000 1.385000 0.445000 ;
      RECT 1.090000  2.275000 1.420000 2.635000 ;
      RECT 1.245000  0.805000 1.455000 0.995000 ;
      RECT 1.245000  0.995000 2.175000 1.355000 ;
      RECT 1.245000  1.355000 1.420000 1.485000 ;
      RECT 1.245000  1.485000 1.415000 1.500000 ;
      RECT 2.035000  0.085000 2.415000 0.445000 ;
      RECT 2.055000  2.275000 2.435000 2.635000 ;
      RECT 2.995000  0.085000 3.375000 0.445000 ;
      RECT 2.995000  2.275000 3.375000 2.635000 ;
      RECT 3.725000  0.495000 3.940000 1.915000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2b_4


MACRO sky130_fd_sc_hdll__and2b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.445000 1.615000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.630000 1.645000 2.275000 1.955000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.505000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.580000 3.080000 2.365000 ;
        RECT 2.705000 0.255000 3.080000 0.775000 ;
        RECT 2.770000 0.775000 3.080000 1.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.590000 ;
      RECT 0.175000  1.785000 0.900000 2.015000 ;
      RECT 0.175000  2.015000 0.345000 2.445000 ;
      RECT 0.515000  2.185000 0.895000 2.635000 ;
      RECT 0.645000  0.280000 0.885000 0.655000 ;
      RECT 0.665000  0.655000 0.885000 0.805000 ;
      RECT 0.665000  0.805000 1.250000 1.135000 ;
      RECT 0.665000  1.135000 0.900000 1.785000 ;
      RECT 1.070000  1.305000 2.505000 1.325000 ;
      RECT 1.070000  1.325000 2.080000 1.475000 ;
      RECT 1.070000  1.475000 1.405000 2.420000 ;
      RECT 1.215000  0.270000 1.385000 0.415000 ;
      RECT 1.215000  0.415000 1.640000 0.610000 ;
      RECT 1.420000  0.610000 1.640000 0.945000 ;
      RECT 1.420000  0.945000 2.505000 1.305000 ;
      RECT 1.635000  2.165000 2.275000 2.635000 ;
      RECT 2.000000  0.085000 2.445000 0.580000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2b_1


MACRO sky130_fd_sc_hdll__and2b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.450000 1.615000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655000 1.645000 2.400000 1.955000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.762000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.575000 1.580000 3.090000 2.365000 ;
        RECT 2.695000 0.255000 3.090000 0.775000 ;
        RECT 2.755000 0.775000 3.090000 1.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.590000 ;
      RECT 0.175000  1.785000 0.905000 2.015000 ;
      RECT 0.175000  2.015000 0.345000 2.445000 ;
      RECT 0.515000  2.185000 0.895000 2.635000 ;
      RECT 0.645000  0.280000 0.885000 0.655000 ;
      RECT 0.670000  0.655000 0.885000 0.805000 ;
      RECT 0.670000  0.805000 1.275000 1.135000 ;
      RECT 0.670000  1.135000 0.905000 1.785000 ;
      RECT 1.095000  1.305000 2.535000 1.325000 ;
      RECT 1.095000  1.325000 2.105000 1.475000 ;
      RECT 1.095000  1.475000 1.430000 2.420000 ;
      RECT 1.215000  0.270000 1.385000 0.415000 ;
      RECT 1.215000  0.415000 1.665000 0.610000 ;
      RECT 1.445000  0.610000 1.665000 0.945000 ;
      RECT 1.445000  0.945000 2.535000 1.305000 ;
      RECT 1.660000  2.165000 2.395000 2.635000 ;
      RECT 2.105000  0.085000 2.475000 0.580000 ;
      RECT 3.325000  0.085000 3.595000 0.720000 ;
      RECT 3.325000  1.680000 3.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2b_2


MACRO sky130_fd_sc_hdll__or4bb_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815000 0.995000 3.570000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.680000 2.125000 3.370000 2.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.810000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.980000 0.995000 1.335000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.463700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.130000 0.415000 4.455000 0.760000 ;
        RECT 4.130000 1.495000 4.455000 2.465000 ;
        RECT 4.235000 0.760000 4.455000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.450000 0.400000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.865000 ;
      RECT 0.085000  1.865000 2.015000 2.035000 ;
      RECT 0.085000  2.035000 0.345000 2.455000 ;
      RECT 0.515000  2.205000 0.895000 2.635000 ;
      RECT 0.705000  0.085000 0.875000 0.825000 ;
      RECT 1.040000  1.525000 1.675000 1.695000 ;
      RECT 1.175000  0.450000 1.345000 0.655000 ;
      RECT 1.175000  0.655000 1.675000 0.825000 ;
      RECT 1.505000  0.825000 1.675000 1.075000 ;
      RECT 1.505000  1.075000 2.155000 1.245000 ;
      RECT 1.505000  1.245000 1.675000 1.525000 ;
      RECT 1.570000  0.085000 1.945000 0.485000 ;
      RECT 1.610000  2.205000 2.405000 2.375000 ;
      RECT 1.845000  1.415000 2.545000 1.585000 ;
      RECT 1.845000  1.585000 2.015000 1.865000 ;
      RECT 2.165000  0.305000 2.335000 0.655000 ;
      RECT 2.165000  0.655000 3.910000 0.825000 ;
      RECT 2.235000  1.785000 3.370000 1.955000 ;
      RECT 2.235000  1.955000 2.405000 2.205000 ;
      RECT 2.375000  0.995000 2.545000 1.415000 ;
      RECT 2.520000  0.085000 2.900000 0.485000 ;
      RECT 3.120000  0.305000 3.290000 0.655000 ;
      RECT 3.200000  1.495000 3.910000 1.665000 ;
      RECT 3.200000  1.665000 3.370000 1.785000 ;
      RECT 3.460000  0.085000 3.890000 0.485000 ;
      RECT 3.590000  1.835000 3.870000 2.635000 ;
      RECT 3.740000  0.825000 3.910000 0.995000 ;
      RECT 3.740000  0.995000 4.030000 1.325000 ;
      RECT 3.740000  1.325000 3.910000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4bb_1


MACRO sky130_fd_sc_hdll__or4bb_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.840000 0.995000 3.595000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705000 2.125000 3.395000 2.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.830000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.995000 1.340000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.155000 0.415000 4.455000 0.760000 ;
        RECT 4.155000 1.495000 4.455000 2.465000 ;
        RECT 4.260000 0.760000 4.455000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.450000 0.405000 0.825000 ;
      RECT 0.085000  0.825000 0.260000 1.865000 ;
      RECT 0.085000  1.865000 2.040000 2.035000 ;
      RECT 0.085000  2.035000 0.345000 2.455000 ;
      RECT 0.515000  2.205000 0.895000 2.635000 ;
      RECT 0.710000  0.085000 0.880000 0.825000 ;
      RECT 1.045000  1.525000 1.700000 1.695000 ;
      RECT 1.180000  0.450000 1.350000 0.655000 ;
      RECT 1.180000  0.655000 1.700000 0.825000 ;
      RECT 1.510000  0.825000 1.700000 1.075000 ;
      RECT 1.510000  1.075000 1.955000 1.245000 ;
      RECT 1.510000  1.245000 1.700000 1.525000 ;
      RECT 1.595000  0.085000 1.970000 0.485000 ;
      RECT 1.635000  2.205000 2.430000 2.375000 ;
      RECT 1.870000  1.415000 2.570000 1.585000 ;
      RECT 1.870000  1.585000 2.040000 1.865000 ;
      RECT 2.190000  0.305000 2.360000 0.655000 ;
      RECT 2.190000  0.655000 3.935000 0.825000 ;
      RECT 2.260000  1.785000 3.395000 1.955000 ;
      RECT 2.260000  1.955000 2.430000 2.205000 ;
      RECT 2.400000  0.995000 2.570000 1.415000 ;
      RECT 2.545000  0.085000 2.925000 0.485000 ;
      RECT 3.145000  0.305000 3.315000 0.655000 ;
      RECT 3.225000  1.495000 3.935000 1.665000 ;
      RECT 3.225000  1.665000 3.395000 1.785000 ;
      RECT 3.485000  0.085000 3.915000 0.485000 ;
      RECT 3.615000  1.835000 3.895000 2.635000 ;
      RECT 3.765000  0.825000 3.935000 0.995000 ;
      RECT 3.765000  0.995000 4.040000 1.325000 ;
      RECT 3.765000  1.325000 3.935000 1.495000 ;
      RECT 4.650000  0.085000 4.820000 0.915000 ;
      RECT 4.650000  1.440000 4.820000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4bb_2


MACRO sky130_fd_sc_hdll__or4bb_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.400000 3.675000 1.615000 ;
        RECT 3.455000 0.995000 3.675000 1.400000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.845000 0.995000 3.145000 2.375000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 0.995000 0.825000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 0.995000 1.335000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.185000 1.455000 5.855000 1.625000 ;
        RECT 4.185000 1.625000 4.435000 2.465000 ;
        RECT 4.225000 0.255000 4.475000 0.725000 ;
        RECT 4.225000 0.725000 5.855000 0.905000 ;
        RECT 5.035000 0.255000 5.415000 0.725000 ;
        RECT 5.125000 1.625000 5.375000 2.465000 ;
        RECT 5.625000 0.905000 5.855000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.095000  0.450000 0.400000 0.825000 ;
      RECT 0.095000  0.825000 0.265000 1.900000 ;
      RECT 0.095000  1.900000 1.395000 2.070000 ;
      RECT 0.095000  2.070000 0.345000 2.455000 ;
      RECT 0.515000  2.240000 0.895000 2.635000 ;
      RECT 0.705000  0.085000 0.875000 0.825000 ;
      RECT 1.040000  1.560000 1.695000 1.730000 ;
      RECT 1.175000  0.450000 1.345000 0.655000 ;
      RECT 1.175000  0.655000 1.695000 0.825000 ;
      RECT 1.225000  2.070000 1.395000 2.295000 ;
      RECT 1.225000  2.295000 2.565000 2.465000 ;
      RECT 1.505000  0.825000 1.695000 0.995000 ;
      RECT 1.505000  0.995000 1.795000 1.325000 ;
      RECT 1.505000  1.325000 1.695000 1.560000 ;
      RECT 1.610000  1.955000 2.225000 2.125000 ;
      RECT 1.615000  0.085000 1.945000 0.480000 ;
      RECT 2.035000  0.655000 4.015000 0.825000 ;
      RECT 2.035000  0.825000 2.225000 1.955000 ;
      RECT 2.245000  0.305000 2.415000 0.655000 ;
      RECT 2.395000  0.995000 2.565000 2.295000 ;
      RECT 2.585000  0.085000 2.965000 0.485000 ;
      RECT 3.185000  0.305000 3.355000 0.655000 ;
      RECT 3.615000  0.085000 3.995000 0.485000 ;
      RECT 3.660000  1.795000 3.910000 2.635000 ;
      RECT 3.845000  0.825000 4.015000 1.075000 ;
      RECT 3.845000  1.075000 5.445000 1.245000 ;
      RECT 4.655000  1.795000 4.905000 2.635000 ;
      RECT 4.695000  0.085000 4.865000 0.555000 ;
      RECT 5.595000  1.795000 5.845000 2.635000 ;
      RECT 5.635000  0.085000 5.805000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or4bb_4


MACRO sky130_fd_sc_hdll__inputiso0p_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.645000 1.835000 1.955000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.445000 1.615000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.580000 3.080000 2.365000 ;
        RECT 2.620000 0.255000 3.080000 0.775000 ;
        RECT 2.905000 0.775000 3.080000 1.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.590000 ;
      RECT 0.175000  1.785000 0.895000 2.015000 ;
      RECT 0.175000  2.015000 0.345000 2.445000 ;
      RECT 0.515000  2.185000 0.895000 2.635000 ;
      RECT 0.645000  0.280000 0.885000 0.805000 ;
      RECT 0.645000  0.805000 1.180000 1.135000 ;
      RECT 0.645000  1.135000 0.895000 1.785000 ;
      RECT 1.065000  1.305000 2.475000 1.325000 ;
      RECT 1.065000  1.325000 1.885000 1.475000 ;
      RECT 1.065000  1.475000 1.335000 2.420000 ;
      RECT 1.165000  0.270000 1.335000 0.415000 ;
      RECT 1.165000  0.415000 1.590000 0.610000 ;
      RECT 1.350000  0.610000 1.590000 0.945000 ;
      RECT 1.350000  0.945000 2.475000 1.305000 ;
      RECT 1.565000  2.165000 2.325000 2.635000 ;
      RECT 2.070000  0.085000 2.400000 0.580000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inputiso0p_1


MACRO sky130_fd_sc_hdll__o31ai_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.740000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.055000 1.930000 1.425000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.150000 1.055000 4.005000 1.425000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 1.055000 6.590000 1.275000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.165000 1.055000 8.585000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.851000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 1.445000 8.625000 1.695000 ;
        RECT 6.420000 1.695000 6.590000 2.465000 ;
        RECT 6.760000 0.645000 8.080000 0.885000 ;
        RECT 6.760000 0.885000 6.995000 1.445000 ;
        RECT 7.360000 1.695000 7.530000 2.465000 ;
        RECT 8.300000 1.695000 8.625000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.090000  0.255000 0.445000 0.715000 ;
      RECT 0.090000  0.715000 6.590000 0.885000 ;
      RECT 0.090000  1.595000 2.325000 1.895000 ;
      RECT 0.090000  1.895000 0.445000 2.465000 ;
      RECT 0.665000  0.085000 0.835000 0.545000 ;
      RECT 0.665000  2.065000 0.835000 2.635000 ;
      RECT 1.005000  0.255000 1.385000 0.715000 ;
      RECT 1.005000  1.895000 1.385000 2.465000 ;
      RECT 1.605000  0.085000 1.775000 0.545000 ;
      RECT 1.605000  2.065000 1.775000 2.635000 ;
      RECT 1.945000  0.255000 2.325000 0.715000 ;
      RECT 1.945000  1.895000 2.325000 2.205000 ;
      RECT 1.945000  2.205000 4.285000 2.465000 ;
      RECT 2.545000  0.085000 2.715000 0.545000 ;
      RECT 2.545000  1.595000 4.005000 1.765000 ;
      RECT 2.545000  1.765000 2.715000 2.035000 ;
      RECT 2.885000  0.255000 3.265000 0.715000 ;
      RECT 2.885000  1.935000 3.265000 2.205000 ;
      RECT 3.485000  0.085000 3.655000 0.545000 ;
      RECT 3.485000  1.765000 4.005000 1.865000 ;
      RECT 3.485000  1.865000 6.200000 2.035000 ;
      RECT 3.825000  0.255000 4.205000 0.715000 ;
      RECT 4.445000  0.085000 5.140000 0.545000 ;
      RECT 4.530000  2.035000 6.200000 2.465000 ;
      RECT 5.360000  0.395000 5.530000 0.715000 ;
      RECT 5.790000  0.085000 6.160000 0.545000 ;
      RECT 6.420000  0.255000 8.585000 0.475000 ;
      RECT 6.420000  0.475000 6.590000 0.715000 ;
      RECT 6.760000  1.890000 7.140000 2.635000 ;
      RECT 7.700000  1.890000 8.080000 2.635000 ;
      RECT 8.300000  0.475000 8.585000 0.885000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o31ai_4


MACRO sky130_fd_sc_hdll__o31ai_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.055000 1.310000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 1.055000 2.420000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.700000 1.055000 3.555000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.630000 0.755000 4.970000 1.325000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.136000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.585000 1.495000 4.965000 1.665000 ;
        RECT 2.585000 1.665000 2.915000 2.125000 ;
        RECT 3.475000 1.665000 3.855000 2.465000 ;
        RECT 4.075000 0.595000 4.455000 1.495000 ;
        RECT 4.625000 1.665000 4.965000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.090000  0.255000 0.445000 0.715000 ;
      RECT 0.090000  0.715000 3.855000 0.885000 ;
      RECT 0.090000  1.495000 2.325000 1.665000 ;
      RECT 0.090000  1.665000 0.445000 2.465000 ;
      RECT 0.665000  0.085000 0.835000 0.545000 ;
      RECT 0.665000  1.835000 0.835000 2.635000 ;
      RECT 1.005000  0.255000 1.385000 0.715000 ;
      RECT 1.005000  1.665000 1.385000 2.465000 ;
      RECT 1.605000  0.085000 2.165000 0.545000 ;
      RECT 1.605000  1.835000 1.775000 2.295000 ;
      RECT 1.605000  2.295000 3.305000 2.465000 ;
      RECT 1.945000  1.665000 2.325000 2.125000 ;
      RECT 2.425000  0.255000 2.755000 0.715000 ;
      RECT 2.925000  0.085000 3.305000 0.545000 ;
      RECT 3.135000  1.835000 3.305000 2.295000 ;
      RECT 3.475000  0.255000 4.965000 0.425000 ;
      RECT 3.475000  0.425000 3.855000 0.715000 ;
      RECT 4.075000  1.835000 4.405000 2.635000 ;
      RECT 4.630000  0.425000 4.965000 0.585000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o31ai_2


MACRO sky130_fd_sc_hdll__o31ai_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.435000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.075000 1.105000 2.465000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.075000 1.695000 1.325000 ;
        RECT 1.455000 1.325000 1.695000 2.405000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 0.995000 2.650000 1.325000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.833500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 0.260000 2.495000 0.825000 ;
        RECT 1.885000 0.825000 2.155000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT -0.015000  2.635000 2.760000 2.805000 ;
      RECT  0.000000 -0.085000 2.760000 0.085000 ;
      RECT  0.085000  1.495000 0.420000 2.635000 ;
      RECT  0.175000  0.085000 0.345000 0.905000 ;
      RECT  0.515000  0.255000 0.895000 0.735000 ;
      RECT  0.515000  0.735000 1.715000 0.905000 ;
      RECT  1.125000  0.085000 1.295000 0.565000 ;
      RECT  1.465000  0.460000 1.715000 0.735000 ;
      RECT  2.355000  1.495000 2.525000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o31ai_1


MACRO sky130_fd_sc_hdll__a21oi_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.895000 0.995000 1.575000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.035000 0.695000 1.495000 ;
        RECT 0.145000 1.495000 2.130000 1.675000 ;
        RECT 1.755000 1.075000 2.130000 1.495000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 0.995000 3.535000 1.625000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.745000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 0.255000 1.400000 0.615000 ;
        RECT 1.005000 0.615000 2.865000 0.785000 ;
        RECT 2.410000 0.785000 2.865000 1.330000 ;
        RECT 2.515000 1.330000 2.865000 2.115000 ;
        RECT 2.545000 0.255000 2.865000 0.615000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.100000  0.085000 0.395000 0.865000 ;
      RECT 0.110000  1.855000 2.345000 2.025000 ;
      RECT 0.110000  2.025000 1.320000 2.105000 ;
      RECT 0.110000  2.105000 0.370000 2.465000 ;
      RECT 0.540000  2.275000 0.920000 2.635000 ;
      RECT 1.150000  2.105000 1.320000 2.465000 ;
      RECT 1.625000  2.195000 1.795000 2.635000 ;
      RECT 1.910000  0.085000 2.290000 0.445000 ;
      RECT 2.015000  2.025000 2.345000 2.285000 ;
      RECT 2.015000  2.285000 3.390000 2.465000 ;
      RECT 3.085000  1.795000 3.390000 2.285000 ;
      RECT 3.095000  0.085000 3.425000 0.825000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21oi_2


MACRO sky130_fd_sc_hdll__a21oi_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815000 1.065000 4.400000 1.310000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.250000 1.065000 2.645000 1.480000 ;
        RECT 2.250000 1.480000 6.070000 1.705000 ;
        RECT 4.675000 1.075000 6.070000 1.480000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.400000 1.035000 ;
        RECT 0.090000 1.035000 1.580000 1.415000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.523000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.630000 1.585000 2.080000 1.705000 ;
        RECT 0.630000 1.705000 1.895000 2.035000 ;
        RECT 0.645000 0.370000 0.835000 0.615000 ;
        RECT 0.645000 0.615000 1.795000 0.695000 ;
        RECT 0.645000 0.695000 4.305000 0.865000 ;
        RECT 1.605000 0.255000 1.795000 0.615000 ;
        RECT 1.750000 0.865000 4.305000 0.895000 ;
        RECT 1.750000 0.895000 2.080000 1.585000 ;
        RECT 2.475000 0.675000 4.305000 0.695000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.805000 ;
      RECT 0.180000  1.795000 0.375000 2.215000 ;
      RECT 0.180000  2.215000 2.315000 2.465000 ;
      RECT 1.005000  0.085000 1.385000 0.445000 ;
      RECT 1.005000  2.205000 2.315000 2.215000 ;
      RECT 1.985000  0.085000 2.315000 0.525000 ;
      RECT 2.115000  1.875000 6.225000 2.105000 ;
      RECT 2.115000  2.105000 2.315000 2.205000 ;
      RECT 2.485000  0.255000 4.785000 0.505000 ;
      RECT 2.485000  2.275000 2.865000 2.635000 ;
      RECT 3.085000  2.105000 3.275000 2.465000 ;
      RECT 3.445000  2.275000 3.825000 2.635000 ;
      RECT 4.045000  2.105000 4.235000 2.465000 ;
      RECT 4.405000  2.275000 4.785000 2.635000 ;
      RECT 4.525000  0.505000 4.785000 0.735000 ;
      RECT 4.525000  0.735000 5.745000 0.905000 ;
      RECT 5.005000  0.085000 5.195000 0.565000 ;
      RECT 5.005000  2.105000 5.185000 2.465000 ;
      RECT 5.365000  0.255000 5.745000 0.735000 ;
      RECT 5.365000  2.275000 5.745000 2.635000 ;
      RECT 5.965000  0.085000 6.225000 0.885000 ;
      RECT 5.965000  2.105000 6.225000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21oi_4


MACRO sky130_fd_sc_hdll__a21oi_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.900000 0.995000 1.295000 1.325000 ;
        RECT 1.065000 0.375000 1.295000 0.995000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 1.820000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.675000 0.335000 1.325000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.489500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.495000 0.730000 1.685000 ;
        RECT 0.095000 1.685000 0.370000 2.455000 ;
        RECT 0.505000 0.645000 0.885000 0.825000 ;
        RECT 0.505000 0.825000 0.730000 1.495000 ;
        RECT 0.660000 0.265000 0.885000 0.645000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.110000  0.085000 0.440000 0.475000 ;
      RECT 0.540000  1.855000 1.895000 2.025000 ;
      RECT 0.540000  2.025000 0.920000 2.455000 ;
      RECT 0.900000  1.525000 1.895000 1.855000 ;
      RECT 1.140000  2.195000 1.335000 2.635000 ;
      RECT 1.515000  2.025000 1.895000 2.455000 ;
      RECT 1.595000  0.085000 1.895000 0.815000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21oi_1


MACRO sky130_fd_sc_hdll__and3b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.745000 0.410000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.915000 2.125000 2.490000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.305000 2.370000 0.765000 ;
        RECT 1.985000 0.765000 2.620000 1.245000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.125000 1.795000 3.590000 2.465000 ;
        RECT 3.165000 0.255000 3.570000 0.715000 ;
        RECT 3.240000 0.715000 3.570000 0.925000 ;
        RECT 3.240000 0.925000 4.040000 1.445000 ;
        RECT 3.240000 1.445000 3.590000 1.795000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.085000 0.355000 0.575000 ;
      RECT 0.085000  1.575000 0.400000 2.635000 ;
      RECT 0.630000  0.305000 0.905000 1.015000 ;
      RECT 0.630000  1.015000 1.465000 1.245000 ;
      RECT 0.630000  1.245000 0.905000 1.905000 ;
      RECT 1.080000  2.130000 1.745000 2.635000 ;
      RECT 1.100000  1.425000 3.020000 1.595000 ;
      RECT 1.100000  1.595000 1.335000 1.960000 ;
      RECT 1.105000  0.305000 1.815000 0.570000 ;
      RECT 1.505000  1.765000 1.885000 1.955000 ;
      RECT 1.505000  1.955000 1.745000 2.130000 ;
      RECT 1.645000  0.570000 1.815000 1.425000 ;
      RECT 2.160000  1.595000 2.350000 1.890000 ;
      RECT 2.610000  0.085000 2.940000 0.580000 ;
      RECT 2.660000  1.790000 2.875000 2.635000 ;
      RECT 2.790000  0.995000 3.020000 1.425000 ;
      RECT 3.760000  0.085000 4.025000 0.745000 ;
      RECT 3.760000  1.625000 4.025000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3b_2


MACRO sky130_fd_sc_hdll__and3b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.955000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.920000 2.125000 2.495000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.280000 0.305000 2.645000 1.255000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.270000 1.765000 3.535000 2.465000 ;
        RECT 3.275000 0.255000 3.535000 0.735000 ;
        RECT 3.365000 0.735000 3.535000 1.765000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.905000 ;
      RECT 0.085000  2.125000 0.345000 2.635000 ;
      RECT 0.515000  0.485000 0.895000 0.905000 ;
      RECT 0.645000  0.905000 0.895000 0.995000 ;
      RECT 0.645000  0.995000 1.520000 1.245000 ;
      RECT 0.645000  1.245000 0.815000 2.465000 ;
      RECT 1.085000  1.425000 3.185000 1.575000 ;
      RECT 1.085000  1.575000 3.050000 1.595000 ;
      RECT 1.085000  1.595000 1.335000 1.940000 ;
      RECT 1.085000  2.130000 1.750000 2.635000 ;
      RECT 1.105000  0.285000 1.945000 0.550000 ;
      RECT 1.505000  1.765000 1.885000 1.955000 ;
      RECT 1.505000  1.955000 1.750000 2.130000 ;
      RECT 1.690000  0.550000 1.945000 1.425000 ;
      RECT 2.155000  1.595000 3.050000 1.890000 ;
      RECT 2.795000  2.090000 3.010000 2.635000 ;
      RECT 2.815000  0.085000 3.105000 0.625000 ;
      RECT 2.965000  0.975000 3.185000 1.425000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3b_1


MACRO sky130_fd_sc_hdll__and3b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 0.615000 4.455000 1.705000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 0.725000 1.285000 1.340000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.490000 0.995000 1.865000 1.340000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.071500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 1.535000 3.995000 1.705000 ;
        RECT 2.485000 0.515000 2.675000 0.615000 ;
        RECT 2.485000 0.615000 3.995000 0.845000 ;
        RECT 3.365000 0.255000 3.635000 0.615000 ;
        RECT 3.570000 0.845000 3.995000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.150000  0.255000 0.635000 0.355000 ;
      RECT 0.150000  0.355000 1.700000 0.545000 ;
      RECT 0.150000  0.545000 0.635000 0.805000 ;
      RECT 0.150000  0.805000 0.370000 1.495000 ;
      RECT 0.150000  1.495000 0.510000 2.165000 ;
      RECT 0.540000  0.995000 0.865000 1.325000 ;
      RECT 0.680000  1.325000 0.865000 1.875000 ;
      RECT 0.680000  1.875000 4.905000 2.105000 ;
      RECT 0.730000  2.275000 1.230000 2.635000 ;
      RECT 1.330000  1.525000 2.205000 1.695000 ;
      RECT 1.520000  0.545000 1.700000 0.615000 ;
      RECT 1.520000  0.615000 2.265000 0.805000 ;
      RECT 1.895000  2.275000 2.225000 2.635000 ;
      RECT 1.930000  0.085000 2.260000 0.445000 ;
      RECT 2.035000  0.805000 2.265000 1.020000 ;
      RECT 2.035000  1.020000 3.400000 1.355000 ;
      RECT 2.035000  1.355000 2.205000 1.525000 ;
      RECT 2.845000  0.085000 3.195000 0.445000 ;
      RECT 2.845000  2.275000 3.230000 2.635000 ;
      RECT 3.805000  0.085000 4.185000 0.445000 ;
      RECT 3.805000  2.275000 4.185000 2.635000 ;
      RECT 4.625000  0.425000 4.905000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3b_4


MACRO sky130_fd_sc_hdll__nor4bb_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.360000 0.995000 3.665000 1.705000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.820000 0.995000 3.130000 2.410000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.830000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.995000 1.340000 1.325000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.660000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.575000 1.955000 2.210000 2.125000 ;
        RECT 1.960000 0.655000 3.340000 0.825000 ;
        RECT 1.960000 0.825000 2.210000 1.955000 ;
        RECT 2.170000 0.300000 2.370000 0.655000 ;
        RECT 3.140000 0.310000 3.340000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.450000 0.405000 0.825000 ;
      RECT 0.085000  0.825000 0.260000 1.885000 ;
      RECT 0.085000  1.885000 1.305000 2.070000 ;
      RECT 0.085000  2.070000 0.345000 2.455000 ;
      RECT 0.515000  2.240000 0.895000 2.635000 ;
      RECT 0.705000  0.085000 0.875000 0.825000 ;
      RECT 1.100000  1.525000 1.790000 1.715000 ;
      RECT 1.135000  2.070000 1.305000 2.295000 ;
      RECT 1.135000  2.295000 2.615000 2.465000 ;
      RECT 1.175000  0.450000 1.345000 0.655000 ;
      RECT 1.175000  0.655000 1.790000 0.825000 ;
      RECT 1.620000  0.085000 1.950000 0.480000 ;
      RECT 1.620000  0.825000 1.790000 1.525000 ;
      RECT 2.380000  0.995000 2.615000 2.295000 ;
      RECT 2.590000  0.085000 2.920000 0.485000 ;
      RECT 3.510000  0.085000 3.990000 0.825000 ;
      RECT 3.510000  1.875000 3.990000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4bb_1


MACRO sky130_fd_sc_hdll__nor4bb_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.12000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.075000 1.075000 10.010000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.650000 1.075000 7.805000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.445000 1.365000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.075000 1.395000 1.325000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  2.374000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 1.415000 3.435000 1.705000 ;
        RECT 2.035000 0.255000 2.415000 0.725000 ;
        RECT 2.035000 0.725000 9.515000 0.905000 ;
        RECT 2.975000 0.255000 3.355000 0.725000 ;
        RECT 3.265000 0.905000 3.435000 1.415000 ;
        RECT 3.915000 0.255000 4.295000 0.725000 ;
        RECT 4.855000 0.255000 5.235000 0.725000 ;
        RECT 6.315000 0.255000 6.695000 0.725000 ;
        RECT 7.255000 0.255000 7.635000 0.725000 ;
        RECT 8.195000 0.255000 8.575000 0.725000 ;
        RECT 9.135000 0.255000 9.515000 0.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.255000  0.445000 0.725000 ;
      RECT 0.085000  0.725000  0.835000 0.895000 ;
      RECT 0.085000  1.535000  0.835000 1.875000 ;
      RECT 0.085000  1.875000  3.825000 2.045000 ;
      RECT 0.085000  2.045000  0.365000 2.465000 ;
      RECT 0.535000  2.215000  0.915000 2.635000 ;
      RECT 0.665000  0.085000  0.835000 0.555000 ;
      RECT 0.665000  0.895000  0.835000 1.535000 ;
      RECT 1.005000  0.255000  1.385000 0.735000 ;
      RECT 1.005000  0.735000  1.735000 0.905000 ;
      RECT 1.005000  1.535000  1.735000 1.705000 ;
      RECT 1.565000  0.905000  1.735000 1.075000 ;
      RECT 1.565000  1.075000  3.095000 1.245000 ;
      RECT 1.565000  1.245000  1.735000 1.535000 ;
      RECT 1.615000  2.215000  3.825000 2.295000 ;
      RECT 1.615000  2.295000  5.695000 2.465000 ;
      RECT 1.695000  0.085000  1.865000 0.555000 ;
      RECT 2.635000  0.085000  2.805000 0.555000 ;
      RECT 3.575000  0.085000  3.745000 0.555000 ;
      RECT 3.655000  1.075000  5.405000 1.285000 ;
      RECT 3.655000  1.285000  3.825000 1.875000 ;
      RECT 4.045000  1.455000  7.595000 1.625000 ;
      RECT 4.045000  1.625000  4.255000 2.125000 ;
      RECT 4.475000  1.795000  4.725000 2.295000 ;
      RECT 4.515000  0.085000  4.685000 0.555000 ;
      RECT 4.945000  1.625000  5.195000 2.125000 ;
      RECT 5.415000  1.795000  5.695000 2.295000 ;
      RECT 5.455000  0.085000  6.145000 0.555000 ;
      RECT 5.880000  1.795000  6.185000 2.295000 ;
      RECT 5.880000  2.295000  8.065000 2.465000 ;
      RECT 6.405000  1.625000  6.655000 2.125000 ;
      RECT 6.875000  1.795000  7.125000 2.295000 ;
      RECT 6.915000  0.085000  7.085000 0.555000 ;
      RECT 7.345000  1.625000  7.595000 2.125000 ;
      RECT 7.815000  1.455000 10.010000 1.625000 ;
      RECT 7.815000  1.625000  8.065000 2.295000 ;
      RECT 7.855000  0.085000  8.025000 0.555000 ;
      RECT 8.285000  1.795000  8.535000 2.635000 ;
      RECT 8.755000  1.625000  9.005000 2.465000 ;
      RECT 8.795000  0.085000  8.965000 0.555000 ;
      RECT 9.225000  1.795000  9.475000 2.635000 ;
      RECT 9.695000  1.625000 10.010000 2.465000 ;
      RECT 9.735000  0.085000 10.010000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4bb_4


MACRO sky130_fd_sc_hdll__nor4bb_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.465000 1.075000 6.330000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.400000 1.075000 5.295000 1.275000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.995000 1.270000 1.325000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.830000 1.695000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.219500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095000 0.255000 2.475000 0.725000 ;
        RECT 2.095000 0.725000 5.835000 0.905000 ;
        RECT 3.035000 0.255000 3.415000 0.725000 ;
        RECT 3.035000 1.445000 4.230000 1.705000 ;
        RECT 3.810000 0.905000 4.230000 1.445000 ;
        RECT 4.515000 0.255000 4.895000 0.725000 ;
        RECT 5.455000 0.255000 5.835000 0.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  0.450000 0.465000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.885000 ;
      RECT 0.085000  1.885000 1.950000 2.055000 ;
      RECT 0.085000  2.055000 0.345000 2.455000 ;
      RECT 0.515000  2.240000 0.895000 2.635000 ;
      RECT 0.685000  0.085000 0.855000 0.825000 ;
      RECT 1.045000  1.525000 1.610000 1.715000 ;
      RECT 1.155000  0.450000 1.350000 0.655000 ;
      RECT 1.155000  0.655000 1.610000 0.825000 ;
      RECT 1.440000  0.825000 1.610000 1.075000 ;
      RECT 1.440000  1.075000 2.475000 1.245000 ;
      RECT 1.440000  1.245000 1.610000 1.525000 ;
      RECT 1.595000  0.085000 1.925000 0.480000 ;
      RECT 1.675000  2.225000 3.885000 2.465000 ;
      RECT 1.780000  1.415000 2.865000 1.585000 ;
      RECT 1.780000  1.585000 1.950000 1.885000 ;
      RECT 2.145000  1.875000 4.895000 2.045000 ;
      RECT 2.695000  0.085000 2.865000 0.555000 ;
      RECT 2.695000  1.075000 3.640000 1.275000 ;
      RECT 2.695000  1.275000 2.865000 1.415000 ;
      RECT 3.635000  0.085000 4.345000 0.555000 ;
      RECT 4.095000  2.215000 5.325000 2.465000 ;
      RECT 4.605000  1.455000 4.895000 1.875000 ;
      RECT 5.115000  0.085000 5.285000 0.555000 ;
      RECT 5.115000  1.455000 6.305000 1.625000 ;
      RECT 5.115000  1.625000 5.325000 2.215000 ;
      RECT 5.545000  1.795000 5.755000 2.635000 ;
      RECT 5.925000  1.625000 6.305000 2.465000 ;
      RECT 6.055000  0.085000 6.330000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4bb_2


MACRO sky130_fd_sc_hdll__or2b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 2.085000 1.835000 2.415000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.325000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.455500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.605000 0.415000 3.090000 0.760000 ;
        RECT 2.605000 1.495000 3.090000 2.465000 ;
        RECT 2.705000 0.760000 3.090000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.110000  0.265000 0.420000 0.735000 ;
      RECT 0.110000  0.735000 0.895000 0.905000 ;
      RECT 0.640000  0.085000 1.375000 0.565000 ;
      RECT 0.645000  0.905000 0.895000 0.995000 ;
      RECT 0.645000  0.995000 1.385000 1.325000 ;
      RECT 0.645000  1.325000 0.815000 1.885000 ;
      RECT 1.040000  1.495000 2.385000 1.665000 ;
      RECT 1.040000  1.665000 1.460000 1.915000 ;
      RECT 1.595000  0.305000 1.765000 0.655000 ;
      RECT 1.595000  0.655000 2.385000 0.825000 ;
      RECT 1.935000  0.085000 2.365000 0.485000 ;
      RECT 2.065000  1.835000 2.345000 2.635000 ;
      RECT 2.215000  0.825000 2.385000 0.995000 ;
      RECT 2.215000  0.995000 2.445000 1.325000 ;
      RECT 2.215000  1.325000 2.385000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2b_1


MACRO sky130_fd_sc_hdll__or2b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.730000 1.075000 2.470000 1.275000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.955000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.475000 0.290000 2.855000 0.735000 ;
        RECT 2.475000 0.735000 4.490000 0.905000 ;
        RECT 2.565000 1.785000 3.755000 1.955000 ;
        RECT 2.565000 1.955000 2.815000 2.465000 ;
        RECT 3.080000 1.445000 4.490000 1.615000 ;
        RECT 3.080000 1.615000 3.755000 1.785000 ;
        RECT 3.415000 0.290000 3.795000 0.735000 ;
        RECT 3.505000 1.955000 3.755000 2.465000 ;
        RECT 4.105000 0.905000 4.490000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  2.125000 0.345000 2.635000 ;
      RECT 0.110000  0.265000 0.420000 0.735000 ;
      RECT 0.110000  0.735000 0.895000 0.905000 ;
      RECT 0.640000  0.085000 1.295000 0.565000 ;
      RECT 0.645000  0.905000 0.895000 0.995000 ;
      RECT 0.645000  0.995000 1.170000 1.325000 ;
      RECT 0.645000  1.325000 0.815000 2.465000 ;
      RECT 1.040000  1.495000 2.860000 1.615000 ;
      RECT 1.040000  1.615000 1.560000 2.465000 ;
      RECT 1.340000  0.735000 1.845000 0.905000 ;
      RECT 1.340000  0.905000 1.560000 1.445000 ;
      RECT 1.340000  1.445000 2.860000 1.495000 ;
      RECT 1.465000  0.305000 1.845000 0.735000 ;
      RECT 2.065000  1.835000 2.345000 2.635000 ;
      RECT 2.130000  0.085000 2.305000 0.905000 ;
      RECT 2.690000  1.075000 3.800000 1.245000 ;
      RECT 2.690000  1.245000 2.860000 1.445000 ;
      RECT 3.035000  2.135000 3.285000 2.635000 ;
      RECT 3.075000  0.085000 3.245000 0.550000 ;
      RECT 3.975000  1.795000 4.225000 2.635000 ;
      RECT 4.015000  0.085000 4.185000 0.550000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2b_4


MACRO sky130_fd_sc_hdll__or2b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 2.085000 1.830000 2.415000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.325000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.811500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 0.415000 3.110000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.105000  0.265000 0.420000 0.735000 ;
      RECT 0.105000  0.735000 0.890000 0.905000 ;
      RECT 0.640000  0.085000 1.370000 0.565000 ;
      RECT 0.645000  0.905000 0.890000 0.995000 ;
      RECT 0.645000  0.995000 1.380000 1.325000 ;
      RECT 0.645000  1.325000 0.815000 1.885000 ;
      RECT 1.035000  1.495000 2.440000 1.665000 ;
      RECT 1.035000  1.665000 1.455000 1.915000 ;
      RECT 1.590000  0.305000 1.760000 0.655000 ;
      RECT 1.590000  0.655000 2.440000 0.825000 ;
      RECT 2.030000  0.085000 2.360000 0.485000 ;
      RECT 2.060000  1.835000 2.340000 2.635000 ;
      RECT 2.270000  0.825000 2.440000 1.495000 ;
      RECT 3.285000  0.085000 3.520000 0.925000 ;
      RECT 3.285000  1.460000 3.520000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2b_2


MACRO sky130_fd_sc_hdll__einvn_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 1.075000 3.535000 1.275000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.516600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.325000 1.385000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.768000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.145000 1.445000 3.535000 1.695000 ;
        RECT 2.445000 0.595000 2.815000 1.445000 ;
        RECT 3.035000 1.695000 3.535000 2.465000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.890000 0.825000 ;
      RECT 0.085000  1.555000 0.945000 1.725000 ;
      RECT 0.085000  1.725000 0.345000 2.465000 ;
      RECT 0.495000  0.825000 0.890000 0.995000 ;
      RECT 0.495000  0.995000 2.180000 1.275000 ;
      RECT 0.495000  1.275000 0.945000 1.555000 ;
      RECT 0.515000  0.085000 0.895000 0.485000 ;
      RECT 0.515000  1.895000 0.945000 2.635000 ;
      RECT 1.065000  0.255000 1.380000 0.655000 ;
      RECT 1.065000  0.655000 2.270000 0.825000 ;
      RECT 1.170000  1.445000 1.925000 1.865000 ;
      RECT 1.170000  1.865000 2.865000 2.085000 ;
      RECT 1.170000  2.085000 1.340000 2.465000 ;
      RECT 1.510000  2.255000 2.475000 2.635000 ;
      RECT 1.600000  0.085000 1.930000 0.485000 ;
      RECT 2.100000  0.255000 3.435000 0.425000 ;
      RECT 2.100000  0.425000 2.270000 0.655000 ;
      RECT 2.695000  2.085000 2.865000 2.465000 ;
      RECT 3.165000  0.425000 3.435000 0.775000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvn_2


MACRO sky130_fd_sc_hdll__einvn_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.520000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.980000 0.620000 5.415000 1.325000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.954300 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.345000 1.325000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.490000 0.620000 4.810000 1.480000 ;
        RECT 3.490000 1.480000 3.870000 2.075000 ;
        RECT 4.430000 1.480000 4.810000 2.075000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.895000 0.825000 ;
      RECT 0.085000  1.495000 0.895000 1.665000 ;
      RECT 0.085000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.895000 0.485000 ;
      RECT 0.515000  0.825000 0.895000 0.995000 ;
      RECT 0.515000  0.995000 3.320000 1.325000 ;
      RECT 0.515000  1.325000 0.895000 1.495000 ;
      RECT 0.515000  1.835000 0.895000 2.635000 ;
      RECT 1.065000  0.255000 1.385000 0.655000 ;
      RECT 1.065000  0.655000 3.295000 0.825000 ;
      RECT 1.065000  1.495000 3.320000 1.665000 ;
      RECT 1.065000  1.665000 1.340000 2.465000 ;
      RECT 1.510000  1.835000 1.890000 2.635000 ;
      RECT 1.605000  0.085000 1.935000 0.485000 ;
      RECT 2.110000  1.665000 2.280000 2.465000 ;
      RECT 2.155000  0.255000 2.325000 0.655000 ;
      RECT 2.450000  1.835000 2.890000 2.635000 ;
      RECT 2.545000  0.085000 2.875000 0.485000 ;
      RECT 3.110000  1.665000 3.320000 2.295000 ;
      RECT 3.110000  2.295000 5.200000 2.465000 ;
      RECT 3.125000  0.255000 5.435000 0.450000 ;
      RECT 3.125000  0.450000 3.295000 0.655000 ;
      RECT 4.090000  1.650000 4.260000 2.295000 ;
      RECT 5.030000  1.650000 5.200000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvn_4


MACRO sky130_fd_sc_hdll__einvn_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.200000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.145000 0.995000 8.650000 1.285000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.631100 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.345000 1.325000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.370000 0.620000 9.095000 0.825000 ;
        RECT 5.370000 1.455000 9.095000 1.625000 ;
        RECT 5.370000 1.625000 5.750000 2.125000 ;
        RECT 6.310000 1.625000 6.690000 2.125000 ;
        RECT 7.250000 1.625000 7.630000 2.125000 ;
        RECT 8.190000 1.625000 8.570000 2.125000 ;
        RECT 8.870000 0.825000 9.095000 1.455000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.090000  0.255000 0.345000 0.655000 ;
      RECT 0.090000  0.655000 0.895000 0.825000 ;
      RECT 0.090000  1.495000 0.895000 1.665000 ;
      RECT 0.090000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.895000 0.485000 ;
      RECT 0.515000  0.825000 0.895000 0.995000 ;
      RECT 0.515000  0.995000 4.975000 1.325000 ;
      RECT 0.515000  1.325000 0.895000 1.495000 ;
      RECT 0.515000  1.835000 0.895000 2.635000 ;
      RECT 1.065000  0.255000 1.385000 0.655000 ;
      RECT 1.065000  0.655000 5.200000 0.825000 ;
      RECT 1.065000  1.495000 5.200000 1.665000 ;
      RECT 1.065000  1.665000 1.340000 2.465000 ;
      RECT 1.510000  1.835000 1.890000 2.635000 ;
      RECT 1.605000  0.085000 1.935000 0.485000 ;
      RECT 2.110000  1.665000 2.280000 2.465000 ;
      RECT 2.155000  0.255000 2.325000 0.655000 ;
      RECT 2.450000  1.835000 2.830000 2.635000 ;
      RECT 2.545000  0.085000 2.875000 0.485000 ;
      RECT 3.050000  1.665000 3.220000 2.465000 ;
      RECT 3.095000  0.255000 3.265000 0.655000 ;
      RECT 3.390000  1.835000 3.770000 2.635000 ;
      RECT 3.485000  0.085000 3.815000 0.485000 ;
      RECT 3.990000  1.665000 4.160000 2.465000 ;
      RECT 4.035000  0.255000 4.205000 0.655000 ;
      RECT 4.330000  1.835000 4.730000 2.635000 ;
      RECT 4.425000  0.085000 4.765000 0.485000 ;
      RECT 4.950000  1.665000 5.200000 2.295000 ;
      RECT 4.950000  2.295000 9.095000 2.465000 ;
      RECT 4.985000  0.255000 9.095000 0.450000 ;
      RECT 4.985000  0.450000 5.200000 0.655000 ;
      RECT 5.970000  1.795000 6.140000 2.295000 ;
      RECT 6.910000  1.795000 7.080000 2.295000 ;
      RECT 7.850000  1.795000 8.020000 2.295000 ;
      RECT 8.790000  1.795000 9.095000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvn_8


MACRO sky130_fd_sc_hdll__einvn_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.430000 0.765000 2.675000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.358200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.510000 1.725000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.471500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.400000 1.785000 2.675000 2.465000 ;
        RECT 1.970000 0.255000 2.675000 0.595000 ;
        RECT 1.970000 0.595000 2.210000 1.785000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.255000 0.370000 0.615000 ;
      RECT 0.085000  0.615000 1.600000 0.785000 ;
      RECT 0.085000  1.895000 0.920000 2.065000 ;
      RECT 0.085000  2.065000 0.370000 2.465000 ;
      RECT 0.540000  0.085000 1.590000 0.445000 ;
      RECT 0.540000  2.235000 0.920000 2.635000 ;
      RECT 0.735000  0.785000 1.600000 0.805000 ;
      RECT 0.735000  1.440000 1.600000 1.615000 ;
      RECT 0.735000  1.615000 0.920000 1.895000 ;
      RECT 1.120000  0.805000 1.600000 1.440000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__einvn_1


MACRO sky130_fd_sc_hdll__clkinvlp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  1.840000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.995000 0.600000 1.665000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.436800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.785000 0.315000 1.545000 0.750000 ;
        RECT 0.785000 0.750000 1.235000 2.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.225000  1.835000 0.555000 2.625000 ;
      RECT 0.225000  2.625000 1.665000 2.635000 ;
      RECT 0.295000  0.085000 0.615000 0.745000 ;
      RECT 1.405000  1.455000 1.665000 2.625000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinvlp_2


MACRO sky130_fd_sc_hdll__clkinvlp_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.330000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.745000 0.425000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.694000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.255000 1.165000 0.680000 ;
        RECT 0.605000 0.680000 0.955000 1.015000 ;
        RECT 0.605000 1.015000 1.985000 1.295000 ;
        RECT 0.605000 1.295000 0.945000 2.465000 ;
        RECT 1.655000 1.295000 1.985000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.575000 ;
      RECT 0.095000  1.495000 0.420000 2.635000 ;
      RECT 1.185000  1.465000 1.460000 2.635000 ;
      RECT 1.675000  0.085000 2.000000 0.775000 ;
      RECT 2.225000  1.465000 2.505000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinvlp_4


MACRO sky130_fd_sc_hdll__nor3_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 2.025000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 1.075000 4.085000 1.285000 ;
        RECT 3.915000 1.285000 4.085000 1.445000 ;
        RECT 3.915000 1.445000 5.715000 1.615000 ;
        RECT 5.545000 1.075000 5.885000 1.285000 ;
        RECT 5.545000 1.285000 5.715000 1.445000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.255000 1.075000 5.315000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.828000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 6.345000 0.905000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 2.415000 0.255000 2.795000 0.725000 ;
        RECT 3.355000 0.255000 3.735000 0.725000 ;
        RECT 3.915000 1.785000 6.345000 1.955000 ;
        RECT 3.915000 1.955000 5.105000 1.965000 ;
        RECT 3.915000 1.965000 4.165000 2.125000 ;
        RECT 4.295000 0.255000 4.675000 0.725000 ;
        RECT 4.855000 1.965000 5.105000 2.125000 ;
        RECT 5.235000 0.255000 5.615000 0.725000 ;
        RECT 6.055000 0.905000 6.345000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.150000  1.455000 2.285000 1.625000 ;
      RECT 0.150000  1.625000 0.405000 2.465000 ;
      RECT 0.625000  1.795000 0.875000 2.635000 ;
      RECT 1.095000  1.625000 1.345000 2.465000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 1.565000  1.795000 1.815000 2.635000 ;
      RECT 2.035000  1.625000 2.285000 2.085000 ;
      RECT 2.035000  2.085000 3.225000 2.465000 ;
      RECT 2.075000  0.085000 2.245000 0.555000 ;
      RECT 2.505000  1.455000 3.695000 1.625000 ;
      RECT 2.505000  1.625000 2.755000 1.915000 ;
      RECT 2.975000  1.795000 3.225000 2.085000 ;
      RECT 3.015000  0.085000 3.185000 0.555000 ;
      RECT 3.445000  1.625000 3.695000 2.295000 ;
      RECT 3.445000  2.295000 5.575000 2.465000 ;
      RECT 3.955000  0.085000 4.125000 0.555000 ;
      RECT 4.385000  2.135000 4.635000 2.295000 ;
      RECT 4.895000  0.085000 5.065000 0.555000 ;
      RECT 5.325000  2.135000 5.575000 2.295000 ;
      RECT 5.795000  2.125000 6.045000 2.465000 ;
      RECT 5.835000  0.085000 6.005000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.695000  2.125000 2.865000 2.295000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.805000  2.125000 5.975000 2.295000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 2.635000 2.065000 2.980000 2.140000 ;
      RECT 2.635000 2.140000 6.040000 2.280000 ;
      RECT 2.635000 2.280000 2.980000 2.335000 ;
      RECT 5.695000 2.065000 6.040000 2.140000 ;
      RECT 5.695000 2.280000 6.040000 2.335000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3_4


MACRO sky130_fd_sc_hdll__nor3_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.740000 0.655000 2.205000 1.665000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.995000 1.075000 1.325000 ;
        RECT 0.595000 1.325000 0.880000 2.005000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.425000 1.325000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.647000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.385000 0.345000 0.655000 ;
        RECT 0.090000 0.655000 1.415000 0.825000 ;
        RECT 0.090000 1.495000 0.425000 2.280000 ;
        RECT 0.090000 2.280000 1.415000 2.450000 ;
        RECT 1.115000 0.385000 1.285000 0.655000 ;
        RECT 1.245000 0.825000 1.415000 2.280000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.515000  0.085000 0.895000 0.485000 ;
      RECT 1.455000  0.085000 2.175000 0.485000 ;
      RECT 1.585000  1.835000 2.175000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3_1


MACRO sky130_fd_sc_hdll__nor3_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 1.075000 1.015000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.235000 1.075000 2.275000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.075000 3.310000 1.285000 ;
        RECT 2.445000 1.285000 2.935000 1.625000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.011500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 3.995000 0.905000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 3.050000 0.255000 3.430000 0.725000 ;
        RECT 3.180000 1.455000 3.995000 1.625000 ;
        RECT 3.180000 1.625000 3.390000 2.125000 ;
        RECT 3.480000 0.905000 3.995000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.150000  1.455000 2.275000 1.625000 ;
      RECT 0.150000  1.625000 0.405000 2.465000 ;
      RECT 0.625000  1.795000 0.875000 2.635000 ;
      RECT 1.095000  1.625000 1.345000 2.465000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 1.565000  1.795000 1.815000 2.295000 ;
      RECT 1.565000  2.295000 3.860000 2.465000 ;
      RECT 2.035000  1.625000 2.275000 2.125000 ;
      RECT 2.075000  0.085000 2.880000 0.555000 ;
      RECT 2.710000  1.795000 2.920000 2.295000 ;
      RECT 3.610000  1.795000 3.860000 2.295000 ;
      RECT 3.650000  0.085000 3.940000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor3_2


MACRO sky130_fd_sc_hdll__isobufsrc_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.660000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.315000 1.065000 ;
        RECT 0.085000 1.065000 0.505000 1.285000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.790000 1.075000 8.880000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  2.889000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.125000 0.255000 2.505000 0.725000 ;
        RECT 2.125000 0.725000 9.565000 0.905000 ;
        RECT 3.065000 0.255000 3.445000 0.725000 ;
        RECT 4.005000 0.255000 4.385000 0.725000 ;
        RECT 4.945000 0.255000 5.325000 0.725000 ;
        RECT 5.885000 0.255000 6.265000 0.725000 ;
        RECT 5.975000 1.445000 9.565000 1.615000 ;
        RECT 5.975000 1.615000 6.225000 2.125000 ;
        RECT 6.825000 0.255000 7.205000 0.725000 ;
        RECT 6.915000 1.615000 7.165000 2.125000 ;
        RECT 7.765000 0.255000 8.145000 0.725000 ;
        RECT 7.855000 1.615000 8.105000 2.125000 ;
        RECT 8.705000 0.255000 9.085000 0.725000 ;
        RECT 8.795000 1.615000 9.045000 2.125000 ;
        RECT 9.050000 0.905000 9.565000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.125000  1.455000 0.345000 2.635000 ;
      RECT 0.485000  0.085000 0.705000 0.895000 ;
      RECT 0.515000  1.455000 0.945000 2.465000 ;
      RECT 0.725000  1.065000 1.235000 1.075000 ;
      RECT 0.725000  1.075000 5.520000 1.285000 ;
      RECT 0.725000  1.285000 0.945000 1.455000 ;
      RECT 0.875000  0.255000 1.235000 1.065000 ;
      RECT 1.165000  1.455000 1.460000 2.635000 ;
      RECT 1.445000  0.085000 1.955000 0.905000 ;
      RECT 1.675000  1.455000 5.755000 1.665000 ;
      RECT 1.675000  1.665000 1.995000 2.465000 ;
      RECT 2.215000  1.835000 2.465000 2.635000 ;
      RECT 2.685000  1.665000 2.935000 2.465000 ;
      RECT 2.725000  0.085000 2.895000 0.555000 ;
      RECT 3.155000  1.835000 3.405000 2.635000 ;
      RECT 3.625000  1.665000 3.875000 2.465000 ;
      RECT 3.665000  0.085000 3.835000 0.555000 ;
      RECT 4.095000  1.835000 4.345000 2.635000 ;
      RECT 4.565000  1.665000 4.815000 2.465000 ;
      RECT 4.605000  0.085000 4.775000 0.555000 ;
      RECT 5.035000  1.835000 5.285000 2.635000 ;
      RECT 5.505000  1.665000 5.755000 2.295000 ;
      RECT 5.505000  2.295000 9.515000 2.465000 ;
      RECT 5.545000  0.085000 5.715000 0.555000 ;
      RECT 6.445000  1.785000 6.695000 2.295000 ;
      RECT 6.485000  0.085000 6.655000 0.555000 ;
      RECT 7.385000  1.785000 7.635000 2.295000 ;
      RECT 7.425000  0.085000 7.595000 0.555000 ;
      RECT 8.325000  1.785000 8.575000 2.295000 ;
      RECT 8.365000  0.085000 8.535000 0.555000 ;
      RECT 9.265000  1.785000 9.515000 2.295000 ;
      RECT 9.305000  0.085000 9.575000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__isobufsrc_8


MACRO sky130_fd_sc_hdll__isobufsrc_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.520000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.845000 1.075000 5.425000 1.320000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.075000 1.950000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  1.477000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 3.735000 0.905000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 2.415000 0.255000 2.795000 0.725000 ;
        RECT 2.545000 0.905000 2.875000 1.445000 ;
        RECT 2.545000 1.445000 3.655000 1.745000 ;
        RECT 2.545000 1.745000 2.715000 2.125000 ;
        RECT 3.355000 0.255000 3.735000 0.725000 ;
        RECT 3.485000 1.745000 3.655000 2.125000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.905000 ;
      RECT 0.085000  1.455000 2.325000 1.665000 ;
      RECT 0.085000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.915000 2.635000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 1.135000  1.665000 1.305000 2.465000 ;
      RECT 1.475000  1.835000 1.775000 2.635000 ;
      RECT 1.945000  1.665000 2.325000 2.295000 ;
      RECT 1.945000  2.295000 4.255000 2.465000 ;
      RECT 2.075000  0.085000 2.245000 0.555000 ;
      RECT 2.885000  1.935000 3.265000 2.295000 ;
      RECT 3.015000  0.085000 3.185000 0.555000 ;
      RECT 3.095000  1.075000 4.675000 1.275000 ;
      RECT 3.825000  1.575000 4.255000 2.295000 ;
      RECT 3.955000  0.085000 4.245000 0.905000 ;
      RECT 4.425000  0.255000 4.755000 0.815000 ;
      RECT 4.425000  0.815000 4.675000 1.075000 ;
      RECT 4.425000  1.275000 4.675000 1.575000 ;
      RECT 4.425000  1.575000 4.755000 2.465000 ;
      RECT 4.975000  0.085000 5.265000 0.905000 ;
      RECT 4.975000  1.495000 5.380000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__isobufsrc_4


MACRO sky130_fd_sc_hdll__isobufsrc_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.725000 0.325000 1.325000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 1.065000 1.425000 1.325000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.478000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.285000 0.255000 1.635000 0.645000 ;
        RECT 1.285000 0.645000 2.205000 0.815000 ;
        RECT 1.755000 1.850000 2.205000 2.465000 ;
        RECT 2.025000 0.815000 2.205000 1.850000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.330000  0.370000 0.675000 0.545000 ;
      RECT 0.415000  1.510000 1.855000 1.680000 ;
      RECT 0.415000  1.680000 0.675000 1.905000 ;
      RECT 0.495000  0.545000 0.675000 1.510000 ;
      RECT 0.905000  0.085000 1.115000 0.895000 ;
      RECT 0.925000  1.855000 1.255000 2.635000 ;
      RECT 1.635000  0.985000 1.855000 1.510000 ;
      RECT 1.805000  0.085000 2.135000 0.475000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__isobufsrc_1


MACRO sky130_fd_sc_hdll__isobufsrc_16
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  18.40000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.315000 0.995000 ;
        RECT 0.085000 0.995000 0.665000 1.325000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  4.440000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.650000 1.075000 17.600000 1.285000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  5.713000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  3.325000 0.255000  3.705000 0.725000 ;
        RECT  3.325000 0.725000 18.305000 0.905000 ;
        RECT  4.265000 0.255000  4.645000 0.725000 ;
        RECT  5.205000 0.255000  5.585000 0.725000 ;
        RECT  6.145000 0.255000  6.525000 0.725000 ;
        RECT  7.085000 0.255000  7.465000 0.725000 ;
        RECT  8.025000 0.255000  8.405000 0.725000 ;
        RECT  8.965000 0.255000  9.345000 0.725000 ;
        RECT  9.905000 0.255000 10.285000 0.725000 ;
        RECT 10.845000 0.255000 11.225000 0.725000 ;
        RECT 10.935000 1.455000 18.305000 1.625000 ;
        RECT 10.935000 1.625000 11.185000 2.125000 ;
        RECT 11.785000 0.255000 12.165000 0.725000 ;
        RECT 11.875000 1.625000 12.125000 2.125000 ;
        RECT 12.725000 0.255000 13.105000 0.725000 ;
        RECT 12.815000 1.625000 13.065000 2.125000 ;
        RECT 13.665000 0.255000 14.045000 0.725000 ;
        RECT 13.755000 1.625000 14.005000 2.125000 ;
        RECT 14.605000 0.255000 14.985000 0.725000 ;
        RECT 14.695000 1.625000 14.945000 2.125000 ;
        RECT 15.545000 0.255000 15.925000 0.725000 ;
        RECT 15.635000 1.625000 15.885000 2.125000 ;
        RECT 16.485000 0.255000 16.865000 0.725000 ;
        RECT 16.575000 1.625000 16.825000 2.125000 ;
        RECT 17.425000 0.255000 17.805000 0.725000 ;
        RECT 17.515000 1.625000 17.765000 2.125000 ;
        RECT 17.770000 0.905000 18.305000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 18.400000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 18.400000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 18.400000 0.085000 ;
      RECT  0.000000  2.635000 18.400000 2.805000 ;
      RECT  0.300000  1.495000  0.515000 2.635000 ;
      RECT  0.485000  0.085000  0.865000 0.825000 ;
      RECT  0.685000  1.495000  1.115000 2.465000 ;
      RECT  0.885000  1.065000  2.385000 1.075000 ;
      RECT  0.885000  1.075000 10.480000 1.285000 ;
      RECT  0.885000  1.285000  1.115000 1.495000 ;
      RECT  1.085000  0.255000  1.345000 1.065000 ;
      RECT  1.335000  1.455000  1.555000 2.635000 ;
      RECT  1.565000  0.085000  1.865000 0.895000 ;
      RECT  1.725000  1.285000  2.155000 2.465000 ;
      RECT  2.085000  0.255000  2.385000 1.065000 ;
      RECT  2.375000  1.455000  2.670000 2.635000 ;
      RECT  2.605000  0.085000  3.155000 0.905000 ;
      RECT  2.875000  1.455000 10.715000 1.665000 ;
      RECT  2.875000  1.665000  3.195000 2.465000 ;
      RECT  3.415000  1.835000  3.665000 2.635000 ;
      RECT  3.885000  1.665000  4.135000 2.465000 ;
      RECT  3.925000  0.085000  4.095000 0.555000 ;
      RECT  4.355000  1.835000  4.605000 2.635000 ;
      RECT  4.825000  1.665000  5.075000 2.465000 ;
      RECT  4.865000  0.085000  5.035000 0.555000 ;
      RECT  5.295000  1.835000  5.545000 2.635000 ;
      RECT  5.765000  1.665000  6.015000 2.465000 ;
      RECT  5.805000  0.085000  5.975000 0.555000 ;
      RECT  6.235000  1.835000  6.485000 2.635000 ;
      RECT  6.705000  1.665000  6.955000 2.465000 ;
      RECT  6.745000  0.085000  6.915000 0.555000 ;
      RECT  7.175000  1.835000  7.425000 2.635000 ;
      RECT  7.645000  1.665000  7.895000 2.465000 ;
      RECT  7.685000  0.085000  7.855000 0.555000 ;
      RECT  8.115000  1.835000  8.365000 2.635000 ;
      RECT  8.585000  1.665000  8.835000 2.465000 ;
      RECT  8.625000  0.085000  8.795000 0.555000 ;
      RECT  9.055000  1.835000  9.305000 2.635000 ;
      RECT  9.525000  1.665000  9.775000 2.465000 ;
      RECT  9.565000  0.085000  9.735000 0.555000 ;
      RECT  9.995000  1.835000 10.245000 2.635000 ;
      RECT 10.465000  1.665000 10.715000 2.295000 ;
      RECT 10.465000  2.295000 18.235000 2.465000 ;
      RECT 10.505000  0.085000 10.675000 0.555000 ;
      RECT 11.405000  1.795000 11.655000 2.295000 ;
      RECT 11.445000  0.085000 11.615000 0.555000 ;
      RECT 12.345000  1.795000 12.595000 2.295000 ;
      RECT 12.385000  0.085000 12.555000 0.555000 ;
      RECT 13.285000  1.795000 13.535000 2.295000 ;
      RECT 13.325000  0.085000 13.495000 0.555000 ;
      RECT 14.225000  1.795000 14.475000 2.295000 ;
      RECT 14.265000  0.085000 14.435000 0.555000 ;
      RECT 15.165000  1.795000 15.415000 2.295000 ;
      RECT 15.205000  0.085000 15.375000 0.555000 ;
      RECT 16.105000  1.795000 16.355000 2.295000 ;
      RECT 16.145000  0.085000 16.315000 0.555000 ;
      RECT 17.045000  1.795000 17.295000 2.295000 ;
      RECT 17.085000  0.085000 17.255000 0.555000 ;
      RECT 17.985000  1.795000 18.235000 2.295000 ;
      RECT 18.025000  0.085000 18.295000 0.555000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
      RECT 17.165000 -0.085000 17.335000 0.085000 ;
      RECT 17.165000  2.635000 17.335000 2.805000 ;
      RECT 17.625000 -0.085000 17.795000 0.085000 ;
      RECT 17.625000  2.635000 17.795000 2.805000 ;
      RECT 18.085000 -0.085000 18.255000 0.085000 ;
      RECT 18.085000  2.635000 18.255000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__isobufsrc_16


MACRO sky130_fd_sc_hdll__isobufsrc_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.800000 1.065000 3.555000 1.275000 ;
        RECT 3.340000 1.275000 3.555000 1.965000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.480000 1.065000 0.970000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.771000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 1.855000 0.895000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 1.525000 0.895000 1.815000 2.125000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.895000 ;
      RECT 0.085000  1.445000 1.345000 1.655000 ;
      RECT 0.085000  1.655000 0.405000 2.465000 ;
      RECT 0.625000  1.825000 0.875000 2.635000 ;
      RECT 1.095000  1.655000 1.345000 2.295000 ;
      RECT 1.095000  2.295000 2.325000 2.465000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 2.035000  1.445000 2.290000 1.890000 ;
      RECT 2.035000  1.890000 2.325000 2.295000 ;
      RECT 2.075000  0.085000 2.245000 0.895000 ;
      RECT 2.075000  1.075000 2.630000 1.245000 ;
      RECT 2.415000  0.725000 2.765000 0.895000 ;
      RECT 2.415000  0.895000 2.630000 1.075000 ;
      RECT 2.460000  1.245000 2.630000 1.445000 ;
      RECT 2.460000  1.445000 2.765000 1.615000 ;
      RECT 2.595000  0.445000 2.765000 0.725000 ;
      RECT 2.595000  1.615000 2.765000 2.460000 ;
      RECT 3.025000  0.085000 3.280000 0.845000 ;
      RECT 3.025000  2.145000 3.275000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__isobufsrc_2


MACRO sky130_fd_sc_hdll__fill_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE SPACER ;
  SYMMETRY X Y R90 ;
  SIZE  0.460000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__fill_1


MACRO sky130_fd_sc_hdll__fill_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE SPACER ;
  SYMMETRY X Y R90 ;
  SIZE  1.840000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__fill_4


MACRO sky130_fd_sc_hdll__fill_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE SPACER ;
  SYMMETRY X Y R90 ;
  SIZE  0.920000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.920000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.920000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.920000 0.085000 ;
      RECT 0.000000  2.635000 0.920000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__fill_2


MACRO sky130_fd_sc_hdll__fill_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE SPACER ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__fill_8


MACRO sky130_fd_sc_hdll__sdfstp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  13.34000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155000 1.055000 3.815000 1.650000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 0.765000 1.485000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.915000 0.275000 13.240000 2.450000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.467400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.580000 1.075000 0.870000 1.120000 ;
        RECT 0.580000 1.120000 2.875000 1.260000 ;
        RECT 0.580000 1.260000 0.870000 1.305000 ;
        RECT 2.585000 1.075000 2.875000 1.120000 ;
        RECT 2.585000 1.260000 2.875000 1.305000 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.375000 1.415000 7.715000 1.460000 ;
        RECT 7.375000 1.460000 9.905000 1.600000 ;
        RECT 7.375000 1.600000 7.715000 1.645000 ;
        RECT 9.565000 1.415000 9.905000 1.460000 ;
        RECT 9.565000 1.600000 9.905000 1.645000 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.340000 0.085000 ;
      RECT  0.000000  2.635000 13.340000 2.805000 ;
      RECT  0.085000  0.085000  0.750000 0.595000 ;
      RECT  0.085000  1.845000  1.225000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.835000 2.635000 ;
      RECT  0.540000  0.765000  0.870000 1.675000 ;
      RECT  0.920000  0.255000  1.845000 0.595000 ;
      RECT  1.055000  2.025000  1.225000 2.255000 ;
      RECT  1.055000  2.255000  2.245000 2.465000 ;
      RECT  1.395000  1.845000  1.845000 2.085000 ;
      RECT  1.655000  0.595000  1.845000 1.845000 ;
      RECT  2.025000  0.085000  2.290000 0.545000 ;
      RECT  2.065000  0.715000  2.720000 0.905000 ;
      RECT  2.065000  0.905000  2.400000 1.770000 ;
      RECT  2.065000  1.770000  2.720000 2.085000 ;
      RECT  2.460000  0.255000  2.720000 0.715000 ;
      RECT  2.470000  2.085000  2.720000 2.465000 ;
      RECT  2.570000  1.075000  2.950000 1.600000 ;
      RECT  2.940000  0.085000  3.350000 0.555000 ;
      RECT  2.940000  2.140000  3.235000 2.635000 ;
      RECT  3.505000  1.830000  4.295000 2.000000 ;
      RECT  3.505000  2.000000  3.675000 2.325000 ;
      RECT  3.520000  0.255000  3.705000 0.715000 ;
      RECT  3.520000  0.715000  4.295000 0.885000 ;
      RECT  3.845000  2.275000  4.225000 2.635000 ;
      RECT  3.925000  0.085000  4.255000 0.545000 ;
      RECT  4.035000  0.885000  4.295000 1.830000 ;
      RECT  4.445000  2.135000  4.790000 2.465000 ;
      RECT  4.475000  0.255000  4.685000 1.085000 ;
      RECT  4.475000  1.085000  4.840000 1.420000 ;
      RECT  4.475000  1.420000  4.790000 2.135000 ;
      RECT  4.855000  0.255000  5.180000 0.780000 ;
      RECT  4.965000  1.590000  5.180000 2.465000 ;
      RECT  5.010000  0.780000  5.180000 1.590000 ;
      RECT  5.435000  2.135000  6.205000 2.465000 ;
      RECT  5.465000  0.255000  5.890000 1.225000 ;
      RECT  5.465000  1.225000  8.315000 1.275000 ;
      RECT  5.465000  1.275000  6.975000 1.395000 ;
      RECT  5.605000  1.575000  5.865000 1.955000 ;
      RECT  6.035000  1.395000  6.205000 2.135000 ;
      RECT  6.060000  0.085000  6.595000 0.465000 ;
      RECT  6.095000  0.635000  7.035000 0.805000 ;
      RECT  6.095000  0.805000  6.475000 1.015000 ;
      RECT  6.425000  1.575000  6.595000 1.935000 ;
      RECT  6.425000  1.935000  7.420000 2.105000 ;
      RECT  6.445000  2.275000  6.830000 2.635000 ;
      RECT  6.785000  0.255000  7.035000 0.635000 ;
      RECT  6.805000  0.975000  8.315000 1.225000 ;
      RECT  7.155000  2.105000  7.420000 2.450000 ;
      RECT  7.190000  1.445000  7.715000 1.765000 ;
      RECT  7.255000  0.085000  8.315000 0.805000 ;
      RECT  7.710000  2.125000  8.625000 2.635000 ;
      RECT  7.885000  1.670000  8.785000 1.955000 ;
      RECT  7.905000  1.275000  8.315000 1.325000 ;
      RECT  8.485000  0.720000  9.850000 0.905000 ;
      RECT  8.485000  0.905000  8.785000 1.670000 ;
      RECT  8.795000  2.125000  9.690000 2.460000 ;
      RECT  8.955000  1.075000  9.290000 1.905000 ;
      RECT  9.025000  0.275000 10.650000 0.545000 ;
      RECT  9.520000  0.905000  9.850000 1.255000 ;
      RECT  9.520000  1.895000 11.255000 2.065000 ;
      RECT  9.520000  2.065000  9.690000 2.125000 ;
      RECT  9.580000  1.425000  9.860000 1.545000 ;
      RECT  9.580000  1.545000 10.695000 1.725000 ;
      RECT  9.860000  2.235000 10.190000 2.635000 ;
      RECT 10.035000  0.855000 10.280000 1.195000 ;
      RECT 10.035000  1.195000 11.685000 1.365000 ;
      RECT 10.395000  2.065000 10.595000 2.450000 ;
      RECT 10.450000  0.545000 10.650000 0.785000 ;
      RECT 10.450000  0.785000 11.285000 1.015000 ;
      RECT 10.835000  0.085000 11.085000 0.545000 ;
      RECT 10.875000  1.605000 11.255000 1.895000 ;
      RECT 10.875000  2.235000 11.255000 2.635000 ;
      RECT 11.345000  0.255000 11.685000 0.585000 ;
      RECT 11.425000  1.365000 11.685000 2.465000 ;
      RECT 11.455000  0.585000 11.685000 1.195000 ;
      RECT 11.855000  0.255000 12.115000 0.995000 ;
      RECT 11.855000  0.995000 12.745000 1.325000 ;
      RECT 11.855000  1.325000 12.195000 2.465000 ;
      RECT 12.285000  0.085000 12.690000 0.550000 ;
      RECT 12.435000  1.845000 12.690000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.640000  1.105000  0.810000 1.275000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.675000  1.445000  1.845000 1.615000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.645000  1.105000  2.815000 1.275000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.125000  1.785000  4.295000 1.955000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.635000  1.100000  4.805000 1.270000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.010000  1.445000  5.180000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.605000  1.785000  5.775000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.435000  1.445000  7.605000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.210000  1.785000  8.380000 1.955000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.050000  1.105000  9.220000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.625000  1.445000  9.795000 1.615000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
    LAYER met1 ;
      RECT 1.615000 1.415000 1.955000 1.460000 ;
      RECT 1.615000 1.460000 5.240000 1.600000 ;
      RECT 1.615000 1.600000 1.955000 1.645000 ;
      RECT 4.065000 1.755000 4.405000 1.800000 ;
      RECT 4.065000 1.800000 8.490000 1.940000 ;
      RECT 4.065000 1.940000 4.405000 1.985000 ;
      RECT 4.575000 1.070000 4.865000 1.120000 ;
      RECT 4.575000 1.120000 9.330000 1.260000 ;
      RECT 4.575000 1.260000 4.865000 1.300000 ;
      RECT 4.950000 1.415000 5.240000 1.460000 ;
      RECT 4.950000 1.600000 5.240000 1.645000 ;
      RECT 5.545000 1.755000 5.885000 1.800000 ;
      RECT 5.545000 1.940000 5.885000 1.985000 ;
      RECT 8.150000 1.755000 8.490000 1.800000 ;
      RECT 8.150000 1.940000 8.490000 1.985000 ;
      RECT 8.940000 1.075000 9.330000 1.120000 ;
      RECT 8.940000 1.260000 9.330000 1.305000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfstp_1


MACRO sky130_fd_sc_hdll__sdfstp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  14.26000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155000 1.055000 3.815000 1.650000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 0.765000 1.485000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.245000 0.275000 13.655000 0.825000 ;
        RECT 13.245000 1.495000 13.655000 2.450000 ;
        RECT 13.350000 0.825000 13.655000 1.495000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.467400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.580000 1.075000 0.870000 1.120000 ;
        RECT 0.580000 1.120000 2.875000 1.260000 ;
        RECT 0.580000 1.260000 0.870000 1.305000 ;
        RECT 2.585000 1.075000 2.875000 1.120000 ;
        RECT 2.585000 1.260000 2.875000 1.305000 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.375000 1.415000  7.715000 1.460000 ;
        RECT 7.375000 1.460000 10.070000 1.600000 ;
        RECT 7.375000 1.600000  7.715000 1.645000 ;
        RECT 9.730000 1.415000 10.070000 1.460000 ;
        RECT 9.730000 1.600000 10.070000 1.645000 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.085000  0.085000  0.750000 0.595000 ;
      RECT  0.085000  1.845000  1.225000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.835000 2.635000 ;
      RECT  0.540000  0.765000  0.870000 1.675000 ;
      RECT  0.920000  0.255000  1.845000 0.595000 ;
      RECT  1.055000  2.025000  1.225000 2.255000 ;
      RECT  1.055000  2.255000  2.245000 2.465000 ;
      RECT  1.395000  1.845000  1.845000 2.085000 ;
      RECT  1.655000  0.595000  1.845000 1.845000 ;
      RECT  2.025000  0.085000  2.290000 0.545000 ;
      RECT  2.065000  0.715000  2.720000 0.905000 ;
      RECT  2.065000  0.905000  2.400000 1.770000 ;
      RECT  2.065000  1.770000  2.720000 2.085000 ;
      RECT  2.460000  0.255000  2.720000 0.715000 ;
      RECT  2.470000  2.085000  2.720000 2.465000 ;
      RECT  2.570000  1.075000  2.950000 1.600000 ;
      RECT  2.940000  0.085000  3.350000 0.555000 ;
      RECT  2.940000  2.140000  3.235000 2.635000 ;
      RECT  3.505000  1.830000  4.295000 2.000000 ;
      RECT  3.505000  2.000000  3.675000 2.325000 ;
      RECT  3.520000  0.255000  3.705000 0.715000 ;
      RECT  3.520000  0.715000  4.295000 0.885000 ;
      RECT  3.845000  2.275000  4.225000 2.635000 ;
      RECT  3.925000  0.085000  4.255000 0.545000 ;
      RECT  4.035000  0.885000  4.295000 1.830000 ;
      RECT  4.445000  2.135000  4.790000 2.465000 ;
      RECT  4.475000  0.255000  4.685000 1.085000 ;
      RECT  4.475000  1.085000  4.840000 1.420000 ;
      RECT  4.475000  1.420000  4.790000 2.135000 ;
      RECT  4.855000  0.255000  5.180000 0.780000 ;
      RECT  4.965000  1.590000  5.180000 2.465000 ;
      RECT  5.010000  0.780000  5.180000 1.590000 ;
      RECT  5.435000  2.135000  6.205000 2.465000 ;
      RECT  5.465000  0.255000  5.890000 1.225000 ;
      RECT  5.465000  1.225000  8.415000 1.275000 ;
      RECT  5.465000  1.275000  6.975000 1.395000 ;
      RECT  5.605000  1.575000  5.865000 1.955000 ;
      RECT  6.035000  1.395000  6.205000 2.135000 ;
      RECT  6.060000  0.085000  6.595000 0.465000 ;
      RECT  6.095000  0.635000  7.035000 0.805000 ;
      RECT  6.095000  0.805000  6.475000 1.015000 ;
      RECT  6.425000  1.575000  6.595000 1.935000 ;
      RECT  6.425000  1.935000  7.420000 2.105000 ;
      RECT  6.445000  2.275000  6.830000 2.635000 ;
      RECT  6.785000  0.255000  7.035000 0.635000 ;
      RECT  6.805000  0.975000  8.415000 1.225000 ;
      RECT  7.155000  2.105000  7.420000 2.450000 ;
      RECT  7.190000  1.445000  7.715000 1.765000 ;
      RECT  7.255000  0.085000  8.415000 0.805000 ;
      RECT  7.710000  2.125000  8.765000 2.635000 ;
      RECT  7.885000  1.670000  8.885000 1.955000 ;
      RECT  8.005000  1.275000  8.415000 1.325000 ;
      RECT  8.585000  0.720000 10.005000 0.905000 ;
      RECT  8.585000  0.905000  8.885000 1.670000 ;
      RECT  8.935000  2.125000  9.840000 2.460000 ;
      RECT  9.175000  1.075000  9.500000 1.905000 ;
      RECT  9.265000  0.275000 10.910000 0.545000 ;
      RECT  9.670000  0.905000 10.005000 1.255000 ;
      RECT  9.670000  1.895000 11.585000 2.065000 ;
      RECT  9.670000  2.065000  9.840000 2.125000 ;
      RECT  9.730000  1.425000 10.035000 1.545000 ;
      RECT  9.730000  1.545000 10.995000 1.725000 ;
      RECT 10.060000  2.235000 10.440000 2.635000 ;
      RECT 10.220000  0.855000 10.480000 1.195000 ;
      RECT 10.220000  1.195000 12.015000 1.365000 ;
      RECT 10.610000  2.065000 11.015000 2.450000 ;
      RECT 10.710000  0.545000 10.910000 0.785000 ;
      RECT 10.710000  0.785000 11.615000 1.015000 ;
      RECT 11.165000  0.085000 11.415000 0.545000 ;
      RECT 11.205000  1.605000 11.585000 1.895000 ;
      RECT 11.205000  2.235000 11.585000 2.635000 ;
      RECT 11.675000  0.255000 12.015000 0.585000 ;
      RECT 11.755000  1.365000 12.015000 2.465000 ;
      RECT 11.785000  0.585000 12.015000 1.195000 ;
      RECT 12.185000  0.255000 12.445000 0.995000 ;
      RECT 12.185000  0.995000 13.125000 1.325000 ;
      RECT 12.185000  1.325000 12.525000 2.465000 ;
      RECT 12.615000  0.085000 13.020000 0.550000 ;
      RECT 12.765000  1.845000 13.020000 2.635000 ;
      RECT 13.825000  0.085000 13.995000 0.885000 ;
      RECT 13.825000  1.495000 13.995000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.640000  1.105000  0.810000 1.275000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.675000  1.445000  1.845000 1.615000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.645000  1.105000  2.815000 1.275000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.125000  1.785000  4.295000 1.955000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.635000  1.100000  4.805000 1.270000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.010000  1.445000  5.180000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.605000  1.785000  5.775000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.435000  1.445000  7.605000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.210000  1.785000  8.380000 1.955000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.280000  1.105000  9.450000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.790000  1.445000  9.960000 1.615000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT 1.615000 1.415000 1.955000 1.460000 ;
      RECT 1.615000 1.460000 5.240000 1.600000 ;
      RECT 1.615000 1.600000 1.955000 1.645000 ;
      RECT 4.065000 1.755000 4.405000 1.800000 ;
      RECT 4.065000 1.800000 8.490000 1.940000 ;
      RECT 4.065000 1.940000 4.405000 1.985000 ;
      RECT 4.575000 1.070000 4.865000 1.120000 ;
      RECT 4.575000 1.120000 9.560000 1.260000 ;
      RECT 4.575000 1.260000 4.865000 1.300000 ;
      RECT 4.950000 1.415000 5.240000 1.460000 ;
      RECT 4.950000 1.600000 5.240000 1.645000 ;
      RECT 5.545000 1.755000 5.885000 1.800000 ;
      RECT 5.545000 1.940000 5.885000 1.985000 ;
      RECT 8.150000 1.755000 8.490000 1.800000 ;
      RECT 8.150000 1.940000 8.490000 1.985000 ;
      RECT 9.170000 1.075000 9.560000 1.120000 ;
      RECT 9.170000 1.260000 9.560000 1.305000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfstp_2


MACRO sky130_fd_sc_hdll__sdfstp_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  15.18000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155000 1.055000 3.815000 1.650000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 0.765000 1.485000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.240000 0.275000 13.570000 0.825000 ;
        RECT 13.240000 1.495000 13.570000 2.450000 ;
        RECT 13.345000 0.825000 13.570000 1.055000 ;
        RECT 13.345000 1.055000 14.610000 1.325000 ;
        RECT 13.345000 1.325000 13.570000 1.495000 ;
        RECT 14.130000 0.255000 14.610000 1.055000 ;
        RECT 14.130000 1.325000 14.610000 2.465000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.467400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.580000 1.075000 0.870000 1.120000 ;
        RECT 0.580000 1.120000 2.875000 1.260000 ;
        RECT 0.580000 1.260000 0.870000 1.305000 ;
        RECT 2.585000 1.075000 2.875000 1.120000 ;
        RECT 2.585000 1.260000 2.875000 1.305000 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.375000 1.415000  7.715000 1.460000 ;
        RECT 7.375000 1.460000 10.070000 1.600000 ;
        RECT 7.375000 1.600000  7.715000 1.645000 ;
        RECT 9.730000 1.415000 10.070000 1.460000 ;
        RECT 9.730000 1.600000 10.070000 1.645000 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.180000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 15.180000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.180000 0.085000 ;
      RECT  0.000000  2.635000 15.180000 2.805000 ;
      RECT  0.085000  0.085000  0.750000 0.595000 ;
      RECT  0.085000  1.845000  1.225000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.835000 2.635000 ;
      RECT  0.540000  0.765000  0.870000 1.675000 ;
      RECT  0.920000  0.255000  1.845000 0.595000 ;
      RECT  1.055000  2.025000  1.225000 2.255000 ;
      RECT  1.055000  2.255000  2.245000 2.465000 ;
      RECT  1.395000  1.845000  1.845000 2.085000 ;
      RECT  1.655000  0.595000  1.845000 1.845000 ;
      RECT  2.025000  0.085000  2.290000 0.545000 ;
      RECT  2.065000  0.715000  2.720000 0.905000 ;
      RECT  2.065000  0.905000  2.400000 1.770000 ;
      RECT  2.065000  1.770000  2.720000 2.085000 ;
      RECT  2.460000  0.255000  2.720000 0.715000 ;
      RECT  2.470000  2.085000  2.720000 2.465000 ;
      RECT  2.570000  1.075000  2.950000 1.600000 ;
      RECT  2.940000  0.085000  3.350000 0.555000 ;
      RECT  2.940000  2.140000  3.235000 2.635000 ;
      RECT  3.505000  1.830000  4.295000 2.000000 ;
      RECT  3.505000  2.000000  3.675000 2.325000 ;
      RECT  3.520000  0.255000  3.705000 0.715000 ;
      RECT  3.520000  0.715000  4.295000 0.885000 ;
      RECT  3.845000  2.275000  4.225000 2.635000 ;
      RECT  3.925000  0.085000  4.255000 0.545000 ;
      RECT  4.035000  0.885000  4.295000 1.830000 ;
      RECT  4.445000  2.135000  4.790000 2.465000 ;
      RECT  4.475000  0.255000  4.685000 1.085000 ;
      RECT  4.475000  1.085000  4.840000 1.420000 ;
      RECT  4.475000  1.420000  4.790000 2.135000 ;
      RECT  4.855000  0.255000  5.180000 0.780000 ;
      RECT  4.965000  1.590000  5.180000 2.465000 ;
      RECT  5.010000  0.780000  5.180000 1.590000 ;
      RECT  5.435000  2.135000  6.205000 2.465000 ;
      RECT  5.465000  0.255000  5.890000 1.225000 ;
      RECT  5.465000  1.225000  8.415000 1.275000 ;
      RECT  5.465000  1.275000  6.975000 1.395000 ;
      RECT  5.605000  1.575000  5.865000 1.955000 ;
      RECT  6.035000  1.395000  6.205000 2.135000 ;
      RECT  6.060000  0.085000  6.595000 0.465000 ;
      RECT  6.095000  0.635000  7.035000 0.805000 ;
      RECT  6.095000  0.805000  6.475000 1.015000 ;
      RECT  6.425000  1.575000  6.595000 1.935000 ;
      RECT  6.425000  1.935000  7.420000 2.105000 ;
      RECT  6.445000  2.275000  6.830000 2.635000 ;
      RECT  6.785000  0.255000  7.035000 0.635000 ;
      RECT  6.805000  0.975000  8.415000 1.225000 ;
      RECT  7.155000  2.105000  7.420000 2.450000 ;
      RECT  7.190000  1.445000  7.715000 1.765000 ;
      RECT  7.255000  0.085000  8.415000 0.805000 ;
      RECT  7.710000  2.125000  8.765000 2.635000 ;
      RECT  7.885000  1.670000  8.885000 1.955000 ;
      RECT  8.005000  1.275000  8.415000 1.325000 ;
      RECT  8.585000  0.720000 10.005000 0.905000 ;
      RECT  8.585000  0.905000  8.885000 1.670000 ;
      RECT  8.935000  2.125000  9.840000 2.460000 ;
      RECT  9.175000  1.075000  9.500000 1.905000 ;
      RECT  9.265000  0.275000 10.910000 0.545000 ;
      RECT  9.670000  0.905000 10.005000 1.255000 ;
      RECT  9.670000  1.895000 11.585000 2.065000 ;
      RECT  9.670000  2.065000  9.840000 2.125000 ;
      RECT  9.730000  1.425000 10.035000 1.545000 ;
      RECT  9.730000  1.545000 10.995000 1.725000 ;
      RECT 10.060000  2.235000 10.440000 2.635000 ;
      RECT 10.220000  0.855000 10.480000 1.195000 ;
      RECT 10.220000  1.195000 12.015000 1.365000 ;
      RECT 10.610000  2.065000 11.015000 2.450000 ;
      RECT 10.710000  0.545000 10.910000 0.785000 ;
      RECT 10.710000  0.785000 11.615000 1.015000 ;
      RECT 11.165000  0.085000 11.415000 0.545000 ;
      RECT 11.205000  1.605000 11.585000 1.895000 ;
      RECT 11.205000  2.235000 11.585000 2.635000 ;
      RECT 11.675000  0.255000 12.015000 0.585000 ;
      RECT 11.755000  1.365000 12.015000 2.465000 ;
      RECT 11.785000  0.585000 12.015000 1.195000 ;
      RECT 12.185000  0.255000 12.445000 0.995000 ;
      RECT 12.185000  0.995000 13.125000 1.325000 ;
      RECT 12.185000  1.325000 12.445000 2.465000 ;
      RECT 12.615000  0.085000 13.020000 0.825000 ;
      RECT 12.615000  1.495000 13.020000 2.635000 ;
      RECT 13.790000  0.085000 13.960000 0.885000 ;
      RECT 13.790000  1.495000 13.960000 2.635000 ;
      RECT 14.780000  0.085000 15.065000 0.885000 ;
      RECT 14.780000  1.495000 15.065000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.640000  1.105000  0.810000 1.275000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.675000  1.445000  1.845000 1.615000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.645000  1.105000  2.815000 1.275000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.125000  1.785000  4.295000 1.955000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.635000  1.100000  4.805000 1.270000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.010000  1.445000  5.180000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.605000  1.785000  5.775000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.435000  1.445000  7.605000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.210000  1.785000  8.380000 1.955000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.280000  1.105000  9.450000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.790000  1.445000  9.960000 1.615000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
    LAYER met1 ;
      RECT 1.615000 1.415000 1.955000 1.460000 ;
      RECT 1.615000 1.460000 5.240000 1.600000 ;
      RECT 1.615000 1.600000 1.955000 1.645000 ;
      RECT 4.065000 1.755000 4.405000 1.800000 ;
      RECT 4.065000 1.800000 8.490000 1.940000 ;
      RECT 4.065000 1.940000 4.405000 1.985000 ;
      RECT 4.575000 1.070000 4.865000 1.120000 ;
      RECT 4.575000 1.120000 9.560000 1.260000 ;
      RECT 4.575000 1.260000 4.865000 1.300000 ;
      RECT 4.950000 1.415000 5.240000 1.460000 ;
      RECT 4.950000 1.600000 5.240000 1.645000 ;
      RECT 5.545000 1.755000 5.885000 1.800000 ;
      RECT 5.545000 1.940000 5.885000 1.985000 ;
      RECT 8.150000 1.755000 8.490000 1.800000 ;
      RECT 8.150000 1.940000 8.490000 1.985000 ;
      RECT 9.170000 1.075000 9.560000 1.120000 ;
      RECT 9.170000 1.260000 9.560000 1.305000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfstp_4


MACRO sky130_fd_sc_hdll__a21o_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.340000 1.010000 4.965000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.010000 4.170000 1.275000 ;
        RECT 3.945000 1.275000 4.170000 1.510000 ;
        RECT 3.945000 1.510000 5.435000 1.680000 ;
        RECT 5.135000 1.055000 5.600000 1.290000 ;
        RECT 5.135000 1.290000 5.435000 1.510000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.500000 0.995000 2.905000 1.525000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.029000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.615000 1.885000 0.785000 ;
        RECT 0.145000 0.785000 0.680000 1.585000 ;
        RECT 0.145000 1.585000 1.885000 1.755000 ;
        RECT 0.675000 1.755000 0.845000 2.185000 ;
        RECT 1.635000 1.755000 1.885000 2.185000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.105000  0.085000 0.445000 0.445000 ;
      RECT 0.115000  1.935000 0.445000 2.635000 ;
      RECT 0.850000  0.995000 2.300000 1.325000 ;
      RECT 1.025000  0.085000 1.405000 0.445000 ;
      RECT 1.025000  1.935000 1.405000 2.635000 ;
      RECT 2.065000  1.515000 2.315000 2.635000 ;
      RECT 2.110000  0.085000 2.885000 0.445000 ;
      RECT 2.130000  0.615000 3.295000 0.670000 ;
      RECT 2.130000  0.670000 4.765000 0.785000 ;
      RECT 2.130000  0.785000 2.300000 0.995000 ;
      RECT 2.655000  1.695000 2.825000 2.295000 ;
      RECT 2.655000  2.295000 3.765000 2.465000 ;
      RECT 3.125000  0.255000 3.295000 0.615000 ;
      RECT 3.125000  0.785000 4.765000 0.840000 ;
      RECT 3.125000  0.840000 3.295000 2.125000 ;
      RECT 3.555000  0.085000 3.885000 0.445000 ;
      RECT 3.585000  1.445000 3.765000 1.850000 ;
      RECT 3.585000  1.850000 5.860000 2.020000 ;
      RECT 3.585000  2.020000 3.765000 2.295000 ;
      RECT 3.935000  2.275000 4.315000 2.635000 ;
      RECT 4.485000  0.405000 4.765000 0.670000 ;
      RECT 4.535000  2.020000 4.705000 2.465000 ;
      RECT 4.875000  2.275000 5.255000 2.635000 ;
      RECT 5.445000  0.085000 5.725000 0.885000 ;
      RECT 5.530000  2.020000 5.860000 2.395000 ;
      RECT 5.605000  1.460000 5.860000 1.850000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_4


MACRO sky130_fd_sc_hdll__a21o_6
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.900000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 1.055000 1.535000 1.290000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.055000 0.695000 1.290000 ;
        RECT 0.525000 1.290000 0.695000 1.460000 ;
        RECT 0.525000 1.460000 1.875000 1.630000 ;
        RECT 1.705000 1.055000 2.045000 1.290000 ;
        RECT 1.705000 1.290000 1.875000 1.460000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 1.055000 3.195000 1.615000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.396500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.905000 0.255000 4.235000 0.695000 ;
        RECT 3.905000 0.695000 6.115000 0.865000 ;
        RECT 3.935000 1.445000 6.085000 1.615000 ;
        RECT 3.935000 1.615000 4.205000 2.465000 ;
        RECT 4.845000 0.255000 5.175000 0.695000 ;
        RECT 4.875000 1.615000 5.145000 2.465000 ;
        RECT 5.625000 0.865000 5.875000 1.445000 ;
        RECT 5.785000 0.255000 6.115000 0.695000 ;
        RECT 5.815000 1.615000 6.085000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.095000  1.460000 0.355000 1.800000 ;
      RECT 0.095000  1.800000 2.275000 1.970000 ;
      RECT 0.095000  1.970000 0.425000 2.465000 ;
      RECT 0.205000  0.085000 0.535000 0.885000 ;
      RECT 0.595000  2.140000 0.865000 2.635000 ;
      RECT 1.035000  0.275000 1.365000 0.675000 ;
      RECT 1.035000  0.675000 3.735000 0.885000 ;
      RECT 1.035000  1.970000 1.365000 2.465000 ;
      RECT 1.535000  2.140000 1.805000 2.635000 ;
      RECT 1.945000  0.085000 2.275000 0.505000 ;
      RECT 1.975000  1.970000 2.275000 2.295000 ;
      RECT 1.975000  2.295000 3.245000 2.465000 ;
      RECT 2.045000  1.460000 2.275000 1.800000 ;
      RECT 2.445000  0.255000 2.745000 0.675000 ;
      RECT 2.445000  0.885000 2.695000 1.790000 ;
      RECT 2.445000  1.790000 2.745000 2.125000 ;
      RECT 2.915000  0.085000 3.735000 0.505000 ;
      RECT 2.915000  1.785000 3.245000 2.295000 ;
      RECT 3.485000  1.495000 3.735000 2.635000 ;
      RECT 3.565000  0.885000 3.735000 1.035000 ;
      RECT 3.565000  1.035000 5.455000 1.275000 ;
      RECT 4.375000  1.785000 4.705000 2.635000 ;
      RECT 4.405000  0.085000 4.675000 0.525000 ;
      RECT 5.315000  1.785000 5.645000 2.635000 ;
      RECT 5.345000  0.085000 5.615000 0.525000 ;
      RECT 6.265000  1.445000 6.595000 2.635000 ;
      RECT 6.285000  0.085000 6.535000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_6


MACRO sky130_fd_sc_hdll__a21o_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.410000 0.365000 2.730000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.160000 0.750000 3.535000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.865000 0.995000 2.240000 1.410000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.629500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.255000 0.825000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  1.665000 0.375000 2.635000 ;
      RECT 0.175000  0.085000 0.345000 0.555000 ;
      RECT 0.995000  0.655000 2.240000 0.825000 ;
      RECT 0.995000  0.825000 1.430000 1.690000 ;
      RECT 0.995000  1.690000 2.040000 1.920000 ;
      RECT 1.055000  2.220000 1.485000 2.635000 ;
      RECT 1.275000  0.085000 1.655000 0.445000 ;
      RECT 1.675000  1.920000 2.040000 2.465000 ;
      RECT 2.050000  0.255000 2.240000 0.655000 ;
      RECT 2.260000  1.670000 3.475000 1.935000 ;
      RECT 2.260000  1.935000 2.485000 2.465000 ;
      RECT 2.705000  2.125000 3.035000 2.635000 ;
      RECT 3.155000  0.085000 3.535000 0.565000 ;
      RECT 3.255000  1.935000 3.475000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_2


MACRO sky130_fd_sc_hdll__a21o_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 1.015000 2.215000 1.325000 ;
        RECT 1.985000 0.375000 2.215000 1.015000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.410000 0.995000 2.660000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.015000 1.610000 1.325000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.265000 0.355000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.525000  1.905000 0.915000 2.635000 ;
      RECT 0.545000  0.635000 1.815000 0.835000 ;
      RECT 0.545000  0.835000 0.885000 1.505000 ;
      RECT 0.545000  1.505000 1.365000 1.725000 ;
      RECT 0.665000  0.085000 1.335000 0.455000 ;
      RECT 1.095000  1.725000 1.365000 2.455000 ;
      RECT 1.515000  0.265000 1.815000 0.635000 ;
      RECT 1.595000  1.505000 2.865000 1.745000 ;
      RECT 1.595000  1.745000 1.825000 2.455000 ;
      RECT 2.005000  1.925000 2.385000 2.635000 ;
      RECT 2.575000  0.085000 2.865000 0.815000 ;
      RECT 2.605000  1.745000 2.865000 2.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_1


MACRO sky130_fd_sc_hdll__a21o_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.820000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 1.055000 1.535000 1.290000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.055000 0.695000 1.290000 ;
        RECT 0.525000 1.290000 0.695000 1.460000 ;
        RECT 0.525000 1.460000 1.875000 1.630000 ;
        RECT 1.705000 1.055000 2.045000 1.290000 ;
        RECT 1.705000 1.290000 1.875000 1.460000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 1.055000 3.195000 1.615000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.862000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.905000 0.255000 4.235000 0.695000 ;
        RECT 3.905000 0.695000 7.055000 0.865000 ;
        RECT 3.935000 1.445000 7.025000 1.615000 ;
        RECT 3.935000 1.615000 4.205000 2.465000 ;
        RECT 4.845000 0.255000 5.175000 0.695000 ;
        RECT 4.875000 1.615000 5.145000 2.465000 ;
        RECT 5.785000 0.255000 6.115000 0.695000 ;
        RECT 5.815000 1.615000 6.085000 2.465000 ;
        RECT 6.545000 0.865000 6.795000 1.445000 ;
        RECT 6.725000 0.255000 7.055000 0.695000 ;
        RECT 6.755000 1.615000 7.025000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.095000  1.460000 0.355000 1.800000 ;
      RECT 0.095000  1.800000 2.275000 1.970000 ;
      RECT 0.095000  1.970000 0.425000 2.465000 ;
      RECT 0.205000  0.085000 0.535000 0.885000 ;
      RECT 0.595000  2.140000 0.865000 2.635000 ;
      RECT 1.035000  0.275000 1.365000 0.675000 ;
      RECT 1.035000  0.675000 3.735000 0.885000 ;
      RECT 1.035000  1.970000 1.365000 2.465000 ;
      RECT 1.535000  2.140000 1.805000 2.635000 ;
      RECT 1.945000  0.085000 2.275000 0.505000 ;
      RECT 1.975000  1.970000 2.275000 2.295000 ;
      RECT 1.975000  2.295000 3.245000 2.465000 ;
      RECT 2.045000  1.460000 2.275000 1.800000 ;
      RECT 2.445000  0.255000 2.745000 0.675000 ;
      RECT 2.445000  0.885000 2.695000 1.790000 ;
      RECT 2.445000  1.790000 2.745000 2.125000 ;
      RECT 2.915000  0.085000 3.735000 0.505000 ;
      RECT 2.915000  1.785000 3.245000 2.295000 ;
      RECT 3.485000  1.495000 3.735000 2.635000 ;
      RECT 3.565000  0.885000 3.735000 1.035000 ;
      RECT 3.565000  1.035000 6.135000 1.275000 ;
      RECT 4.375000  1.785000 4.705000 2.635000 ;
      RECT 4.405000  0.085000 4.675000 0.525000 ;
      RECT 5.315000  1.785000 5.645000 2.635000 ;
      RECT 5.345000  0.085000 5.615000 0.525000 ;
      RECT 6.255000  1.785000 6.585000 2.635000 ;
      RECT 6.285000  0.085000 6.555000 0.525000 ;
      RECT 7.215000  1.445000 7.525000 2.635000 ;
      RECT 7.225000  0.085000 7.475000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_8


MACRO sky130_fd_sc_hdll__dlygate4sd1_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.605000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.830000 0.255000 3.120000 0.825000 ;
        RECT 2.860000 1.495000 3.120000 2.465000 ;
        RECT 2.950000 0.825000 3.120000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.785000 0.945000 2.005000 ;
      RECT 0.085000  2.005000 0.380000 2.465000 ;
      RECT 0.095000  0.255000 0.380000 0.715000 ;
      RECT 0.095000  0.715000 0.945000 0.885000 ;
      RECT 0.600000  0.085000 0.815000 0.545000 ;
      RECT 0.600000  2.175000 0.815000 2.635000 ;
      RECT 0.775000  0.885000 0.945000 0.995000 ;
      RECT 0.775000  0.995000 1.080000 1.325000 ;
      RECT 0.775000  1.325000 0.945000 1.785000 ;
      RECT 0.985000  0.255000 1.420000 0.545000 ;
      RECT 0.985000  2.175000 1.420000 2.465000 ;
      RECT 1.250000  0.545000 1.420000 1.075000 ;
      RECT 1.250000  1.075000 2.000000 1.275000 ;
      RECT 1.250000  1.275000 1.420000 2.175000 ;
      RECT 1.615000  0.255000 1.840000 0.735000 ;
      RECT 1.615000  0.735000 2.610000 0.905000 ;
      RECT 1.615000  1.575000 2.610000 1.745000 ;
      RECT 1.615000  1.745000 1.840000 2.430000 ;
      RECT 2.145000  0.085000 2.555000 0.565000 ;
      RECT 2.145000  1.915000 2.515000 2.635000 ;
      RECT 2.400000  0.905000 2.610000 0.995000 ;
      RECT 2.400000  0.995000 2.730000 1.325000 ;
      RECT 2.400000  1.325000 2.610000 1.575000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlygate4sd1_1


MACRO sky130_fd_sc_hdll__mux2i_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.200000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 0.995000 1.235000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.355000 0.995000 4.050000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.387500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.245000 1.075000 6.530000 1.290000 ;
        RECT 6.360000 1.290000 6.530000 1.425000 ;
        RECT 6.360000 1.425000 8.650000 1.595000 ;
        RECT 8.480000 0.995000 8.650000 1.425000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  2.339500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.315000 4.185000 0.485000 ;
        RECT 0.095000 0.485000 0.320000 2.255000 ;
        RECT 0.095000 2.255000 4.185000 2.425000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.515000  0.655000 1.850000 0.825000 ;
      RECT 0.515000  1.575000 6.130000 1.745000 ;
      RECT 1.455000  0.825000 1.850000 0.935000 ;
      RECT 2.395000  0.655000 6.035000 0.825000 ;
      RECT 2.395000  1.915000 7.915000 2.085000 ;
      RECT 4.375000  0.085000 4.705000 0.465000 ;
      RECT 4.375000  2.255000 4.705000 2.635000 ;
      RECT 4.925000  0.255000 5.095000 0.655000 ;
      RECT 5.265000  0.085000 5.645000 0.465000 ;
      RECT 5.265000  2.255000 5.645000 2.635000 ;
      RECT 5.865000  0.255000 6.035000 0.655000 ;
      RECT 6.205000  0.085000 6.580000 0.590000 ;
      RECT 6.205000  2.255000 6.585000 2.635000 ;
      RECT 6.800000  0.255000 6.975000 0.715000 ;
      RECT 6.800000  0.715000 7.915000 0.905000 ;
      RECT 6.800000  0.905000 7.100000 0.935000 ;
      RECT 6.805000  1.795000 6.975000 1.915000 ;
      RECT 6.805000  2.085000 6.975000 2.465000 ;
      RECT 7.145000  2.255000 7.525000 2.635000 ;
      RECT 7.245000  0.085000 7.495000 0.545000 ;
      RECT 7.430000  1.075000 8.310000 1.245000 ;
      RECT 7.745000  0.510000 7.915000 0.715000 ;
      RECT 7.745000  1.795000 7.915000 1.915000 ;
      RECT 7.745000  2.085000 7.915000 2.465000 ;
      RECT 8.090000  0.655000 9.045000 0.825000 ;
      RECT 8.090000  0.825000 8.310000 1.075000 ;
      RECT 8.235000  0.085000 8.565000 0.465000 ;
      RECT 8.235000  2.255000 8.565000 2.635000 ;
      RECT 8.785000  0.255000 9.045000 0.655000 ;
      RECT 8.785000  1.795000 9.045000 2.465000 ;
      RECT 8.870000  0.825000 9.045000 1.795000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.680000  0.765000 1.850000 0.935000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.800000  0.765000 6.970000 0.935000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 1.620000 0.735000 1.910000 0.780000 ;
      RECT 1.620000 0.780000 7.030000 0.920000 ;
      RECT 1.620000 0.920000 1.910000 0.965000 ;
      RECT 6.690000 0.735000 7.030000 0.780000 ;
      RECT 6.690000 0.920000 7.030000 0.965000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2i_4


MACRO sky130_fd_sc_hdll__mux2i_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.520000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.720000 1.075000 4.025000 1.275000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.710000 0.995000 5.085000 1.615000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.832500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.830000 1.325000 ;
        RECT 0.630000 0.725000 0.830000 0.995000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  1.796300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965000 0.295000 5.425000 0.465000 ;
        RECT 2.965000 2.255000 5.425000 2.425000 ;
        RECT 5.200000 1.785000 5.425000 2.255000 ;
        RECT 5.255000 0.465000 5.425000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.675000 ;
      RECT 0.085000  0.675000 0.260000 1.495000 ;
      RECT 0.085000  1.495000 1.545000 1.665000 ;
      RECT 0.085000  1.665000 0.260000 2.135000 ;
      RECT 0.085000  2.135000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.885000 0.545000 ;
      RECT 0.515000  2.255000 0.895000 2.635000 ;
      RECT 0.985000  1.835000 1.885000 2.005000 ;
      RECT 1.115000  0.575000 1.355000 0.935000 ;
      RECT 1.325000  1.155000 2.185000 1.325000 ;
      RECT 1.325000  1.325000 1.545000 1.495000 ;
      RECT 1.455000  2.255000 1.835000 2.635000 ;
      RECT 1.585000  0.085000 1.835000 0.885000 ;
      RECT 1.715000  1.495000 3.765000 1.665000 ;
      RECT 1.715000  1.665000 1.885000 1.835000 ;
      RECT 1.805000  1.075000 2.185000 1.155000 ;
      RECT 2.055000  0.295000 2.225000 0.735000 ;
      RECT 2.055000  0.735000 3.765000 0.905000 ;
      RECT 2.055000  2.135000 2.280000 2.465000 ;
      RECT 2.110000  1.835000 3.135000 1.915000 ;
      RECT 2.110000  1.915000 4.750000 2.005000 ;
      RECT 2.110000  2.005000 2.280000 2.135000 ;
      RECT 2.525000  0.085000 2.695000 0.545000 ;
      RECT 2.525000  2.175000 2.775000 2.635000 ;
      RECT 2.965000  2.005000 4.750000 2.085000 ;
      RECT 3.385000  0.655000 3.765000 0.735000 ;
      RECT 3.385000  1.665000 3.765000 1.715000 ;
      RECT 4.200000  0.655000 4.745000 0.825000 ;
      RECT 4.200000  0.825000 4.505000 0.935000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.170000  0.765000 1.340000 0.935000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.200000  0.765000 4.370000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
    LAYER met1 ;
      RECT 1.110000 0.735000 1.400000 0.780000 ;
      RECT 1.110000 0.780000 4.480000 0.920000 ;
      RECT 1.110000 0.920000 1.400000 0.965000 ;
      RECT 4.140000 0.735000 4.480000 0.780000 ;
      RECT 4.140000 0.920000 4.480000 0.965000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2i_2


MACRO sky130_fd_sc_hdll__mux2i_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.060000 0.420000 1.285000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 0.995000 1.265000 1.325000 ;
        RECT 1.065000 1.325000 1.265000 2.110000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 0.760000 3.750000 1.620000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  0.465500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.595000 0.835000 1.455000 ;
        RECT 0.605000 1.455000 0.890000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.255000 1.855000 0.425000 ;
      RECT 0.085000  0.425000 0.440000 0.465000 ;
      RECT 0.085000  0.465000 0.345000 0.885000 ;
      RECT 0.120000  1.455000 0.420000 2.295000 ;
      RECT 0.120000  2.295000 1.725000 2.465000 ;
      RECT 1.005000  0.655000 1.750000 0.715000 ;
      RECT 1.005000  0.715000 2.700000 0.825000 ;
      RECT 1.065000  0.425000 1.855000 0.465000 ;
      RECT 1.485000  1.075000 3.195000 1.310000 ;
      RECT 1.505000  1.480000 2.745000 1.650000 ;
      RECT 1.505000  1.650000 1.725000 2.295000 ;
      RECT 1.575000  0.825000 2.700000 0.885000 ;
      RECT 1.895000  1.835000 2.175000 2.635000 ;
      RECT 2.025000  0.085000 2.195000 0.525000 ;
      RECT 2.365000  1.650000 2.745000 2.465000 ;
      RECT 2.465000  0.255000 2.700000 0.715000 ;
      RECT 2.930000  0.255000 3.195000 1.075000 ;
      RECT 2.970000  1.310000 3.195000 2.465000 ;
      RECT 3.475000  1.835000 3.770000 2.635000 ;
      RECT 3.515000  0.085000 3.735000 0.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2i_1


MACRO sky130_fd_sc_hdll__o2bb2ai_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.435000 1.285000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.280000 0.825000 0.995000 ;
        RECT 0.605000 0.995000 1.100000 1.325000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 1.075000 3.245000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.150000 1.075000 2.615000 1.275000 ;
        RECT 2.445000 1.275000 2.615000 2.425000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.485500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.610000 0.430000 1.930000 0.790000 ;
        RECT 1.760000 0.790000 1.930000 1.445000 ;
        RECT 1.760000 1.445000 2.275000 1.665000 ;
        RECT 1.950000 1.665000 2.275000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.815000 ;
      RECT 0.150000  1.455000 0.400000 2.635000 ;
      RECT 0.620000  1.495000 1.440000 1.665000 ;
      RECT 0.620000  1.665000 0.870000 2.465000 ;
      RECT 1.000000  0.280000 1.440000 0.825000 ;
      RECT 1.090000  1.835000 1.780000 2.635000 ;
      RECT 1.270000  0.825000 1.440000 0.995000 ;
      RECT 1.270000  0.995000 1.580000 1.325000 ;
      RECT 1.270000  1.325000 1.440000 1.495000 ;
      RECT 2.100000  0.425000 2.350000 0.725000 ;
      RECT 2.100000  0.725000 3.240000 0.905000 ;
      RECT 2.520000  0.085000 2.690000 0.555000 ;
      RECT 2.860000  0.275000 3.240000 0.725000 ;
      RECT 2.950000  1.455000 3.200000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2ai_1


MACRO sky130_fd_sc_hdll__o2bb2ai_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.04000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 1.075000 3.905000 1.285000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 2.025000 1.285000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.845000 1.075000 10.940000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.065000 1.075000 8.675000 1.285000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.608500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.865000 0.645000 6.805000 0.905000 ;
        RECT 4.875000 1.455000 8.465000 1.625000 ;
        RECT 4.875000 1.625000 5.125000 2.465000 ;
        RECT 5.815000 1.625000 6.065000 2.465000 ;
        RECT 6.475000 0.905000 6.805000 1.455000 ;
        RECT 7.275000 1.625000 7.525000 2.125000 ;
        RECT 8.215000 1.625000 8.465000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.085000  0.645000  1.855000 0.905000 ;
      RECT  0.085000  0.905000  0.255000 1.455000 ;
      RECT  0.085000  1.455000  4.315000 1.625000 ;
      RECT  0.100000  0.255000  2.325000 0.475000 ;
      RECT  0.155000  1.795000  0.405000 2.635000 ;
      RECT  0.625000  1.625000  0.875000 2.465000 ;
      RECT  1.095000  1.795000  1.345000 2.635000 ;
      RECT  1.565000  1.625000  1.815000 2.465000 ;
      RECT  2.035000  1.795000  2.285000 2.635000 ;
      RECT  2.075000  0.475000  2.325000 0.725000 ;
      RECT  2.075000  0.725000  4.205000 0.905000 ;
      RECT  2.505000  1.625000  2.755000 2.465000 ;
      RECT  2.545000  0.085000  2.715000 0.555000 ;
      RECT  2.885000  0.255000  3.265000 0.725000 ;
      RECT  2.975000  1.795000  3.225000 2.635000 ;
      RECT  3.445000  1.625000  3.695000 2.465000 ;
      RECT  3.485000  0.085000  3.655000 0.555000 ;
      RECT  3.825000  0.255000  4.205000 0.725000 ;
      RECT  3.915000  1.795000  4.655000 2.635000 ;
      RECT  4.145000  1.075000  6.305000 1.285000 ;
      RECT  4.145000  1.285000  4.315000 1.455000 ;
      RECT  4.460000  0.255000  7.145000 0.475000 ;
      RECT  4.460000  0.475000  4.645000 0.835000 ;
      RECT  5.345000  1.795000  5.595000 2.635000 ;
      RECT  6.285000  1.795000  6.535000 2.635000 ;
      RECT  6.775000  1.795000  7.055000 2.295000 ;
      RECT  6.775000  2.295000  8.935000 2.465000 ;
      RECT  6.975000  0.475000  7.145000 0.735000 ;
      RECT  6.975000  0.735000 10.855000 0.905000 ;
      RECT  7.315000  0.085000  7.485000 0.555000 ;
      RECT  7.655000  0.255000  8.035000 0.725000 ;
      RECT  7.655000  0.725000 10.855000 0.735000 ;
      RECT  7.745000  1.795000  7.995000 2.295000 ;
      RECT  8.255000  0.085000  8.425000 0.555000 ;
      RECT  8.595000  0.255000  8.975000 0.725000 ;
      RECT  8.685000  1.455000 10.875000 1.625000 ;
      RECT  8.685000  1.625000  8.935000 2.295000 ;
      RECT  9.155000  1.795000  9.405000 2.635000 ;
      RECT  9.195000  0.085000  9.365000 0.555000 ;
      RECT  9.535000  0.255000  9.915000 0.725000 ;
      RECT  9.625000  1.625000  9.875000 2.465000 ;
      RECT 10.095000  1.795000 10.345000 2.635000 ;
      RECT 10.135000  0.085000 10.305000 0.555000 ;
      RECT 10.475000  0.255000 10.855000 0.725000 ;
      RECT 10.565000  1.625000 10.875000 2.465000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2ai_4


MACRO sky130_fd_sc_hdll__o2bb2ai_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.675000 1.445000 ;
        RECT 0.090000 1.445000 2.145000 1.615000 ;
        RECT 1.765000 1.075000 2.145000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845000 1.075000 1.500000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.650000 1.075000 4.040000 1.445000 ;
        RECT 3.650000 1.445000 5.460000 1.615000 ;
        RECT 5.130000 1.075000 5.460000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.260000 1.075000 4.900000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.788000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895000 0.645000 3.275000 1.075000 ;
        RECT 2.895000 1.075000 3.465000 1.785000 ;
        RECT 2.895000 1.785000 4.680000 1.955000 ;
        RECT 2.895000 1.955000 3.235000 2.465000 ;
        RECT 4.430000 1.955000 4.680000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.150000  1.795000 0.400000 2.635000 ;
      RECT 0.195000  0.085000 0.365000 0.895000 ;
      RECT 0.535000  0.305000 1.855000 0.475000 ;
      RECT 0.535000  0.475000 0.835000 0.895000 ;
      RECT 0.625000  1.785000 2.485000 1.965000 ;
      RECT 0.625000  1.965000 0.875000 2.465000 ;
      RECT 1.005000  0.645000 1.385000 0.725000 ;
      RECT 1.005000  0.725000 2.485000 0.905000 ;
      RECT 1.095000  2.135000 1.345000 2.635000 ;
      RECT 2.035000  0.085000 2.205000 0.555000 ;
      RECT 2.035000  2.135000 2.725000 2.635000 ;
      RECT 2.315000  0.905000 2.485000 0.995000 ;
      RECT 2.315000  0.995000 2.725000 1.325000 ;
      RECT 2.315000  1.325000 2.485000 1.785000 ;
      RECT 2.475000  0.255000 3.780000 0.475000 ;
      RECT 2.475000  0.475000 2.725000 0.555000 ;
      RECT 3.455000  2.125000 3.740000 2.635000 ;
      RECT 3.495000  0.475000 3.780000 0.735000 ;
      RECT 3.495000  0.735000 5.660000 0.905000 ;
      RECT 3.960000  2.125000 4.210000 2.295000 ;
      RECT 3.960000  2.295000 5.150000 2.465000 ;
      RECT 4.000000  0.085000 4.170000 0.555000 ;
      RECT 4.340000  0.255000 4.720000 0.725000 ;
      RECT 4.340000  0.725000 5.660000 0.735000 ;
      RECT 4.900000  1.785000 5.150000 2.295000 ;
      RECT 4.940000  0.085000 5.110000 0.555000 ;
      RECT 5.280000  0.255000 5.660000 0.725000 ;
      RECT 5.415000  1.795000 5.620000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2ai_2


MACRO sky130_fd_sc_hdll__nor2b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.520000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.075000 1.950000 1.275000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.075000 5.425000 1.320000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  1.444500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 3.735000 0.905000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 2.415000 0.255000 2.795000 0.725000 ;
        RECT 2.545000 0.905000 2.875000 1.415000 ;
        RECT 2.545000 1.415000 3.655000 1.745000 ;
        RECT 2.545000 1.745000 2.715000 2.125000 ;
        RECT 3.355000 0.255000 3.735000 0.725000 ;
        RECT 3.485000 1.745000 3.655000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.905000 ;
      RECT 0.085000  1.455000 2.325000 1.665000 ;
      RECT 0.085000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.915000 2.635000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 1.135000  1.665000 1.305000 2.465000 ;
      RECT 1.475000  1.835000 1.775000 2.635000 ;
      RECT 1.945000  1.665000 2.325000 2.295000 ;
      RECT 1.945000  2.295000 4.225000 2.465000 ;
      RECT 2.075000  0.085000 2.245000 0.555000 ;
      RECT 2.885000  1.935000 3.265000 2.295000 ;
      RECT 3.015000  0.085000 3.185000 0.555000 ;
      RECT 3.065000  1.075000 4.755000 1.245000 ;
      RECT 3.825000  1.575000 4.225000 2.295000 ;
      RECT 3.955000  0.085000 4.125000 0.905000 ;
      RECT 4.395000  0.255000 4.755000 1.075000 ;
      RECT 4.395000  1.245000 4.755000 2.465000 ;
      RECT 4.975000  0.085000 5.265000 0.905000 ;
      RECT 4.975000  1.495000 5.380000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2b_4


MACRO sky130_fd_sc_hdll__nor2b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.065000 1.285000 1.325000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.975000 0.785000 1.745000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135000 0.255000 1.515000 0.725000 ;
        RECT 1.135000 0.725000 2.215000 0.895000 ;
        RECT 1.655000 1.850000 2.215000 2.465000 ;
        RECT 2.035000 0.895000 2.215000 1.850000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.095000  0.290000 0.345000 1.915000 ;
      RECT 0.095000  1.915000 1.485000 2.085000 ;
      RECT 0.675000  0.085000 0.965000 0.625000 ;
      RECT 0.775000  2.255000 1.105000 2.635000 ;
      RECT 1.315000  1.495000 1.655000 1.665000 ;
      RECT 1.315000  1.665000 1.485000 1.915000 ;
      RECT 1.485000  1.075000 1.865000 1.325000 ;
      RECT 1.485000  1.325000 1.655000 1.495000 ;
      RECT 1.735000  0.085000 2.120000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2b_1


MACRO sky130_fd_sc_hdll__nor2b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.480000 1.065000 1.260000 1.275000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.960000 1.065000 3.535000 1.275000 ;
        RECT 3.270000 1.275000 3.535000 1.965000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.738500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.935000 0.725000 ;
        RECT 0.535000 0.725000 1.855000 0.895000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 1.565000 0.895000 1.815000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.895000 ;
      RECT 0.085000  1.445000 1.345000 1.655000 ;
      RECT 0.085000  1.655000 0.405000 2.465000 ;
      RECT 0.625000  1.825000 0.875000 2.635000 ;
      RECT 1.095000  1.655000 1.345000 2.295000 ;
      RECT 1.095000  2.295000 2.325000 2.465000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 2.035000  1.445000 2.325000 2.295000 ;
      RECT 2.075000  0.085000 2.245000 0.895000 ;
      RECT 2.075000  1.075000 2.765000 1.245000 ;
      RECT 2.595000  0.445000 2.765000 1.075000 ;
      RECT 2.595000  1.245000 2.765000 2.460000 ;
      RECT 3.185000  0.085000 3.440000 0.845000 ;
      RECT 3.185000  2.145000 3.435000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2b_2


MACRO sky130_fd_sc_hdll__muxb4to1_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  25.76000 BY  2.720000 ;
  SITE unithd ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 1.055000 1.785000 1.325000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.095000 1.055000 12.485000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.275000 1.055000 14.665000 1.325000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 23.975000 1.055000 25.365000 1.325000 ;
    END
  END D[3]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 0.995000 6.355000 1.325000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.525000 0.995000 7.120000 1.325000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.640000 0.995000 19.235000 1.325000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.405000 0.995000 20.000000 1.325000 ;
    END
  END S[3]
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  2.985000 1.755000  3.275000 1.800000 ;
        RECT  2.985000 1.800000 22.775000 1.940000 ;
        RECT  2.985000 1.940000  3.275000 1.985000 ;
        RECT  3.925000 1.755000  4.215000 1.800000 ;
        RECT  3.925000 1.940000  4.215000 1.985000 ;
        RECT  8.665000 1.755000  8.955000 1.800000 ;
        RECT  8.665000 1.940000  8.955000 1.985000 ;
        RECT  9.605000 1.755000  9.895000 1.800000 ;
        RECT  9.605000 1.940000  9.895000 1.985000 ;
        RECT 15.865000 1.755000 16.155000 1.800000 ;
        RECT 15.865000 1.940000 16.155000 1.985000 ;
        RECT 16.805000 1.755000 17.095000 1.800000 ;
        RECT 16.805000 1.940000 17.095000 1.985000 ;
        RECT 21.545000 1.755000 21.835000 1.800000 ;
        RECT 21.545000 1.940000 21.835000 1.985000 ;
        RECT 22.485000 1.755000 22.775000 1.800000 ;
        RECT 22.485000 1.940000 22.775000 1.985000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 25.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 25.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 25.760000 0.085000 ;
      RECT  0.000000  2.635000 25.760000 2.805000 ;
      RECT  0.125000  1.495000  0.395000 2.635000 ;
      RECT  0.145000  0.085000  0.395000 0.885000 ;
      RECT  0.565000  0.255000  0.895000 0.715000 ;
      RECT  0.565000  0.715000  2.695000 0.885000 ;
      RECT  0.565000  1.495000  2.795000 1.665000 ;
      RECT  0.565000  1.665000  0.895000 2.465000 ;
      RECT  1.065000  0.085000  1.335000 0.545000 ;
      RECT  1.065000  1.835000  1.335000 2.635000 ;
      RECT  1.505000  0.255000  1.835000 0.715000 ;
      RECT  1.505000  1.665000  1.835000 2.465000 ;
      RECT  2.005000  0.085000  2.255000 0.545000 ;
      RECT  2.005000  1.835000  2.275000 2.635000 ;
      RECT  2.425000  0.255000  4.455000 0.425000 ;
      RECT  2.425000  0.425000  2.695000 0.715000 ;
      RECT  2.495000  1.665000  2.795000 2.295000 ;
      RECT  2.495000  2.295000  4.705000 2.465000 ;
      RECT  2.865000  0.595000  3.195000 0.885000 ;
      RECT  2.965000  0.885000  3.195000 1.065000 ;
      RECT  2.965000  1.065000  4.235000 1.365000 ;
      RECT  2.965000  1.365000  3.295000 2.125000 ;
      RECT  3.365000  0.425000  3.535000 0.770000 ;
      RECT  3.465000  1.535000  3.735000 2.295000 ;
      RECT  3.705000  0.595000  4.035000 1.065000 ;
      RECT  3.905000  1.365000  4.235000 2.125000 ;
      RECT  4.205000  0.425000  4.455000 0.770000 ;
      RECT  4.405000  1.065000  5.590000 1.395000 ;
      RECT  4.405000  1.565000  4.705000 2.295000 ;
      RECT  4.950000  1.605000  5.225000 2.635000 ;
      RECT  4.960000  0.085000  5.250000 0.610000 ;
      RECT  5.420000  0.280000  5.670000 0.825000 ;
      RECT  5.420000  0.825000  5.590000 1.065000 ;
      RECT  5.420000  1.395000  5.590000 1.605000 ;
      RECT  5.420000  1.605000  5.750000 2.465000 ;
      RECT  5.880000  0.085000  6.170000 0.610000 ;
      RECT  5.920000  1.605000  6.220000 2.635000 ;
      RECT  6.660000  1.605000  6.960000 2.635000 ;
      RECT  6.710000  0.085000  7.000000 0.610000 ;
      RECT  7.130000  1.605000  7.460000 2.465000 ;
      RECT  7.210000  0.280000  7.460000 0.825000 ;
      RECT  7.290000  0.825000  7.460000 1.065000 ;
      RECT  7.290000  1.065000  8.475000 1.395000 ;
      RECT  7.290000  1.395000  7.460000 1.605000 ;
      RECT  7.630000  0.085000  7.920000 0.610000 ;
      RECT  7.655000  1.605000  7.930000 2.635000 ;
      RECT  8.175000  1.565000  8.475000 2.295000 ;
      RECT  8.175000  2.295000 10.385000 2.465000 ;
      RECT  8.425000  0.255000 10.455000 0.425000 ;
      RECT  8.425000  0.425000  8.675000 0.770000 ;
      RECT  8.645000  1.065000  9.915000 1.365000 ;
      RECT  8.645000  1.365000  8.975000 2.125000 ;
      RECT  8.845000  0.595000  9.175000 1.065000 ;
      RECT  9.145000  1.535000  9.415000 2.295000 ;
      RECT  9.345000  0.425000  9.515000 0.770000 ;
      RECT  9.585000  1.365000  9.915000 2.125000 ;
      RECT  9.685000  0.595000 10.015000 0.885000 ;
      RECT  9.685000  0.885000  9.915000 1.065000 ;
      RECT 10.085000  1.495000 12.315000 1.665000 ;
      RECT 10.085000  1.665000 10.385000 2.295000 ;
      RECT 10.185000  0.425000 10.455000 0.715000 ;
      RECT 10.185000  0.715000 12.315000 0.885000 ;
      RECT 10.605000  1.835000 10.875000 2.635000 ;
      RECT 10.625000  0.085000 10.875000 0.545000 ;
      RECT 11.045000  0.255000 11.375000 0.715000 ;
      RECT 11.045000  1.665000 11.375000 2.465000 ;
      RECT 11.545000  0.085000 11.815000 0.545000 ;
      RECT 11.545000  1.835000 11.815000 2.635000 ;
      RECT 11.985000  0.255000 12.315000 0.715000 ;
      RECT 11.985000  1.665000 12.315000 2.465000 ;
      RECT 12.485000  0.085000 12.735000 0.885000 ;
      RECT 12.485000  1.495000 12.755000 2.635000 ;
      RECT 13.005000  1.495000 13.275000 2.635000 ;
      RECT 13.025000  0.085000 13.275000 0.885000 ;
      RECT 13.445000  0.255000 13.775000 0.715000 ;
      RECT 13.445000  0.715000 15.575000 0.885000 ;
      RECT 13.445000  1.495000 15.675000 1.665000 ;
      RECT 13.445000  1.665000 13.775000 2.465000 ;
      RECT 13.945000  0.085000 14.215000 0.545000 ;
      RECT 13.945000  1.835000 14.215000 2.635000 ;
      RECT 14.385000  0.255000 14.715000 0.715000 ;
      RECT 14.385000  1.665000 14.715000 2.465000 ;
      RECT 14.885000  0.085000 15.135000 0.545000 ;
      RECT 14.885000  1.835000 15.155000 2.635000 ;
      RECT 15.305000  0.255000 17.335000 0.425000 ;
      RECT 15.305000  0.425000 15.575000 0.715000 ;
      RECT 15.375000  1.665000 15.675000 2.295000 ;
      RECT 15.375000  2.295000 17.585000 2.465000 ;
      RECT 15.745000  0.595000 16.075000 0.885000 ;
      RECT 15.845000  0.885000 16.075000 1.065000 ;
      RECT 15.845000  1.065000 17.115000 1.365000 ;
      RECT 15.845000  1.365000 16.175000 2.125000 ;
      RECT 16.245000  0.425000 16.415000 0.770000 ;
      RECT 16.345000  1.535000 16.615000 2.295000 ;
      RECT 16.585000  0.595000 16.915000 1.065000 ;
      RECT 16.785000  1.365000 17.115000 2.125000 ;
      RECT 17.085000  0.425000 17.335000 0.770000 ;
      RECT 17.285000  1.065000 18.470000 1.395000 ;
      RECT 17.285000  1.565000 17.585000 2.295000 ;
      RECT 17.830000  1.605000 18.105000 2.635000 ;
      RECT 17.840000  0.085000 18.130000 0.610000 ;
      RECT 18.300000  0.280000 18.550000 0.825000 ;
      RECT 18.300000  0.825000 18.470000 1.065000 ;
      RECT 18.300000  1.395000 18.470000 1.605000 ;
      RECT 18.300000  1.605000 18.630000 2.465000 ;
      RECT 18.760000  0.085000 19.050000 0.610000 ;
      RECT 18.800000  1.605000 19.100000 2.635000 ;
      RECT 19.540000  1.605000 19.840000 2.635000 ;
      RECT 19.590000  0.085000 19.880000 0.610000 ;
      RECT 20.010000  1.605000 20.340000 2.465000 ;
      RECT 20.090000  0.280000 20.340000 0.825000 ;
      RECT 20.170000  0.825000 20.340000 1.065000 ;
      RECT 20.170000  1.065000 21.355000 1.395000 ;
      RECT 20.170000  1.395000 20.340000 1.605000 ;
      RECT 20.510000  0.085000 20.800000 0.610000 ;
      RECT 20.535000  1.605000 20.810000 2.635000 ;
      RECT 21.055000  1.565000 21.355000 2.295000 ;
      RECT 21.055000  2.295000 23.265000 2.465000 ;
      RECT 21.305000  0.255000 23.335000 0.425000 ;
      RECT 21.305000  0.425000 21.555000 0.770000 ;
      RECT 21.525000  1.065000 22.795000 1.365000 ;
      RECT 21.525000  1.365000 21.855000 2.125000 ;
      RECT 21.725000  0.595000 22.055000 1.065000 ;
      RECT 22.025000  1.535000 22.295000 2.295000 ;
      RECT 22.225000  0.425000 22.395000 0.770000 ;
      RECT 22.465000  1.365000 22.795000 2.125000 ;
      RECT 22.565000  0.595000 22.895000 0.885000 ;
      RECT 22.565000  0.885000 22.795000 1.065000 ;
      RECT 22.965000  1.495000 25.195000 1.665000 ;
      RECT 22.965000  1.665000 23.265000 2.295000 ;
      RECT 23.065000  0.425000 23.335000 0.715000 ;
      RECT 23.065000  0.715000 25.195000 0.885000 ;
      RECT 23.485000  1.835000 23.755000 2.635000 ;
      RECT 23.505000  0.085000 23.755000 0.545000 ;
      RECT 23.925000  0.255000 24.255000 0.715000 ;
      RECT 23.925000  1.665000 24.255000 2.465000 ;
      RECT 24.425000  0.085000 24.695000 0.545000 ;
      RECT 24.425000  1.835000 24.695000 2.635000 ;
      RECT 24.865000  0.255000 25.195000 0.715000 ;
      RECT 24.865000  1.665000 25.195000 2.465000 ;
      RECT 25.365000  0.085000 25.615000 0.885000 ;
      RECT 25.365000  1.495000 25.635000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.045000  1.785000  3.215000 1.955000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  3.985000  1.785000  4.155000 1.955000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.725000  1.785000  8.895000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.665000  1.785000  9.835000 1.955000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 15.925000  1.785000 16.095000 1.955000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
      RECT 16.865000  1.785000 17.035000 1.955000 ;
      RECT 17.165000 -0.085000 17.335000 0.085000 ;
      RECT 17.165000  2.635000 17.335000 2.805000 ;
      RECT 17.625000 -0.085000 17.795000 0.085000 ;
      RECT 17.625000  2.635000 17.795000 2.805000 ;
      RECT 18.085000 -0.085000 18.255000 0.085000 ;
      RECT 18.085000  2.635000 18.255000 2.805000 ;
      RECT 18.545000 -0.085000 18.715000 0.085000 ;
      RECT 18.545000  2.635000 18.715000 2.805000 ;
      RECT 19.005000 -0.085000 19.175000 0.085000 ;
      RECT 19.005000  2.635000 19.175000 2.805000 ;
      RECT 19.465000 -0.085000 19.635000 0.085000 ;
      RECT 19.465000  2.635000 19.635000 2.805000 ;
      RECT 19.925000 -0.085000 20.095000 0.085000 ;
      RECT 19.925000  2.635000 20.095000 2.805000 ;
      RECT 20.385000 -0.085000 20.555000 0.085000 ;
      RECT 20.385000  2.635000 20.555000 2.805000 ;
      RECT 20.845000 -0.085000 21.015000 0.085000 ;
      RECT 20.845000  2.635000 21.015000 2.805000 ;
      RECT 21.305000 -0.085000 21.475000 0.085000 ;
      RECT 21.305000  2.635000 21.475000 2.805000 ;
      RECT 21.605000  1.785000 21.775000 1.955000 ;
      RECT 21.765000 -0.085000 21.935000 0.085000 ;
      RECT 21.765000  2.635000 21.935000 2.805000 ;
      RECT 22.225000 -0.085000 22.395000 0.085000 ;
      RECT 22.225000  2.635000 22.395000 2.805000 ;
      RECT 22.545000  1.785000 22.715000 1.955000 ;
      RECT 22.685000 -0.085000 22.855000 0.085000 ;
      RECT 22.685000  2.635000 22.855000 2.805000 ;
      RECT 23.145000 -0.085000 23.315000 0.085000 ;
      RECT 23.145000  2.635000 23.315000 2.805000 ;
      RECT 23.605000 -0.085000 23.775000 0.085000 ;
      RECT 23.605000  2.635000 23.775000 2.805000 ;
      RECT 24.065000 -0.085000 24.235000 0.085000 ;
      RECT 24.065000  2.635000 24.235000 2.805000 ;
      RECT 24.525000 -0.085000 24.695000 0.085000 ;
      RECT 24.525000  2.635000 24.695000 2.805000 ;
      RECT 24.985000 -0.085000 25.155000 0.085000 ;
      RECT 24.985000  2.635000 25.155000 2.805000 ;
      RECT 25.445000 -0.085000 25.615000 0.085000 ;
      RECT 25.445000  2.635000 25.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb4to1_4


MACRO sky130_fd_sc_hdll__muxb4to1_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.740000 BY  2.720000 ;
  SITE unithd ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.335000 1.055000 0.730000 1.325000 ;
        RECT 0.560000 0.395000 0.835000 0.625000 ;
        RECT 0.560000 0.625000 0.730000 1.055000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 0.395000 4.040000 0.625000 ;
        RECT 3.870000 0.625000 4.040000 1.055000 ;
        RECT 3.870000 1.055000 4.265000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 1.055000 4.870000 1.325000 ;
        RECT 4.700000 0.395000 4.975000 0.625000 ;
        RECT 4.700000 0.625000 4.870000 1.055000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.905000 0.395000 8.180000 0.625000 ;
        RECT 8.010000 0.625000 8.180000 1.055000 ;
        RECT 8.010000 1.055000 8.405000 1.325000 ;
    END
  END D[3]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 0.945000 2.155000 1.295000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.945000 2.795000 1.295000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.945000 0.945000 6.295000 1.295000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.585000 0.945000 6.935000 1.295000 ;
    END
  END S[3]
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.005000 1.755000 1.295000 1.800000 ;
        RECT 1.005000 1.800000 7.735000 1.940000 ;
        RECT 1.005000 1.940000 1.295000 1.985000 ;
        RECT 3.305000 1.755000 3.595000 1.800000 ;
        RECT 3.305000 1.940000 3.595000 1.985000 ;
        RECT 5.145000 1.755000 5.435000 1.800000 ;
        RECT 5.145000 1.940000 5.435000 1.985000 ;
        RECT 7.445000 1.755000 7.735000 1.800000 ;
        RECT 7.445000 1.940000 7.735000 1.985000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.095000  1.495000 0.425000 2.635000 ;
      RECT 0.130000  0.085000 0.390000 0.885000 ;
      RECT 0.900000  0.835000 1.290000 1.005000 ;
      RECT 0.900000  1.005000 1.070000 1.755000 ;
      RECT 0.900000  1.755000 1.295000 1.805000 ;
      RECT 0.900000  1.805000 1.420000 1.985000 ;
      RECT 1.045000  0.330000 1.290000 0.835000 ;
      RECT 1.090000  1.985000 1.420000 2.465000 ;
      RECT 1.240000  1.175000 1.630000 1.465000 ;
      RECT 1.240000  1.465000 1.940000 1.505000 ;
      RECT 1.460000  0.585000 1.900000 0.755000 ;
      RECT 1.460000  0.755000 1.630000 1.175000 ;
      RECT 1.460000  1.505000 1.940000 1.635000 ;
      RECT 1.610000  1.635000 1.940000 2.465000 ;
      RECT 1.650000  0.330000 1.900000 0.585000 ;
      RECT 2.135000  0.085000 2.465000 0.660000 ;
      RECT 2.165000  1.465000 2.465000 2.635000 ;
      RECT 2.660000  1.465000 3.360000 1.505000 ;
      RECT 2.660000  1.505000 3.140000 1.635000 ;
      RECT 2.660000  1.635000 2.990000 2.465000 ;
      RECT 2.700000  0.330000 2.950000 0.585000 ;
      RECT 2.700000  0.585000 3.140000 0.755000 ;
      RECT 2.970000  0.755000 3.140000 1.175000 ;
      RECT 2.970000  1.175000 3.360000 1.465000 ;
      RECT 3.180000  1.805000 3.700000 1.985000 ;
      RECT 3.180000  1.985000 3.510000 2.465000 ;
      RECT 3.305000  1.755000 3.700000 1.805000 ;
      RECT 3.310000  0.330000 3.555000 0.835000 ;
      RECT 3.310000  0.835000 3.700000 1.005000 ;
      RECT 3.530000  1.005000 3.700000 1.755000 ;
      RECT 4.175000  1.495000 4.565000 2.635000 ;
      RECT 4.210000  0.085000 4.530000 0.885000 ;
      RECT 5.040000  0.835000 5.430000 1.005000 ;
      RECT 5.040000  1.005000 5.210000 1.755000 ;
      RECT 5.040000  1.755000 5.435000 1.805000 ;
      RECT 5.040000  1.805000 5.560000 1.985000 ;
      RECT 5.185000  0.330000 5.430000 0.835000 ;
      RECT 5.230000  1.985000 5.560000 2.465000 ;
      RECT 5.380000  1.175000 5.770000 1.465000 ;
      RECT 5.380000  1.465000 6.080000 1.505000 ;
      RECT 5.600000  0.585000 6.040000 0.755000 ;
      RECT 5.600000  0.755000 5.770000 1.175000 ;
      RECT 5.600000  1.505000 6.080000 1.635000 ;
      RECT 5.750000  1.635000 6.080000 2.465000 ;
      RECT 5.790000  0.330000 6.040000 0.585000 ;
      RECT 6.275000  0.085000 6.605000 0.660000 ;
      RECT 6.275000  1.465000 6.575000 2.635000 ;
      RECT 6.800000  1.465000 7.500000 1.505000 ;
      RECT 6.800000  1.505000 7.280000 1.635000 ;
      RECT 6.800000  1.635000 7.130000 2.465000 ;
      RECT 6.840000  0.330000 7.090000 0.585000 ;
      RECT 6.840000  0.585000 7.280000 0.755000 ;
      RECT 7.110000  0.755000 7.280000 1.175000 ;
      RECT 7.110000  1.175000 7.500000 1.465000 ;
      RECT 7.320000  1.805000 7.840000 1.985000 ;
      RECT 7.320000  1.985000 7.650000 2.465000 ;
      RECT 7.445000  1.755000 7.840000 1.805000 ;
      RECT 7.450000  0.330000 7.695000 0.835000 ;
      RECT 7.450000  0.835000 7.840000 1.005000 ;
      RECT 7.670000  1.005000 7.840000 1.755000 ;
      RECT 8.315000  1.495000 8.645000 2.635000 ;
      RECT 8.350000  0.085000 8.610000 0.885000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  1.785000 1.235000 1.955000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  1.785000 3.535000 1.955000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  1.785000 5.375000 1.955000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  1.785000 7.675000 1.955000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb4to1_1


MACRO sky130_fd_sc_hdll__muxb4to1_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  12.88000 BY  2.720000 ;
  SITE unithd ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.055000 0.915000 1.325000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.525000 1.055000 6.345000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 1.055000 7.355000 1.325000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.965000 1.055000 12.785000 1.325000 ;
    END
  END D[3]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 1.025000 3.125000 1.295000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.025000 3.650000 1.295000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.230000 1.025000 9.565000 1.295000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.755000 1.025000 10.090000 1.295000 ;
    END
  END S[3]
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  1.465000 1.755000  1.755000 1.800000 ;
        RECT  1.465000 1.800000 11.415000 1.940000 ;
        RECT  1.465000 1.940000  1.755000 1.985000 ;
        RECT  4.685000 1.755000  4.975000 1.800000 ;
        RECT  4.685000 1.940000  4.975000 1.985000 ;
        RECT  7.905000 1.755000  8.195000 1.800000 ;
        RECT  7.905000 1.940000  8.195000 1.985000 ;
        RECT 11.125000 1.755000 11.415000 1.800000 ;
        RECT 11.125000 1.940000 11.415000 1.985000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.880000 0.085000 ;
      RECT  0.000000  2.635000 12.880000 2.805000 ;
      RECT  0.095000  1.495000  1.285000 1.665000 ;
      RECT  0.095000  1.665000  0.395000 2.210000 ;
      RECT  0.095000  2.210000  0.425000 2.465000 ;
      RECT  0.145000  0.255000  0.475000 0.715000 ;
      RECT  0.145000  0.715000  1.335000 0.885000 ;
      RECT  0.565000  1.835000  0.895000 2.105000 ;
      RECT  0.595000  2.105000  0.895000 2.635000 ;
      RECT  0.645000  0.085000  0.860000 0.545000 ;
      RECT  1.030000  0.255000  2.175000 0.425000 ;
      RECT  1.030000  0.425000  1.335000 0.715000 ;
      RECT  1.030000  0.885000  1.335000 0.925000 ;
      RECT  1.115000  1.665000  1.285000 2.295000 ;
      RECT  1.115000  2.295000  2.280000 2.465000 ;
      RECT  1.465000  1.755000  1.895000 2.125000 ;
      RECT  1.505000  0.595000  1.835000 0.885000 ;
      RECT  1.585000  0.885000  1.755000 1.755000 ;
      RECT  2.005000  0.425000  2.175000 0.770000 ;
      RECT  2.100000  1.205000  2.515000 1.305000 ;
      RECT  2.100000  1.305000  2.620000 1.465000 ;
      RECT  2.100000  1.465000  2.880000 1.475000 ;
      RECT  2.110000  1.645000  2.280000 2.295000 ;
      RECT  2.345000  0.585000  2.925000 0.755000 ;
      RECT  2.345000  0.755000  2.515000 1.205000 ;
      RECT  2.450000  1.475000  2.880000 1.635000 ;
      RECT  2.550000  1.635000  2.880000 2.465000 ;
      RECT  2.675000  0.330000  2.925000 0.585000 ;
      RECT  3.055000  1.465000  3.385000 2.635000 ;
      RECT  3.095000  0.085000  3.345000 0.660000 ;
      RECT  3.515000  0.330000  3.765000 0.585000 ;
      RECT  3.515000  0.585000  4.095000 0.755000 ;
      RECT  3.560000  1.465000  4.340000 1.475000 ;
      RECT  3.560000  1.475000  3.990000 1.635000 ;
      RECT  3.560000  1.635000  3.890000 2.465000 ;
      RECT  3.820000  1.305000  4.340000 1.465000 ;
      RECT  3.925000  0.755000  4.095000 1.205000 ;
      RECT  3.925000  1.205000  4.340000 1.305000 ;
      RECT  4.160000  1.645000  4.330000 2.295000 ;
      RECT  4.160000  2.295000  5.325000 2.465000 ;
      RECT  4.265000  0.255000  5.410000 0.425000 ;
      RECT  4.265000  0.425000  4.435000 0.770000 ;
      RECT  4.545000  1.755000  4.975000 2.125000 ;
      RECT  4.605000  0.595000  4.935000 0.885000 ;
      RECT  4.685000  0.885000  4.855000 1.755000 ;
      RECT  5.105000  0.425000  5.410000 0.715000 ;
      RECT  5.105000  0.715000  6.295000 0.885000 ;
      RECT  5.105000  0.885000  5.410000 0.925000 ;
      RECT  5.155000  1.495000  6.345000 1.665000 ;
      RECT  5.155000  1.665000  5.325000 2.295000 ;
      RECT  5.545000  1.835000  5.875000 2.105000 ;
      RECT  5.545000  2.105000  5.845000 2.635000 ;
      RECT  5.580000  0.085000  5.795000 0.545000 ;
      RECT  5.965000  0.255000  6.295000 0.715000 ;
      RECT  6.015000  2.210000  6.345000 2.465000 ;
      RECT  6.045000  1.665000  6.345000 2.210000 ;
      RECT  6.535000  1.495000  7.725000 1.665000 ;
      RECT  6.535000  1.665000  6.835000 2.210000 ;
      RECT  6.535000  2.210000  6.865000 2.465000 ;
      RECT  6.585000  0.255000  6.915000 0.715000 ;
      RECT  6.585000  0.715000  7.775000 0.885000 ;
      RECT  7.005000  1.835000  7.335000 2.105000 ;
      RECT  7.035000  2.105000  7.335000 2.635000 ;
      RECT  7.085000  0.085000  7.300000 0.545000 ;
      RECT  7.470000  0.255000  8.615000 0.425000 ;
      RECT  7.470000  0.425000  7.775000 0.715000 ;
      RECT  7.470000  0.885000  7.775000 0.925000 ;
      RECT  7.555000  1.665000  7.725000 2.295000 ;
      RECT  7.555000  2.295000  8.720000 2.465000 ;
      RECT  7.905000  1.755000  8.335000 2.125000 ;
      RECT  7.945000  0.595000  8.275000 0.885000 ;
      RECT  8.025000  0.885000  8.195000 1.755000 ;
      RECT  8.445000  0.425000  8.615000 0.770000 ;
      RECT  8.540000  1.205000  8.955000 1.305000 ;
      RECT  8.540000  1.305000  9.060000 1.465000 ;
      RECT  8.540000  1.465000  9.320000 1.475000 ;
      RECT  8.550000  1.645000  8.720000 2.295000 ;
      RECT  8.785000  0.585000  9.365000 0.755000 ;
      RECT  8.785000  0.755000  8.955000 1.205000 ;
      RECT  8.890000  1.475000  9.320000 1.635000 ;
      RECT  8.990000  1.635000  9.320000 2.465000 ;
      RECT  9.115000  0.330000  9.365000 0.585000 ;
      RECT  9.495000  1.465000  9.825000 2.635000 ;
      RECT  9.535000  0.085000  9.785000 0.660000 ;
      RECT  9.955000  0.330000 10.205000 0.585000 ;
      RECT  9.955000  0.585000 10.535000 0.755000 ;
      RECT 10.000000  1.465000 10.780000 1.475000 ;
      RECT 10.000000  1.475000 10.430000 1.635000 ;
      RECT 10.000000  1.635000 10.330000 2.465000 ;
      RECT 10.260000  1.305000 10.780000 1.465000 ;
      RECT 10.365000  0.755000 10.535000 1.205000 ;
      RECT 10.365000  1.205000 10.780000 1.305000 ;
      RECT 10.600000  1.645000 10.770000 2.295000 ;
      RECT 10.600000  2.295000 11.765000 2.465000 ;
      RECT 10.705000  0.255000 11.850000 0.425000 ;
      RECT 10.705000  0.425000 10.875000 0.770000 ;
      RECT 10.985000  1.755000 11.415000 2.125000 ;
      RECT 11.045000  0.595000 11.375000 0.885000 ;
      RECT 11.125000  0.885000 11.295000 1.755000 ;
      RECT 11.545000  0.425000 11.850000 0.715000 ;
      RECT 11.545000  0.715000 12.735000 0.885000 ;
      RECT 11.545000  0.885000 11.850000 0.925000 ;
      RECT 11.595000  1.495000 12.785000 1.665000 ;
      RECT 11.595000  1.665000 11.765000 2.295000 ;
      RECT 11.985000  1.835000 12.315000 2.105000 ;
      RECT 11.985000  2.105000 12.285000 2.635000 ;
      RECT 12.020000  0.085000 12.235000 0.545000 ;
      RECT 12.405000  0.255000 12.735000 0.715000 ;
      RECT 12.455000  2.210000 12.785000 2.465000 ;
      RECT 12.485000  1.665000 12.785000 2.210000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.785000  1.695000 1.955000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.785000  4.915000 1.955000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  1.785000  8.135000 1.955000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  1.785000 11.355000 1.955000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb4to1_2


MACRO sky130_fd_sc_hdll__sdfbbp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  15.64000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.155000 1.325000 4.475000 2.375000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.260000 0.255000 15.545000 0.825000 ;
        RECT 15.260000 1.605000 15.545000 2.465000 ;
        RECT 15.310000 0.825000 15.545000 1.605000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.595800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.715000 0.255000 14.115000 0.715000 ;
        RECT 13.715000 1.630000 14.095000 2.465000 ;
        RECT 13.820000 0.715000 14.115000 1.520000 ;
        RECT 13.820000 1.520000 14.095000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.515000 1.095000 13.090000 1.325000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.490000 1.025000 1.765000 1.685000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.277200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.760000 2.255000 0.765000 ;
        RECT 1.935000 0.765000 2.605000 1.015000 ;
        RECT 1.935000 1.015000 2.255000 1.695000 ;
        RECT 1.975000 0.345000 2.255000 0.760000 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  6.525000 0.735000  6.815000 0.780000 ;
        RECT  6.525000 0.780000 10.945000 0.920000 ;
        RECT  6.525000 0.920000  6.815000 0.965000 ;
        RECT 10.655000 0.735000 10.945000 0.780000 ;
        RECT 10.655000 0.920000 10.945000 0.965000 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 15.640000 0.085000 ;
        RECT  0.515000  0.085000  0.895000 0.465000 ;
        RECT  1.555000  0.085000  1.805000 0.635000 ;
        RECT  3.620000  0.085000  3.950000 0.445000 ;
        RECT  6.385000  0.085000  6.555000 0.525000 ;
        RECT  8.290000  0.085000  8.675000 0.465000 ;
        RECT 10.410000  0.085000 10.720000 0.525000 ;
        RECT 13.100000  0.085000 13.430000 0.805000 ;
        RECT 14.750000  0.085000 15.040000 0.545000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.640000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 15.640000 2.805000 ;
        RECT  0.515000 2.135000  0.895000 2.635000 ;
        RECT  1.555000 1.885000  1.885000 2.635000 ;
        RECT  3.510000 2.215000  3.890000 2.635000 ;
        RECT  6.205000 2.205000  6.585000 2.635000 ;
        RECT  7.825000 1.915000  8.155000 2.635000 ;
        RECT 10.520000 2.255000 10.900000 2.635000 ;
        RECT 11.940000 2.255000 13.430000 2.635000 ;
        RECT 14.745000 1.765000 15.040000 2.635000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 15.640000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.170000 0.345000  0.345000 0.635000 ;
      RECT  0.170000 0.635000  0.885000 0.805000 ;
      RECT  0.170000 1.795000  0.885000 1.965000 ;
      RECT  0.170000 1.965000  0.345000 2.465000 ;
      RECT  0.655000 0.805000  0.885000 1.795000 ;
      RECT  1.115000 0.345000  1.320000 2.465000 ;
      RECT  2.385000 1.875000  2.765000 2.385000 ;
      RECT  2.550000 0.265000  2.955000 0.595000 ;
      RECT  2.550000 1.185000  3.275000 1.365000 ;
      RECT  2.550000 1.365000  2.765000 1.875000 ;
      RECT  2.785000 0.595000  2.955000 1.075000 ;
      RECT  2.785000 1.075000  3.275000 1.185000 ;
      RECT  2.945000 1.575000  3.895000 1.745000 ;
      RECT  2.945000 1.745000  3.265000 1.905000 ;
      RECT  3.095000 1.905000  3.265000 2.465000 ;
      RECT  3.125000 0.305000  3.325000 0.625000 ;
      RECT  3.125000 0.625000  3.895000 0.765000 ;
      RECT  3.125000 0.765000  4.070000 0.795000 ;
      RECT  3.725000 0.795000  4.070000 1.095000 ;
      RECT  3.725000 1.095000  3.895000 1.575000 ;
      RECT  4.645000 0.305000  4.815000 2.465000 ;
      RECT  4.985000 0.705000  5.245000 1.575000 ;
      RECT  4.985000 1.575000  5.575000 1.955000 ;
      RECT  5.035000 2.250000  5.915000 2.420000 ;
      RECT  5.100000 0.265000  6.215000 0.465000 ;
      RECT  5.425000 0.645000  5.825000 1.015000 ;
      RECT  5.745000 1.195000  6.215000 1.235000 ;
      RECT  5.745000 1.235000  7.195000 1.405000 ;
      RECT  5.745000 1.405000  5.915000 2.250000 ;
      RECT  5.995000 0.465000  6.215000 1.195000 ;
      RECT  6.085000 1.575000  6.385000 1.785000 ;
      RECT  6.085000 1.785000  7.585000 2.035000 ;
      RECT  6.385000 0.735000  6.795000 1.065000 ;
      RECT  6.775000 0.255000  8.045000 0.425000 ;
      RECT  6.775000 0.425000  7.105000 0.465000 ;
      RECT  6.935000 2.035000  7.105000 2.375000 ;
      RECT  6.945000 1.405000  7.195000 1.485000 ;
      RECT  6.975000 1.155000  7.195000 1.235000 ;
      RECT  7.275000 0.595000  7.655000 0.765000 ;
      RECT  7.415000 0.765000  7.655000 0.895000 ;
      RECT  7.415000 0.895000  8.875000 1.065000 ;
      RECT  7.415000 1.065000  7.585000 1.785000 ;
      RECT  7.805000 1.235000  8.135000 1.415000 ;
      RECT  7.805000 1.415000  8.910000 1.655000 ;
      RECT  7.850000 0.425000  8.045000 0.715000 ;
      RECT  8.445000 1.065000  8.875000 1.235000 ;
      RECT  9.110000 1.575000  9.345000 1.985000 ;
      RECT  9.170000 0.705000  9.510000 1.125000 ;
      RECT  9.170000 1.125000  9.890000 1.305000 ;
      RECT  9.300000 2.250000 10.230000 2.420000 ;
      RECT  9.415000 0.265000 10.230000 0.465000 ;
      RECT  9.635000 1.305000  9.890000 1.905000 ;
      RECT 10.060000 0.465000 10.230000 1.235000 ;
      RECT 10.060000 1.235000 11.510000 1.405000 ;
      RECT 10.060000 1.405000 10.230000 2.250000 ;
      RECT 10.400000 1.575000 10.700000 1.915000 ;
      RECT 10.400000 1.915000 13.430000 2.085000 ;
      RECT 10.655000 0.735000 11.080000 1.065000 ;
      RECT 10.980000 0.255000 12.300000 0.425000 ;
      RECT 10.980000 0.425000 11.380000 0.465000 ;
      RECT 11.190000 2.085000 11.360000 2.375000 ;
      RECT 11.290000 1.075000 11.510000 1.235000 ;
      RECT 11.535000 0.645000 11.915000 0.815000 ;
      RECT 11.730000 0.815000 11.915000 1.915000 ;
      RECT 12.125000 0.425000 12.300000 0.585000 ;
      RECT 12.130000 0.755000 12.815000 0.925000 ;
      RECT 12.130000 0.925000 12.345000 1.575000 ;
      RECT 12.130000 1.575000 12.905000 1.745000 ;
      RECT 12.615000 0.265000 12.815000 0.755000 ;
      RECT 13.260000 0.995000 13.525000 1.325000 ;
      RECT 13.260000 1.325000 13.430000 1.915000 ;
      RECT 14.265000 1.725000 14.520000 2.415000 ;
      RECT 14.315000 0.255000 14.520000 0.995000 ;
      RECT 14.315000 0.995000 15.090000 1.325000 ;
      RECT 14.315000 1.325000 14.520000 1.725000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.655000  1.785000  0.825000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.150000  0.765000  1.320000 0.935000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.105000  1.105000  3.275000 1.275000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.645000  1.105000  4.815000 1.275000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.145000  1.785000  5.315000 1.955000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.655000  0.765000  5.825000 0.935000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  0.765000  6.755000 0.935000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.715000  1.445000  8.885000 1.615000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.175000  1.105000  9.345000 1.275000 ;
      RECT  9.175000  1.785000  9.345000 1.955000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.715000  0.765000 10.885000 0.935000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.165000  1.445000 12.335000 1.615000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
    LAYER met1 ;
      RECT  0.595000 1.755000  0.885000 1.800000 ;
      RECT  0.595000 1.800000  9.405000 1.940000 ;
      RECT  0.595000 1.940000  0.885000 1.985000 ;
      RECT  1.090000 0.735000  1.380000 0.780000 ;
      RECT  1.090000 0.780000  5.885000 0.920000 ;
      RECT  1.090000 0.920000  1.380000 0.965000 ;
      RECT  3.045000 1.075000  3.335000 1.120000 ;
      RECT  3.045000 1.120000  4.875000 1.260000 ;
      RECT  3.045000 1.260000  3.335000 1.305000 ;
      RECT  4.585000 1.075000  4.875000 1.120000 ;
      RECT  4.585000 1.260000  4.875000 1.305000 ;
      RECT  5.085000 1.755000  5.375000 1.800000 ;
      RECT  5.085000 1.940000  5.375000 1.985000 ;
      RECT  5.595000 0.735000  5.885000 0.780000 ;
      RECT  5.595000 0.920000  5.885000 0.965000 ;
      RECT  5.670000 0.965000  5.885000 1.120000 ;
      RECT  5.670000 1.120000  9.405000 1.260000 ;
      RECT  8.655000 1.415000  8.945000 1.460000 ;
      RECT  8.655000 1.460000 12.395000 1.600000 ;
      RECT  8.655000 1.600000  8.945000 1.645000 ;
      RECT  9.115000 1.075000  9.405000 1.120000 ;
      RECT  9.115000 1.260000  9.405000 1.305000 ;
      RECT  9.115000 1.755000  9.405000 1.800000 ;
      RECT  9.115000 1.940000  9.405000 1.985000 ;
      RECT 12.105000 1.415000 12.395000 1.460000 ;
      RECT 12.105000 1.600000 12.395000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfbbp_1


MACRO sky130_fd_sc_hdll__nand2b_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 0.995000 0.850000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 1.075000 3.095000 1.275000 ;
        RECT 2.905000 1.275000 3.095000 1.655000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.825500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135000 1.835000 2.615000 2.005000 ;
        RECT 1.135000 2.005000 1.465000 2.465000 ;
        RECT 1.455000 0.635000 1.785000 1.835000 ;
        RECT 2.285000 2.005000 2.615000 2.465000 ;
        RECT 2.340000 1.495000 2.615000 1.835000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.110000  0.510000 0.345000 0.840000 ;
      RECT 0.110000  0.840000 0.280000 1.495000 ;
      RECT 0.110000  1.495000 1.190000 1.665000 ;
      RECT 0.110000  1.665000 0.410000 1.860000 ;
      RECT 0.595000  0.085000 0.765000 0.775000 ;
      RECT 0.630000  1.835000 0.885000 2.635000 ;
      RECT 1.020000  0.995000 1.190000 1.495000 ;
      RECT 1.035000  0.255000 2.205000 0.465000 ;
      RECT 1.725000  2.175000 2.100000 2.635000 ;
      RECT 1.955000  0.465000 2.205000 0.695000 ;
      RECT 1.955000  0.695000 3.095000 0.905000 ;
      RECT 2.425000  0.085000 2.595000 0.525000 ;
      RECT 2.765000  0.255000 3.095000 0.695000 ;
      RECT 2.845000  1.835000 3.015000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2b_2


MACRO sky130_fd_sc_hdll__nand2b_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.420000 1.315000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 1.075000 1.185000 1.315000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.491500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 1.835000 2.190000 2.005000 ;
        RECT 1.050000 2.005000 1.430000 2.465000 ;
        RECT 1.360000 0.255000 2.190000 0.545000 ;
        RECT 1.820000 0.545000 2.190000 1.835000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.090000  0.525000 0.360000 0.735000 ;
      RECT 0.090000  0.735000 1.620000 0.905000 ;
      RECT 0.090000  1.495000 1.620000 1.665000 ;
      RECT 0.090000  1.665000 0.370000 1.825000 ;
      RECT 0.630000  0.085000 0.960000 0.545000 ;
      RECT 0.630000  1.835000 0.880000 2.635000 ;
      RECT 1.450000  0.905000 1.620000 1.495000 ;
      RECT 1.650000  2.175000 1.865000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2b_1


MACRO sky130_fd_sc_hdll__nand2b_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.520000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.075000 5.390000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.576000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 0.635000 2.840000 0.905000 ;
        RECT 1.505000 1.445000 4.720000 1.665000 ;
        RECT 1.505000 1.665000 1.885000 2.465000 ;
        RECT 2.445000 1.665000 2.840000 2.465000 ;
        RECT 2.575000 0.905000 2.840000 1.445000 ;
        RECT 3.400000 1.665000 3.780000 2.465000 ;
        RECT 4.340000 1.665000 4.720000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.715000 ;
      RECT 0.090000  0.715000 0.830000 0.905000 ;
      RECT 0.090000  1.445000 0.830000 1.665000 ;
      RECT 0.090000  1.665000 0.425000 2.465000 ;
      RECT 0.645000  0.085000 0.840000 0.545000 ;
      RECT 0.645000  1.835000 1.335000 2.635000 ;
      RECT 0.660000  0.905000 0.830000 1.075000 ;
      RECT 0.660000  1.075000 2.355000 1.275000 ;
      RECT 0.660000  1.275000 0.830000 1.445000 ;
      RECT 1.020000  1.445000 1.335000 1.835000 ;
      RECT 1.085000  0.255000 3.310000 0.465000 ;
      RECT 1.085000  0.465000 1.335000 0.905000 ;
      RECT 2.105000  1.835000 2.275000 2.635000 ;
      RECT 3.060000  0.465000 3.310000 0.715000 ;
      RECT 3.060000  0.715000 5.300000 0.905000 ;
      RECT 3.060000  1.835000 3.230000 2.635000 ;
      RECT 3.530000  0.085000 3.700000 0.545000 ;
      RECT 3.870000  0.255000 4.250000 0.715000 ;
      RECT 4.000000  1.835000 4.170000 2.635000 ;
      RECT 4.470000  0.085000 4.710000 0.545000 ;
      RECT 4.970000  0.255000 5.300000 0.715000 ;
      RECT 4.970000  1.495000 5.300000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2b_4


MACRO sky130_fd_sc_hdll__nand2_6
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 1.055000 5.155000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 1.055000 2.765000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.495000 5.595000 1.665000 ;
        RECT 0.565000 1.665000 0.895000 2.465000 ;
        RECT 1.505000 1.665000 1.835000 2.465000 ;
        RECT 2.445000 1.665000 2.775000 2.465000 ;
        RECT 3.335000 0.635000 5.595000 0.885000 ;
        RECT 3.335000 0.885000 3.635000 1.495000 ;
        RECT 3.385000 1.665000 3.715000 2.465000 ;
        RECT 4.325000 1.665000 4.655000 2.465000 ;
        RECT 5.265000 1.665000 5.595000 2.465000 ;
        RECT 5.325000 0.885000 5.595000 1.055000 ;
        RECT 5.325000 1.055000 5.915000 1.325000 ;
        RECT 5.325000 1.325000 5.595000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.715000 ;
      RECT 0.090000  0.715000 3.165000 0.885000 ;
      RECT 0.125000  1.495000 0.395000 2.635000 ;
      RECT 0.595000  0.085000 0.865000 0.545000 ;
      RECT 1.035000  0.255000 1.365000 0.715000 ;
      RECT 1.065000  1.835000 1.335000 2.635000 ;
      RECT 1.535000  0.085000 1.805000 0.545000 ;
      RECT 1.975000  0.255000 2.305000 0.715000 ;
      RECT 2.005000  1.835000 2.275000 2.635000 ;
      RECT 2.475000  0.085000 2.745000 0.545000 ;
      RECT 2.915000  0.255000 6.065000 0.465000 ;
      RECT 2.915000  0.465000 3.165000 0.715000 ;
      RECT 2.945000  1.835000 3.215000 2.635000 ;
      RECT 3.885000  1.835000 4.155000 2.635000 ;
      RECT 4.825000  1.835000 5.095000 2.635000 ;
      RECT 5.765000  0.465000 6.065000 0.885000 ;
      RECT 5.765000  1.495000 6.035000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_6


MACRO sky130_fd_sc_hdll__nand2_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.280000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.740000 1.075000 7.005000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.510000 1.075000 3.715000 1.295000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  3.184500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.465000 7.475000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.465000 ;
        RECT 1.455000 1.665000 1.835000 2.465000 ;
        RECT 2.395000 1.665000 2.775000 2.465000 ;
        RECT 3.335000 1.665000 3.715000 2.465000 ;
        RECT 4.040000 1.075000 4.570000 1.465000 ;
        RECT 4.275000 0.655000 7.475000 0.905000 ;
        RECT 4.275000 0.905000 4.570000 1.075000 ;
        RECT 4.275000 1.665000 4.655000 2.465000 ;
        RECT 5.215000 1.665000 5.595000 2.465000 ;
        RECT 6.155000 1.665000 6.535000 2.465000 ;
        RECT 7.095000 1.665000 7.475000 2.465000 ;
        RECT 7.225000 0.905000 7.475000 1.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 4.105000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.645000  0.085000 0.815000 0.565000 ;
      RECT 0.985000  0.255000 1.365000 0.735000 ;
      RECT 1.115000  1.835000 1.285000 2.635000 ;
      RECT 1.585000  0.085000 1.755000 0.565000 ;
      RECT 1.925000  0.255000 2.305000 0.735000 ;
      RECT 2.055000  1.835000 2.225000 2.635000 ;
      RECT 2.525000  0.085000 2.695000 0.565000 ;
      RECT 2.865000  0.255000 3.245000 0.735000 ;
      RECT 2.995000  1.835000 3.165000 2.635000 ;
      RECT 3.465000  0.085000 3.635000 0.565000 ;
      RECT 3.805000  0.255000 8.070000 0.485000 ;
      RECT 3.805000  0.485000 4.105000 0.735000 ;
      RECT 3.935000  1.835000 4.105000 2.635000 ;
      RECT 4.875000  1.835000 5.045000 2.635000 ;
      RECT 5.815000  1.835000 5.985000 2.635000 ;
      RECT 6.755000  1.835000 6.925000 2.635000 ;
      RECT 7.695000  0.485000 8.070000 0.905000 ;
      RECT 7.715000  1.495000 8.070000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_8


MACRO sky130_fd_sc_hdll__nand2_12
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.96000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  3.330000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.625000 1.055000 10.695000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  3.330000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.335000 1.055000 5.765000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  4.858000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.565000 1.495000 11.235000 1.665000 ;
        RECT  0.565000 1.665000  0.895000 2.465000 ;
        RECT  1.505000 1.665000  1.835000 2.465000 ;
        RECT  2.445000 1.665000  2.775000 2.465000 ;
        RECT  3.385000 1.665000  3.715000 2.465000 ;
        RECT  4.325000 1.665000  4.655000 2.465000 ;
        RECT  5.265000 1.665000  5.595000 2.465000 ;
        RECT  6.045000 1.055000  6.455000 1.495000 ;
        RECT  6.155000 0.635000 11.235000 0.885000 ;
        RECT  6.155000 0.885000  6.455000 1.055000 ;
        RECT  6.205000 1.665000  6.535000 2.465000 ;
        RECT  7.145000 1.665000  7.475000 2.465000 ;
        RECT  8.085000 1.665000  8.415000 2.465000 ;
        RECT  9.025000 1.665000  9.355000 2.465000 ;
        RECT  9.965000 1.665000 10.295000 2.465000 ;
        RECT 10.905000 1.665000 11.235000 2.465000 ;
        RECT 10.965000 0.885000 11.235000 1.055000 ;
        RECT 10.965000 1.055000 11.435000 1.325000 ;
        RECT 10.965000 1.325000 11.235000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.090000  0.255000  0.425000 0.715000 ;
      RECT  0.090000  0.715000  5.985000 0.885000 ;
      RECT  0.125000  1.495000  0.395000 2.635000 ;
      RECT  0.595000  0.085000  0.865000 0.545000 ;
      RECT  1.035000  0.255000  1.365000 0.715000 ;
      RECT  1.065000  1.835000  1.335000 2.635000 ;
      RECT  1.535000  0.085000  1.805000 0.545000 ;
      RECT  1.975000  0.255000  2.305000 0.715000 ;
      RECT  2.005000  1.835000  2.275000 2.635000 ;
      RECT  2.475000  0.085000  2.745000 0.545000 ;
      RECT  2.915000  0.255000  3.245000 0.715000 ;
      RECT  2.945000  1.835000  3.215000 2.635000 ;
      RECT  3.415000  0.085000  3.685000 0.545000 ;
      RECT  3.855000  0.255000  4.185000 0.715000 ;
      RECT  3.885000  1.835000  4.155000 2.635000 ;
      RECT  4.355000  0.085000  4.625000 0.545000 ;
      RECT  4.795000  0.255000  5.125000 0.715000 ;
      RECT  4.825000  1.835000  5.095000 2.635000 ;
      RECT  5.295000  0.085000  5.565000 0.545000 ;
      RECT  5.735000  0.255000 11.705000 0.465000 ;
      RECT  5.735000  0.465000  5.985000 0.715000 ;
      RECT  5.765000  1.835000  6.035000 2.635000 ;
      RECT  6.705000  1.835000  6.975000 2.635000 ;
      RECT  7.645000  1.835000  7.915000 2.635000 ;
      RECT  8.585000  1.835000  8.855000 2.635000 ;
      RECT  9.525000  1.835000  9.795000 2.635000 ;
      RECT 10.465000  1.835000 10.735000 2.635000 ;
      RECT 11.405000  1.495000 11.675000 2.635000 ;
      RECT 11.455000  0.465000 11.705000 0.885000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_12


MACRO sky130_fd_sc_hdll__nand2_16
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  15.64000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  4.440000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.505000 1.055000 14.275000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  4.440000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 1.055000 7.525000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  6.499000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.565000 1.495000 14.995000 1.665000 ;
        RECT  0.565000 1.665000  0.895000 2.465000 ;
        RECT  1.505000 1.665000  1.835000 2.465000 ;
        RECT  2.445000 1.665000  2.775000 2.465000 ;
        RECT  3.385000 1.665000  3.715000 2.465000 ;
        RECT  4.325000 1.665000  4.655000 2.465000 ;
        RECT  5.265000 1.665000  5.595000 2.465000 ;
        RECT  6.205000 1.665000  6.535000 2.465000 ;
        RECT  7.145000 1.665000  7.475000 2.465000 ;
        RECT  7.925000 1.055000  8.335000 1.495000 ;
        RECT  8.035000 0.635000 14.995000 0.885000 ;
        RECT  8.035000 0.885000  8.335000 1.055000 ;
        RECT  8.085000 1.665000  8.415000 2.465000 ;
        RECT  9.025000 1.665000  9.355000 2.465000 ;
        RECT  9.965000 1.665000 10.295000 2.465000 ;
        RECT 10.905000 1.665000 11.235000 2.465000 ;
        RECT 11.845000 1.665000 12.175000 2.465000 ;
        RECT 12.785000 1.665000 13.115000 2.465000 ;
        RECT 13.725000 1.665000 14.055000 2.465000 ;
        RECT 14.665000 1.665000 14.995000 2.465000 ;
        RECT 14.725000 0.885000 14.995000 1.055000 ;
        RECT 14.725000 1.055000 15.115000 1.325000 ;
        RECT 14.725000 1.325000 14.995000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.640000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 15.640000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.640000 0.085000 ;
      RECT  0.000000  2.635000 15.640000 2.805000 ;
      RECT  0.095000  0.255000  0.425000 0.715000 ;
      RECT  0.095000  0.715000  7.865000 0.885000 ;
      RECT  0.125000  1.495000  0.395000 2.635000 ;
      RECT  0.595000  0.085000  0.865000 0.545000 ;
      RECT  1.035000  0.255000  1.365000 0.715000 ;
      RECT  1.065000  1.835000  1.335000 2.635000 ;
      RECT  1.535000  0.085000  1.805000 0.545000 ;
      RECT  1.975000  0.255000  2.305000 0.715000 ;
      RECT  2.005000  1.835000  2.275000 2.635000 ;
      RECT  2.475000  0.085000  2.745000 0.545000 ;
      RECT  2.915000  0.255000  3.245000 0.715000 ;
      RECT  2.945000  1.835000  3.215000 2.635000 ;
      RECT  3.415000  0.085000  3.685000 0.545000 ;
      RECT  3.855000  0.255000  4.185000 0.715000 ;
      RECT  3.885000  1.835000  4.155000 2.635000 ;
      RECT  4.355000  0.085000  4.625000 0.545000 ;
      RECT  4.795000  0.255000  5.125000 0.715000 ;
      RECT  4.825000  1.835000  5.095000 2.635000 ;
      RECT  5.295000  0.085000  5.565000 0.545000 ;
      RECT  5.735000  0.255000  6.065000 0.715000 ;
      RECT  5.765000  1.835000  6.035000 2.635000 ;
      RECT  6.235000  0.085000  6.505000 0.545000 ;
      RECT  6.675000  0.255000  7.005000 0.715000 ;
      RECT  6.705000  1.835000  6.975000 2.635000 ;
      RECT  7.175000  0.085000  7.445000 0.545000 ;
      RECT  7.615000  0.255000 15.465000 0.465000 ;
      RECT  7.615000  0.465000  7.865000 0.715000 ;
      RECT  7.645000  1.835000  7.915000 2.635000 ;
      RECT  8.585000  1.835000  8.855000 2.635000 ;
      RECT  9.525000  1.835000  9.795000 2.635000 ;
      RECT 10.465000  1.835000 10.735000 2.635000 ;
      RECT 11.405000  1.835000 11.675000 2.635000 ;
      RECT 12.345000  1.835000 12.615000 2.635000 ;
      RECT 13.285000  1.835000 13.555000 2.635000 ;
      RECT 14.225000  1.835000 14.495000 2.635000 ;
      RECT 15.165000  1.495000 15.435000 2.635000 ;
      RECT 15.215000  0.465000 15.465000 0.885000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_16


MACRO sky130_fd_sc_hdll__nand2_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  1.840000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.990000 1.075000 1.375000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.055000 0.430000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.491500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 1.485000 0.915000 2.465000 ;
        RECT 0.650000 0.255000 1.395000 0.885000 ;
        RECT 0.650000 0.885000 0.820000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.085000 0.395000 0.885000 ;
      RECT 0.085000  1.495000 0.365000 2.635000 ;
      RECT 1.135000  1.495000 1.395000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_1


MACRO sky130_fd_sc_hdll__nand2_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 1.075000 4.115000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.880000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.608500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.495000 3.715000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.465000 ;
        RECT 1.455000 1.665000 1.835000 2.465000 ;
        RECT 2.395000 0.635000 3.715000 0.805000 ;
        RECT 2.395000 0.805000 2.695000 1.495000 ;
        RECT 2.395000 1.665000 2.775000 2.465000 ;
        RECT 3.335000 1.665000 3.715000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.715000 ;
      RECT 0.090000  0.715000 2.225000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.645000  0.085000 0.815000 0.545000 ;
      RECT 0.985000  0.255000 1.365000 0.715000 ;
      RECT 1.115000  1.835000 1.285000 2.635000 ;
      RECT 1.585000  0.085000 1.755000 0.545000 ;
      RECT 1.925000  0.255000 4.185000 0.465000 ;
      RECT 1.925000  0.465000 2.225000 0.715000 ;
      RECT 2.055000  1.835000 2.225000 2.635000 ;
      RECT 2.995000  1.835000 3.165000 2.635000 ;
      RECT 3.935000  0.465000 4.185000 0.885000 ;
      RECT 3.935000  1.835000 4.185000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_4


MACRO sky130_fd_sc_hdll__nand2_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.780000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.895000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.820500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.495000 2.230000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.465000 ;
        RECT 1.455000 0.655000 2.230000 0.905000 ;
        RECT 1.455000 1.665000 1.835000 2.465000 ;
        RECT 1.950000 0.905000 2.230000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.255000 0.425000 0.715000 ;
      RECT 0.085000  0.715000 1.285000 0.885000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.645000  0.085000 0.815000 0.545000 ;
      RECT 0.985000  0.255000 2.305000 0.485000 ;
      RECT 0.985000  0.485000 1.285000 0.715000 ;
      RECT 1.115000  1.835000 1.285000 2.635000 ;
      RECT 2.055000  1.835000 2.310000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand2_2


MACRO sky130_fd_sc_hdll__xor2_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.04000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 3.100000 1.275000 ;
        RECT 2.880000 1.275000 3.100000 1.445000 ;
        RECT 2.880000 1.445000 6.815000 1.615000 ;
        RECT 6.595000 1.075000 8.120000 1.275000 ;
        RECT 6.595000 1.275000 6.815000 1.445000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.270000 1.075000 5.500000 1.105000 ;
        RECT 3.270000 1.105000 6.340000 1.275000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.318500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  8.650000 0.725000  9.480000 0.735000 ;
        RECT  8.650000 0.735000 10.955000 0.905000 ;
        RECT  8.680000 1.445000 10.955000 1.625000 ;
        RECT  8.680000 1.625000  9.910000 1.665000 ;
        RECT  8.680000 1.665000  8.970000 2.125000 ;
        RECT  9.100000 0.255000  9.480000 0.725000 ;
        RECT  9.660000 1.665000  9.910000 2.125000 ;
        RECT 10.040000 0.255000 10.420000 0.735000 ;
        RECT 10.550000 1.625000 10.955000 2.465000 ;
        RECT 10.635000 0.905000 10.955000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.085000  0.085000  0.360000 0.565000 ;
      RECT  0.085000  0.735000  3.730000 0.905000 ;
      RECT  0.085000  0.905000  0.255000 1.445000 ;
      RECT  0.085000  1.445000  2.670000 1.615000 ;
      RECT  0.085000  1.785000  2.280000 2.005000 ;
      RECT  0.085000  2.005000  0.400000 2.465000 ;
      RECT  0.530000  0.255000  0.910000 0.725000 ;
      RECT  0.530000  0.725000  3.730000 0.735000 ;
      RECT  0.620000  2.175000  0.870000 2.635000 ;
      RECT  1.090000  2.005000  1.340000 2.465000 ;
      RECT  1.130000  0.085000  1.300000 0.555000 ;
      RECT  1.470000  0.255000  1.850000 0.725000 ;
      RECT  1.560000  2.175000  1.810000 2.635000 ;
      RECT  2.030000  2.005000  2.280000 2.295000 ;
      RECT  2.030000  2.295000  4.160000 2.465000 ;
      RECT  2.070000  0.085000  2.240000 0.555000 ;
      RECT  2.410000  0.255000  2.790000 0.725000 ;
      RECT  2.500000  1.615000  2.670000 1.785000 ;
      RECT  2.500000  1.785000  3.690000 1.955000 ;
      RECT  2.500000  1.955000  2.750000 2.125000 ;
      RECT  2.970000  2.125000  3.220000 2.295000 ;
      RECT  3.010000  0.085000  3.180000 0.555000 ;
      RECT  3.350000  0.255000  3.730000 0.725000 ;
      RECT  3.440000  1.955000  3.690000 2.125000 ;
      RECT  3.910000  1.795000  4.160000 2.295000 ;
      RECT  3.950000  0.085000  4.220000 0.895000 ;
      RECT  4.390000  0.255000  6.600000 0.475000 ;
      RECT  4.430000  1.785000  8.440000 2.005000 ;
      RECT  4.430000  2.005000  4.680000 2.465000 ;
      RECT  4.565000  0.645000  6.130000 0.905000 ;
      RECT  4.900000  2.175000  5.150000 2.635000 ;
      RECT  5.370000  2.005000  5.620000 2.465000 ;
      RECT  5.650000  0.905000  6.130000 0.935000 ;
      RECT  5.840000  2.175000  6.090000 2.635000 ;
      RECT  6.310000  2.005000  6.560000 2.465000 ;
      RECT  6.350000  0.475000  6.600000 0.725000 ;
      RECT  6.350000  0.725000  8.480000 0.905000 ;
      RECT  6.780000  2.175000  7.030000 2.635000 ;
      RECT  6.820000  0.085000  6.990000 0.555000 ;
      RECT  7.160000  0.255000  7.540000 0.725000 ;
      RECT  7.250000  1.455000  7.500000 1.785000 ;
      RECT  7.250000  2.005000  7.500000 2.465000 ;
      RECT  7.720000  2.175000  7.970000 2.635000 ;
      RECT  7.760000  0.085000  7.930000 0.555000 ;
      RECT  8.010000  1.445000  8.510000 1.615000 ;
      RECT  8.100000  0.255000  8.480000 0.725000 ;
      RECT  8.190000  2.005000  8.440000 2.295000 ;
      RECT  8.190000  2.295000 10.380000 2.465000 ;
      RECT  8.340000  1.075000 10.130000 1.275000 ;
      RECT  8.340000  1.275000  8.510000 1.445000 ;
      RECT  8.760000  0.085000  8.930000 0.555000 ;
      RECT  9.190000  1.835000  9.440000 2.295000 ;
      RECT  9.700000  0.085000  9.870000 0.555000 ;
      RECT 10.130000  1.795000 10.380000 2.295000 ;
      RECT 10.640000  0.085000 10.810000 0.555000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.185000  1.445000  2.355000 1.615000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.705000  0.725000  5.875000 0.895000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.305000  1.445000  8.475000 1.615000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.765000  0.725000  8.935000 0.895000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 2.125000 1.415000 2.415000 1.460000 ;
      RECT 2.125000 1.460000 8.535000 1.600000 ;
      RECT 2.125000 1.600000 2.415000 1.645000 ;
      RECT 5.645000 0.695000 5.935000 0.780000 ;
      RECT 5.645000 0.780000 8.995000 0.925000 ;
      RECT 8.245000 1.415000 8.535000 1.460000 ;
      RECT 8.245000 1.600000 8.535000 1.645000 ;
      RECT 8.705000 0.695000 8.995000 0.780000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor2_4


MACRO sky130_fd_sc_hdll__xor2_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.680000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.075000 1.500000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.445000 ;
        RECT 0.425000 1.445000 1.890000 1.615000 ;
        RECT 1.720000 1.075000 2.155000 1.245000 ;
        RECT 1.720000 1.245000 1.890000 1.445000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.880000 0.315000 3.085000 0.485000 ;
        RECT 2.915000 0.485000 3.085000 1.365000 ;
        RECT 2.915000 1.365000 3.545000 1.535000 ;
        RECT 3.225000 1.535000 3.545000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.655000 2.745000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.785000 ;
      RECT 0.085000  1.785000 0.465000 2.465000 ;
      RECT 0.135000  0.085000 0.465000 0.475000 ;
      RECT 0.685000  0.335000 0.855000 0.655000 ;
      RECT 1.035000  0.085000 1.415000 0.475000 ;
      RECT 1.165000  1.785000 1.335000 2.635000 ;
      RECT 1.505000  1.785000 2.855000 1.955000 ;
      RECT 1.505000  1.955000 1.885000 2.465000 ;
      RECT 2.115000  2.125000 2.285000 2.635000 ;
      RECT 2.455000  1.955000 2.855000 2.465000 ;
      RECT 2.515000  0.825000 2.745000 1.325000 ;
      RECT 3.255000  0.085000 3.545000 0.920000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor2_1


MACRO sky130_fd_sc_hdll__xor2_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.075000 0.925000 1.275000 ;
        RECT 0.755000 1.275000 0.925000 1.445000 ;
        RECT 0.755000 1.445000 2.080000 1.615000 ;
        RECT 1.860000 1.075000 3.530000 1.275000 ;
        RECT 1.860000 1.275000 2.080000 1.445000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.105000 1.075000 1.395000 1.120000 ;
        RECT 1.105000 1.120000 4.055000 1.260000 ;
        RECT 1.105000 1.260000 1.395000 1.305000 ;
        RECT 3.765000 1.075000 4.055000 1.120000 ;
        RECT 3.765000 1.260000 4.055000 1.305000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.806800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.975000 0.645000 4.305000 0.725000 ;
        RECT 3.975000 0.725000 6.350000 0.905000 ;
        RECT 5.385000 0.645000 5.765000 0.725000 ;
        RECT 5.475000 1.415000 6.350000 1.625000 ;
        RECT 5.475000 1.625000 5.725000 2.125000 ;
        RECT 5.985000 0.905000 6.350000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.120000  0.725000 1.850000 0.905000 ;
      RECT 0.120000  0.905000 0.290000 1.785000 ;
      RECT 0.120000  1.785000 2.420000 1.955000 ;
      RECT 0.120000  2.135000 0.400000 2.465000 ;
      RECT 0.145000  2.125000 0.315000 2.135000 ;
      RECT 0.190000  0.085000 0.360000 0.555000 ;
      RECT 0.530000  0.255000 0.910000 0.725000 ;
      RECT 0.620000  2.135000 0.870000 2.635000 ;
      RECT 1.090000  2.135000 1.340000 2.295000 ;
      RECT 1.090000  2.295000 2.280000 2.465000 ;
      RECT 1.130000  0.085000 1.300000 0.555000 ;
      RECT 1.145000  1.075000 1.690000 1.275000 ;
      RECT 1.165000  2.125000 1.335000 2.135000 ;
      RECT 1.470000  0.255000 1.850000 0.725000 ;
      RECT 1.560000  1.955000 1.810000 2.125000 ;
      RECT 2.030000  2.135000 2.280000 2.295000 ;
      RECT 2.070000  0.085000 2.240000 0.555000 ;
      RECT 2.250000  1.445000 5.185000 1.615000 ;
      RECT 2.250000  1.615000 2.420000 1.785000 ;
      RECT 2.485000  2.125000 2.800000 2.465000 ;
      RECT 2.510000  0.255000 2.840000 0.725000 ;
      RECT 2.510000  0.725000 3.700000 0.905000 ;
      RECT 2.590000  1.785000 5.255000 1.955000 ;
      RECT 2.590000  1.955000 2.800000 2.125000 ;
      RECT 3.020000  2.135000 3.270000 2.635000 ;
      RECT 3.060000  0.085000 3.230000 0.555000 ;
      RECT 3.400000  0.255000 4.780000 0.475000 ;
      RECT 3.400000  0.475000 3.700000 0.725000 ;
      RECT 3.490000  1.955000 3.740000 2.465000 ;
      RECT 3.720000  1.075000 4.490000 1.275000 ;
      RECT 3.960000  2.135000 4.265000 2.635000 ;
      RECT 4.485000  1.955000 5.255000 2.295000 ;
      RECT 4.485000  2.295000 6.195000 2.465000 ;
      RECT 5.015000  1.075000 5.725000 1.245000 ;
      RECT 5.015000  1.245000 5.185000 1.445000 ;
      RECT 5.045000  0.085000 5.215000 0.555000 ;
      RECT 5.945000  1.795000 6.195000 2.295000 ;
      RECT 5.985000  0.085000 6.155000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.125000 0.315000 2.295000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.165000  1.105000 1.335000 1.275000 ;
      RECT 1.165000  2.125000 1.335000 2.295000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  1.105000 3.995000 1.275000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.085000 2.095000 0.375000 2.140000 ;
      RECT 0.085000 2.140000 1.395000 2.280000 ;
      RECT 0.085000 2.280000 0.375000 2.325000 ;
      RECT 1.105000 2.095000 1.395000 2.140000 ;
      RECT 1.105000 2.280000 1.395000 2.325000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor2_2


MACRO sky130_fd_sc_hdll__a31oi_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.740000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.225000 0.995000 6.020000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.135000 0.995000 3.950000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.995000 1.885000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.270000 0.995000 7.605000 1.630000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.613500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.425000 0.635000 8.435000 0.805000 ;
        RECT 6.725000 1.915000 8.085000 2.085000 ;
        RECT 7.325000 0.255000 7.495000 0.635000 ;
        RECT 7.845000 0.805000 8.085000 1.915000 ;
        RECT 8.265000 0.255000 8.435000 0.635000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 4.185000 0.805000 ;
      RECT 0.175000  1.495000 6.005000 1.665000 ;
      RECT 0.175000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.895000 0.465000 ;
      RECT 0.515000  1.915000 0.895000 2.635000 ;
      RECT 1.115000  0.255000 1.285000 0.635000 ;
      RECT 1.115000  1.665000 1.285000 2.465000 ;
      RECT 1.455000  0.085000 1.835000 0.465000 ;
      RECT 1.455000  1.915000 1.835000 2.635000 ;
      RECT 2.055000  0.255000 2.225000 0.635000 ;
      RECT 2.055000  1.665000 2.225000 2.465000 ;
      RECT 2.395000  0.295000 6.165000 0.465000 ;
      RECT 2.395000  1.915000 2.775000 2.635000 ;
      RECT 2.995000  1.665000 3.165000 2.465000 ;
      RECT 3.335000  1.915000 3.715000 2.635000 ;
      RECT 3.935000  1.665000 4.105000 2.465000 ;
      RECT 4.295000  1.915000 4.675000 2.635000 ;
      RECT 4.895000  1.665000 5.065000 2.465000 ;
      RECT 5.235000  2.255000 5.615000 2.635000 ;
      RECT 5.835000  1.665000 6.005000 2.255000 ;
      RECT 5.835000  2.255000 8.515000 2.425000 ;
      RECT 5.835000  2.425000 6.005000 2.465000 ;
      RECT 6.725000  0.085000 7.105000 0.465000 ;
      RECT 7.665000  0.085000 8.045000 0.465000 ;
      RECT 8.265000  1.495000 8.515000 2.255000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31oi_4


MACRO sky130_fd_sc_hdll__a31oi_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.760000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.445000 1.695000 1.665000 ;
        RECT 1.370000 0.995000 1.695000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.335000 1.165000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.435000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 0.995000 2.650000 1.325000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.523800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 0.295000 2.155000 0.825000 ;
        RECT 1.985000 0.825000 2.155000 1.495000 ;
        RECT 1.985000 1.495000 2.410000 2.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  0.085000 0.430000 0.815000 ;
      RECT 0.090000  1.495000 0.420000 2.635000 ;
      RECT 0.640000  1.835000 1.815000 2.005000 ;
      RECT 0.640000  2.005000 0.815000 2.415000 ;
      RECT 1.035000  2.175000 1.365000 2.635000 ;
      RECT 1.620000  2.005000 1.815000 2.415000 ;
      RECT 2.325000  0.085000 2.585000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31oi_1


MACRO sky130_fd_sc_hdll__a31oi_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.060000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.330000 0.995000 3.090000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.150000 0.995000 1.905000 1.615000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.995000 0.870000 1.615000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.220000 1.075000 4.940000 1.275000 ;
        RECT 4.715000 1.275000 4.940000 1.625000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.007000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545000 0.655000 4.955000 0.825000 ;
        RECT 3.330000 0.825000 4.955000 0.845000 ;
        RECT 3.330000 0.845000 3.645000 1.445000 ;
        RECT 3.330000 1.445000 4.485000 1.615000 ;
        RECT 3.605000 0.255000 3.775000 0.655000 ;
        RECT 4.155000 1.615000 4.485000 2.115000 ;
        RECT 4.575000 0.295000 4.955000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.095000  0.655000 2.305000 0.825000 ;
      RECT 0.175000  1.785000 3.855000 1.955000 ;
      RECT 0.175000  1.955000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.895000 0.465000 ;
      RECT 0.515000  2.125000 0.895000 2.635000 ;
      RECT 1.115000  1.955000 1.285000 2.465000 ;
      RECT 1.455000  0.295000 3.375000 0.465000 ;
      RECT 1.455000  2.125000 1.835000 2.635000 ;
      RECT 2.055000  1.955000 2.225000 2.465000 ;
      RECT 2.560000  2.125000 3.280000 2.635000 ;
      RECT 3.685000  1.955000 3.855000 2.295000 ;
      RECT 3.685000  2.295000 4.875000 2.465000 ;
      RECT 4.025000  0.085000 4.405000 0.465000 ;
      RECT 4.705000  1.795000 4.875000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31oi_2


MACRO sky130_fd_sc_hdll__dlxtn_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.360000 BY  2.720000 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 0.955000 1.890000 1.325000 ;
    END
  END D
  PIN GATE_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN Q
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.595000 0.415000 5.895000 0.745000 ;
        RECT 5.595000 1.495000 5.895000 2.455000 ;
        RECT 5.710000 0.745000 5.895000 0.995000 ;
        RECT 5.710000 0.995000 7.235000 1.325000 ;
        RECT 5.710000 1.325000 5.895000 1.495000 ;
        RECT 6.535000 0.385000 6.805000 0.995000 ;
        RECT 6.535000 1.325000 6.805000 2.455000 ;
    END
  END Q
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.890000 0.805000 ;
      RECT 0.175000  1.795000 0.890000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.895000 0.465000 ;
      RECT 0.515000  2.135000 0.895000 2.635000 ;
      RECT 0.660000  0.805000 0.890000 1.795000 ;
      RECT 1.115000  0.345000 1.285000 2.465000 ;
      RECT 1.555000  1.495000 2.290000 1.665000 ;
      RECT 1.555000  1.665000 1.885000 2.415000 ;
      RECT 1.635000  0.345000 1.805000 0.615000 ;
      RECT 1.635000  0.615000 2.290000 0.765000 ;
      RECT 1.635000  0.765000 2.540000 0.785000 ;
      RECT 1.975000  0.085000 2.355000 0.445000 ;
      RECT 2.105000  1.835000 2.420000 2.635000 ;
      RECT 2.120000  0.785000 2.540000 1.095000 ;
      RECT 2.120000  1.095000 2.290000 1.495000 ;
      RECT 2.670000  1.355000 2.955000 2.005000 ;
      RECT 2.915000  0.705000 3.345000 1.035000 ;
      RECT 3.025000  2.255000 3.950000 2.425000 ;
      RECT 3.090000  0.365000 3.950000 0.535000 ;
      RECT 3.175000  1.035000 3.345000 1.415000 ;
      RECT 3.175000  1.415000 3.565000 1.995000 ;
      RECT 3.780000  0.535000 3.950000 0.995000 ;
      RECT 3.780000  0.995000 4.500000 1.325000 ;
      RECT 3.780000  1.325000 3.950000 2.255000 ;
      RECT 4.120000  0.085000 4.290000 0.610000 ;
      RECT 4.120000  2.135000 4.290000 2.635000 ;
      RECT 4.140000  1.535000 4.860000 1.865000 ;
      RECT 4.640000  1.865000 4.860000 2.435000 ;
      RECT 4.670000  0.415000 4.860000 0.995000 ;
      RECT 4.670000  0.995000 5.490000 1.325000 ;
      RECT 4.670000  1.325000 4.860000 1.535000 ;
      RECT 5.090000  0.085000 5.375000 0.715000 ;
      RECT 5.090000  1.495000 5.375000 2.635000 ;
      RECT 6.065000  0.085000 6.315000 0.825000 ;
      RECT 6.065000  1.495000 6.315000 2.635000 ;
      RECT 7.005000  0.085000 7.175000 0.715000 ;
      RECT 7.005000  1.495000 7.175000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.660000  1.400000 0.830000 1.570000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.115000  1.770000 1.285000 1.940000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.670000  1.770000 2.840000 1.940000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.175000  1.400000 3.345000 1.570000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 0.600000 1.370000 0.890000 1.460000 ;
      RECT 0.600000 1.460000 3.410000 1.600000 ;
      RECT 1.055000 1.740000 1.345000 1.800000 ;
      RECT 1.055000 1.800000 2.900000 1.940000 ;
      RECT 1.055000 1.940000 1.345000 1.970000 ;
      RECT 2.610000 1.740000 2.900000 1.800000 ;
      RECT 2.610000 1.940000 2.900000 1.970000 ;
      RECT 3.115000 1.370000 3.410000 1.460000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlxtn_4


MACRO sky130_fd_sc_hdll__dlxtn_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.980000 BY  2.720000 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.955000 1.890000 1.325000 ;
    END
  END D
  PIN GATE_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN Q
    ANTENNADIFFAREA  0.554500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.590000 0.415000 5.875000 2.455000 ;
    END
  END Q
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.830000 0.805000 ;
      RECT 0.175000  1.795000 0.830000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.895000 0.465000 ;
      RECT 0.515000  2.135000 0.895000 2.635000 ;
      RECT 0.660000  0.805000 0.830000 1.070000 ;
      RECT 0.660000  1.070000 0.890000 1.400000 ;
      RECT 0.660000  1.400000 0.830000 1.795000 ;
      RECT 1.115000  0.345000 1.285000 1.685000 ;
      RECT 1.115000  1.685000 1.340000 2.465000 ;
      RECT 1.555000  1.495000 2.290000 1.665000 ;
      RECT 1.555000  1.665000 1.885000 2.415000 ;
      RECT 1.635000  0.345000 1.805000 0.615000 ;
      RECT 1.635000  0.615000 2.290000 0.765000 ;
      RECT 1.635000  0.765000 2.540000 0.785000 ;
      RECT 1.975000  0.085000 2.355000 0.445000 ;
      RECT 2.105000  1.835000 2.420000 2.635000 ;
      RECT 2.120000  0.785000 2.540000 1.095000 ;
      RECT 2.120000  1.095000 2.290000 1.495000 ;
      RECT 2.670000  1.355000 2.955000 2.005000 ;
      RECT 2.885000  0.705000 3.340000 1.035000 ;
      RECT 3.005000  0.365000 3.850000 0.535000 ;
      RECT 3.020000  2.255000 3.850000 2.425000 ;
      RECT 3.170000  1.035000 3.340000 1.415000 ;
      RECT 3.170000  1.415000 3.510000 1.995000 ;
      RECT 3.680000  0.535000 3.850000 0.995000 ;
      RECT 3.680000  0.995000 4.430000 1.325000 ;
      RECT 3.680000  1.325000 3.850000 2.255000 ;
      RECT 4.020000  0.085000 4.300000 0.825000 ;
      RECT 4.050000  2.135000 4.350000 2.635000 ;
      RECT 4.070000  1.535000 4.790000 1.865000 ;
      RECT 4.570000  0.415000 4.790000 0.825000 ;
      RECT 4.570000  1.865000 4.790000 2.435000 ;
      RECT 4.620000  0.825000 4.790000 0.995000 ;
      RECT 4.620000  0.995000 5.420000 1.325000 ;
      RECT 4.620000  1.325000 4.790000 1.535000 ;
      RECT 5.020000  0.085000 5.290000 0.825000 ;
      RECT 5.020000  1.495000 5.290000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.660000  1.445000 0.830000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.170000  1.785000 1.340000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.670000  1.785000 2.840000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.175000  1.445000 3.345000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 0.600000 1.415000 0.890000 1.460000 ;
      RECT 0.600000 1.460000 3.405000 1.600000 ;
      RECT 0.600000 1.600000 0.890000 1.645000 ;
      RECT 1.110000 1.755000 1.400000 1.800000 ;
      RECT 1.110000 1.800000 2.900000 1.940000 ;
      RECT 1.110000 1.940000 1.400000 1.985000 ;
      RECT 2.610000 1.755000 2.900000 1.800000 ;
      RECT 2.610000 1.940000 2.900000 1.985000 ;
      RECT 3.115000 1.415000 3.405000 1.460000 ;
      RECT 3.115000 1.600000 3.405000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlxtn_1


MACRO sky130_fd_sc_hdll__dlxtn_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.955000 1.890000 1.325000 ;
    END
  END D
  PIN GATE_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN Q
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.625000 0.415000 5.910000 0.825000 ;
        RECT 5.625000 1.495000 5.910000 2.455000 ;
        RECT 5.740000 0.825000 5.910000 0.995000 ;
        RECT 5.740000 0.995000 6.345000 1.325000 ;
        RECT 5.740000 1.325000 5.910000 1.495000 ;
    END
  END Q
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.830000 0.805000 ;
      RECT 0.175000  1.795000 0.830000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.895000 0.465000 ;
      RECT 0.515000  2.135000 0.895000 2.635000 ;
      RECT 0.660000  0.805000 0.830000 1.070000 ;
      RECT 0.660000  1.070000 0.890000 1.400000 ;
      RECT 0.660000  1.400000 0.830000 1.795000 ;
      RECT 1.115000  0.345000 1.285000 1.685000 ;
      RECT 1.115000  1.685000 1.340000 2.465000 ;
      RECT 1.555000  1.495000 2.290000 1.665000 ;
      RECT 1.555000  1.665000 1.885000 2.415000 ;
      RECT 1.635000  0.345000 1.805000 0.615000 ;
      RECT 1.635000  0.615000 2.290000 0.765000 ;
      RECT 1.635000  0.765000 2.540000 0.785000 ;
      RECT 1.975000  0.085000 2.355000 0.445000 ;
      RECT 2.105000  1.835000 2.420000 2.635000 ;
      RECT 2.120000  0.785000 2.540000 1.095000 ;
      RECT 2.120000  1.095000 2.290000 1.495000 ;
      RECT 2.670000  1.355000 2.955000 2.005000 ;
      RECT 2.915000  0.705000 3.340000 1.035000 ;
      RECT 3.085000  0.365000 3.795000 0.535000 ;
      RECT 3.145000  2.255000 3.945000 2.425000 ;
      RECT 3.170000  1.035000 3.340000 1.415000 ;
      RECT 3.170000  1.415000 3.510000 1.995000 ;
      RECT 3.625000  0.535000 3.795000 0.995000 ;
      RECT 3.625000  0.995000 4.545000 1.165000 ;
      RECT 3.775000  1.165000 4.545000 1.325000 ;
      RECT 3.775000  1.325000 3.945000 2.255000 ;
      RECT 4.035000  0.085000 4.415000 0.825000 ;
      RECT 4.165000  2.135000 4.465000 2.635000 ;
      RECT 4.185000  1.535000 4.905000 1.865000 ;
      RECT 4.685000  0.415000 4.905000 0.825000 ;
      RECT 4.685000  1.865000 4.905000 2.435000 ;
      RECT 4.735000  0.825000 4.905000 0.995000 ;
      RECT 4.735000  0.995000 5.535000 1.325000 ;
      RECT 4.735000  1.325000 4.905000 1.535000 ;
      RECT 5.135000  0.085000 5.405000 0.825000 ;
      RECT 5.135000  1.495000 5.405000 2.635000 ;
      RECT 6.095000  0.085000 6.355000 0.550000 ;
      RECT 6.095000  1.755000 6.345000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.660000  1.445000 0.830000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.170000  1.785000 1.340000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.670000  1.785000 2.840000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.175000  1.445000 3.345000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.600000 1.415000 0.890000 1.460000 ;
      RECT 0.600000 1.460000 3.405000 1.600000 ;
      RECT 0.600000 1.600000 0.890000 1.645000 ;
      RECT 1.110000 1.755000 1.400000 1.800000 ;
      RECT 1.110000 1.800000 2.900000 1.940000 ;
      RECT 1.110000 1.940000 1.400000 1.985000 ;
      RECT 2.610000 1.755000 2.900000 1.800000 ;
      RECT 2.610000 1.940000 2.900000 1.985000 ;
      RECT 3.115000 1.415000 3.405000 1.460000 ;
      RECT 3.115000 1.600000 3.405000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlxtn_2


MACRO sky130_fd_sc_hdll__a21boi_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.360000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.865000 1.065000 5.440000 1.310000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.300000 1.065000 3.695000 1.480000 ;
        RECT 3.300000 1.480000 7.120000 1.705000 ;
        RECT 5.725000 1.075000 7.120000 1.480000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 1.075000 0.670000 1.615000 ;
        RECT 0.450000 0.995000 0.670000 1.075000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.490500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.375000 0.370000 1.565000 0.615000 ;
        RECT 1.375000 0.615000 2.525000 0.695000 ;
        RECT 1.375000 0.695000 5.385000 0.865000 ;
        RECT 1.680000 1.585000 3.130000 1.705000 ;
        RECT 1.680000 1.705000 2.945000 2.035000 ;
        RECT 2.335000 0.255000 2.525000 0.615000 ;
        RECT 2.820000 0.865000 5.385000 0.895000 ;
        RECT 2.820000 0.895000 3.130000 1.585000 ;
        RECT 3.555000 0.675000 5.385000 0.695000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.090000  0.255000 0.445000 0.615000 ;
      RECT 0.090000  0.615000 1.155000 0.795000 ;
      RECT 0.095000  1.785000 1.010000 2.005000 ;
      RECT 0.095000  2.005000 0.425000 2.465000 ;
      RECT 0.645000  2.175000 0.905000 2.635000 ;
      RECT 0.770000  0.085000 1.155000 0.445000 ;
      RECT 0.840000  0.795000 1.155000 1.035000 ;
      RECT 0.840000  1.035000 2.620000 1.345000 ;
      RECT 0.840000  1.345000 1.010000 1.785000 ;
      RECT 1.180000  1.795000 1.425000 2.215000 ;
      RECT 1.180000  2.215000 3.365000 2.465000 ;
      RECT 1.785000  0.085000 2.165000 0.445000 ;
      RECT 2.055000  2.205000 3.365000 2.215000 ;
      RECT 2.745000  0.085000 3.385000 0.525000 ;
      RECT 3.165000  1.875000 7.240000 2.105000 ;
      RECT 3.165000  2.105000 3.365000 2.205000 ;
      RECT 3.535000  2.275000 3.915000 2.635000 ;
      RECT 3.565000  0.255000 5.865000 0.505000 ;
      RECT 4.495000  2.275000 4.875000 2.635000 ;
      RECT 5.095000  2.105000 5.285000 2.465000 ;
      RECT 5.455000  2.275000 5.835000 2.635000 ;
      RECT 5.605000  0.505000 5.865000 0.735000 ;
      RECT 5.605000  0.735000 6.825000 0.905000 ;
      RECT 6.050000  2.105000 6.235000 2.465000 ;
      RECT 6.085000  0.085000 6.275000 0.565000 ;
      RECT 6.415000  2.275000 6.795000 2.635000 ;
      RECT 6.445000  0.255000 6.825000 0.735000 ;
      RECT 6.990000  2.105000 7.240000 2.465000 ;
      RECT 7.000000  0.085000 7.240000 0.885000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21boi_4


MACRO sky130_fd_sc_hdll__a21boi_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855000 0.995000 3.565000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 1.075000 2.675000 1.245000 ;
        RECT 2.300000 1.245000 2.675000 1.495000 ;
        RECT 2.300000 1.495000 4.085000 1.675000 ;
        RECT 3.735000 0.995000 4.085000 1.495000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.765000 0.425000 1.805000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.712500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.255000 1.870000 0.615000 ;
        RECT 1.525000 0.615000 3.360000 0.785000 ;
        RECT 1.525000 0.785000 1.865000 2.115000 ;
        RECT 2.980000 0.255000 3.360000 0.615000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.095000  2.080000 0.425000 2.635000 ;
      RECT 0.265000  0.360000 0.825000 0.530000 ;
      RECT 0.645000  0.530000 0.825000 1.070000 ;
      RECT 0.645000  1.070000 1.355000 1.285000 ;
      RECT 0.645000  1.285000 0.825000 2.265000 ;
      RECT 1.085000  0.085000 1.325000 0.885000 ;
      RECT 1.100000  1.795000 1.350000 2.285000 ;
      RECT 1.100000  2.285000 2.415000 2.465000 ;
      RECT 2.035000  1.855000 4.320000 2.025000 ;
      RECT 2.035000  2.025000 2.415000 2.285000 ;
      RECT 2.140000  0.085000 2.470000 0.445000 ;
      RECT 2.635000  2.195000 2.805000 2.635000 ;
      RECT 3.110000  2.025000 4.320000 2.105000 ;
      RECT 3.110000  2.105000 3.280000 2.465000 ;
      RECT 3.460000  2.275000 3.840000 2.635000 ;
      RECT 3.990000  0.085000 4.330000 0.785000 ;
      RECT 4.060000  2.105000 4.320000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21boi_2


MACRO sky130_fd_sc_hdll__a21boi_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.375000 2.240000 1.345000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.650000 0.995000 3.125000 1.345000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.975000 0.335000 1.665000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.676000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.045000 1.780000 1.345000 ;
        RECT 1.065000 1.345000 1.525000 2.455000 ;
        RECT 1.440000 0.265000 1.780000 1.045000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.095000  1.835000 0.855000 2.005000 ;
      RECT 0.095000  2.005000 0.355000 2.435000 ;
      RECT 0.365000  0.265000 0.855000 0.715000 ;
      RECT 0.515000  0.715000 0.855000 1.835000 ;
      RECT 0.525000  2.175000 0.895000 2.635000 ;
      RECT 1.025000  0.085000 1.255000 0.865000 ;
      RECT 1.745000  1.525000 3.005000 1.725000 ;
      RECT 1.745000  1.725000 1.935000 2.455000 ;
      RECT 2.105000  1.905000 2.485000 2.635000 ;
      RECT 2.715000  0.085000 3.075000 0.815000 ;
      RECT 2.835000  1.725000 3.005000 2.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21boi_1


MACRO sky130_fd_sc_hdll__clkbuf_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  5.520000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.486000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 0.400000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.775400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.570000 0.280000 1.830000 0.735000 ;
        RECT 1.570000 0.735000 5.230000 0.905000 ;
        RECT 1.570000 1.495000 5.230000 1.735000 ;
        RECT 1.570000 1.735000 1.830000 2.460000 ;
        RECT 2.530000 0.280000 2.790000 0.735000 ;
        RECT 2.530000 1.735000 2.790000 2.460000 ;
        RECT 3.490000 0.280000 3.750000 0.735000 ;
        RECT 3.490000 1.735000 3.750000 2.460000 ;
        RECT 4.160000 0.905000 5.230000 1.495000 ;
        RECT 4.450000 0.280000 4.710000 0.735000 ;
        RECT 4.450000 1.735000 4.710000 2.460000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.095000  1.525000 0.390000 2.635000 ;
      RECT 0.145000  0.085000 0.390000 0.545000 ;
      RECT 0.620000  0.265000 0.870000 1.075000 ;
      RECT 0.620000  1.075000 3.990000 1.325000 ;
      RECT 0.620000  1.325000 0.870000 2.460000 ;
      RECT 1.090000  0.085000 1.350000 0.610000 ;
      RECT 1.090000  1.525000 1.350000 2.635000 ;
      RECT 2.050000  0.085000 2.310000 0.565000 ;
      RECT 2.050000  1.905000 2.310000 2.635000 ;
      RECT 3.010000  0.085000 3.270000 0.565000 ;
      RECT 3.010000  1.905000 3.270000 2.635000 ;
      RECT 3.970000  0.085000 4.230000 0.565000 ;
      RECT 3.970000  1.905000 4.230000 2.635000 ;
      RECT 4.930000  0.085000 5.230000 0.565000 ;
      RECT 4.930000  1.905000 5.225000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_8


MACRO sky130_fd_sc_hdll__clkbuf_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  3.220000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.243000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.755000 0.825000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.898200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.345000 1.405000 0.735000 ;
        RECT 1.050000 0.735000 2.910000 0.905000 ;
        RECT 1.145000 1.835000 2.365000 2.005000 ;
        RECT 1.145000 2.005000 1.405000 2.465000 ;
        RECT 2.105000 0.345000 2.365000 0.735000 ;
        RECT 2.105000 1.415000 2.910000 1.650000 ;
        RECT 2.105000 1.650000 2.365000 1.835000 ;
        RECT 2.105000 2.005000 2.365000 2.465000 ;
        RECT 2.410000 0.905000 2.910000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.255000 0.385000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 1.215000 1.665000 ;
      RECT 0.085000  1.665000 0.395000 2.465000 ;
      RECT 0.605000  0.085000 0.880000 0.565000 ;
      RECT 0.615000  1.835000 0.925000 2.635000 ;
      RECT 0.995000  1.075000 2.240000 1.245000 ;
      RECT 0.995000  1.245000 1.215000 1.495000 ;
      RECT 1.625000  0.085000 1.880000 0.565000 ;
      RECT 1.625000  2.175000 1.880000 2.635000 ;
      RECT 2.545000  1.845000 2.875000 2.635000 ;
      RECT 2.585000  0.085000 2.865000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_4


MACRO sky130_fd_sc_hdll__clkbuf_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  2.300000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.243000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.745000 0.835000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.445400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.140000 0.255000 1.345000 0.655000 ;
        RECT 1.140000 0.655000 1.875000 0.825000 ;
        RECT 1.160000 1.855000 1.875000 2.030000 ;
        RECT 1.160000 2.030000 1.345000 2.435000 ;
        RECT 1.485000 0.825000 1.875000 1.855000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 1.315000 1.665000 ;
      RECT 0.085000  1.665000 0.355000 2.435000 ;
      RECT 0.525000  1.855000 0.905000 2.635000 ;
      RECT 0.605000  0.085000 0.880000 0.565000 ;
      RECT 1.015000  0.995000 1.315000 1.495000 ;
      RECT 1.515000  0.085000 1.900000 0.485000 ;
      RECT 1.515000  2.210000 1.900000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_2


MACRO sky130_fd_sc_hdll__clkbuf_6
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.486000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 0.395000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.212300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 0.255000 1.835000 0.735000 ;
        RECT 1.505000 0.735000 4.075000 0.905000 ;
        RECT 1.505000 1.495000 4.075000 1.665000 ;
        RECT 1.505000 1.665000 1.835000 2.460000 ;
        RECT 2.445000 0.255000 2.775000 0.735000 ;
        RECT 2.445000 1.665000 2.775000 2.460000 ;
        RECT 3.385000 0.255000 3.715000 0.735000 ;
        RECT 3.385000 1.665000 3.715000 2.460000 ;
        RECT 3.745000 0.905000 4.075000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.095000  1.495000 0.395000 2.635000 ;
      RECT 0.145000  0.085000 0.395000 0.545000 ;
      RECT 0.565000  0.265000 0.895000 1.075000 ;
      RECT 0.565000  1.075000 3.390000 1.325000 ;
      RECT 0.565000  1.325000 0.895000 2.465000 ;
      RECT 1.065000  0.085000 1.335000 0.610000 ;
      RECT 1.065000  1.495000 1.335000 2.635000 ;
      RECT 2.005000  0.085000 2.275000 0.565000 ;
      RECT 2.005000  1.835000 2.275000 2.635000 ;
      RECT 2.945000  0.085000 3.215000 0.565000 ;
      RECT 2.945000  1.835000 3.215000 2.635000 ;
      RECT 3.885000  0.085000 4.155000 0.565000 ;
      RECT 3.885000  1.835000 4.155000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_6


MACRO sky130_fd_sc_hdll__clkbuf_12
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.280000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.972000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.075000 1.320000 1.305000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.420400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.475000 7.445000 1.665000 ;
        RECT 2.445000 1.665000 2.745000 2.465000 ;
        RECT 2.475000 0.280000 2.745000 0.715000 ;
        RECT 2.475000 0.715000 7.445000 0.905000 ;
        RECT 3.415000 0.280000 3.685000 0.715000 ;
        RECT 3.415000 1.665000 3.685000 2.465000 ;
        RECT 4.355000 0.280000 4.625000 0.715000 ;
        RECT 4.355000 1.665000 4.625000 2.465000 ;
        RECT 5.295000 0.280000 5.565000 0.715000 ;
        RECT 5.295000 1.665000 5.565000 2.465000 ;
        RECT 6.235000 0.280000 6.505000 0.715000 ;
        RECT 6.235000 1.665000 6.505000 2.465000 ;
        RECT 6.960000 0.905000 7.445000 1.475000 ;
        RECT 7.175000 0.280000 7.445000 0.715000 ;
        RECT 7.175000 1.665000 7.445000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.610000 ;
      RECT 0.095000  1.495000 0.395000 2.635000 ;
      RECT 0.565000  1.495000 1.805000 1.665000 ;
      RECT 0.565000  1.665000 0.895000 2.465000 ;
      RECT 0.570000  1.475000 1.805000 1.495000 ;
      RECT 0.595000  0.280000 0.865000 0.715000 ;
      RECT 0.595000  0.715000 1.805000 0.905000 ;
      RECT 1.035000  0.085000 1.365000 0.545000 ;
      RECT 1.065000  1.835000 1.335000 2.635000 ;
      RECT 1.535000  0.280000 1.805000 0.715000 ;
      RECT 1.535000  0.905000 1.805000 1.075000 ;
      RECT 1.535000  1.075000 6.685000 1.305000 ;
      RECT 1.535000  1.305000 1.805000 1.475000 ;
      RECT 1.535000  1.665000 1.805000 2.465000 ;
      RECT 1.975000  0.085000 2.305000 0.545000 ;
      RECT 1.975000  1.475000 2.275000 2.635000 ;
      RECT 2.915000  0.085000 3.245000 0.545000 ;
      RECT 2.915000  1.835000 3.245000 2.635000 ;
      RECT 3.855000  0.085000 4.185000 0.545000 ;
      RECT 3.855000  1.835000 4.185000 2.635000 ;
      RECT 4.795000  0.085000 5.125000 0.545000 ;
      RECT 4.795000  1.835000 5.125000 2.635000 ;
      RECT 5.735000  0.085000 6.065000 0.545000 ;
      RECT 5.735000  1.835000 6.065000 2.635000 ;
      RECT 6.675000  0.085000 7.005000 0.545000 ;
      RECT 6.675000  1.835000 7.005000 2.635000 ;
      RECT 7.615000  0.085000 7.945000 0.610000 ;
      RECT 7.615000  1.465000 7.945000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_12


MACRO sky130_fd_sc_hdll__clkbuf_16
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.12000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.972000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.400000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.529800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.530000 0.280000  2.790000 0.735000 ;
        RECT 2.530000 0.735000 10.025000 0.905000 ;
        RECT 2.530000 1.495000 10.025000 1.720000 ;
        RECT 2.530000 1.720000  8.535000 1.735000 ;
        RECT 2.530000 1.735000  2.790000 2.460000 ;
        RECT 3.490000 0.280000  3.750000 0.735000 ;
        RECT 3.490000 1.735000  3.750000 2.460000 ;
        RECT 4.450000 0.280000  4.710000 0.735000 ;
        RECT 4.450000 1.735000  4.710000 2.460000 ;
        RECT 5.345000 0.280000  5.670000 0.735000 ;
        RECT 5.410000 1.735000  5.670000 2.460000 ;
        RECT 6.355000 0.280000  6.615000 0.735000 ;
        RECT 6.355000 1.735000  6.615000 2.460000 ;
        RECT 7.315000 0.280000  7.575000 0.735000 ;
        RECT 7.315000 1.735000  7.575000 2.460000 ;
        RECT 8.275000 0.280000  8.535000 0.735000 ;
        RECT 8.275000 1.735000  8.535000 2.460000 ;
        RECT 8.760000 0.905000 10.025000 1.495000 ;
        RECT 9.245000 0.280000  9.505000 0.735000 ;
        RECT 9.245000 1.720000  9.535000 2.460000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.085000  0.390000 0.595000 ;
      RECT 0.095000  1.825000  0.390000 2.635000 ;
      RECT 0.620000  0.265000  0.870000 1.075000 ;
      RECT 0.620000  1.075000  8.540000 1.325000 ;
      RECT 0.620000  1.325000  0.865000 2.465000 ;
      RECT 1.090000  0.085000  1.350000 0.610000 ;
      RECT 1.090000  1.825000  1.350000 2.635000 ;
      RECT 1.580000  0.265000  1.830000 1.075000 ;
      RECT 1.580000  1.325000  1.830000 2.460000 ;
      RECT 2.050000  0.085000  2.310000 0.645000 ;
      RECT 2.050000  1.835000  2.310000 2.630000 ;
      RECT 2.050000  2.630000  9.025000 2.635000 ;
      RECT 3.010000  0.085000  3.270000 0.565000 ;
      RECT 3.010000  1.905000  3.270000 2.630000 ;
      RECT 3.970000  0.085000  4.230000 0.565000 ;
      RECT 3.970000  1.905000  4.230000 2.630000 ;
      RECT 4.930000  0.085000  5.175000 0.565000 ;
      RECT 4.930000  1.905000  5.190000 2.630000 ;
      RECT 5.890000  0.085000  6.135000 0.565000 ;
      RECT 5.890000  1.905000  6.135000 2.630000 ;
      RECT 6.845000  0.085000  7.095000 0.565000 ;
      RECT 6.850000  1.905000  7.095000 2.630000 ;
      RECT 7.805000  0.085000  8.055000 0.565000 ;
      RECT 7.810000  1.905000  8.055000 2.630000 ;
      RECT 8.765000  0.085000  9.025000 0.565000 ;
      RECT 8.770000  1.905000  9.025000 2.630000 ;
      RECT 9.725000  0.085000 10.025000 0.565000 ;
      RECT 9.755000  1.890000 10.025000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_16


MACRO sky130_fd_sc_hdll__clkbuf_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  1.840000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.220200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.365000 0.985000 1.745000 1.355000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.374500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.345000 0.760000 ;
        RECT 0.085000 0.760000 0.255000 1.560000 ;
        RECT 0.085000 1.560000 0.355000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.425000  1.060000 0.760000 1.390000 ;
      RECT 0.525000  0.085000 1.275000 0.465000 ;
      RECT 0.525000  1.875000 1.275000 2.635000 ;
      RECT 0.540000  0.635000 1.625000 0.805000 ;
      RECT 0.540000  0.805000 0.760000 1.060000 ;
      RECT 0.540000  1.390000 0.760000 1.535000 ;
      RECT 0.540000  1.535000 1.665000 1.705000 ;
      RECT 1.455000  0.255000 1.625000 0.635000 ;
      RECT 1.495000  1.705000 1.665000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkbuf_1


MACRO sky130_fd_sc_hdll__sdfxtp_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.96000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.745000 1.355000 3.150000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.030000 0.305000 10.410000 0.735000 ;
        RECT 10.030000 0.735000 11.850000 0.905000 ;
        RECT 10.030000 1.505000 11.850000 1.675000 ;
        RECT 10.030000 1.675000 10.410000 2.395000 ;
        RECT 10.980000 0.305000 11.360000 0.735000 ;
        RECT 10.980000 1.675000 11.360000 2.395000 ;
        RECT 11.550000 0.905000 11.850000 1.505000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.035000 4.095000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.880000 0.615000 3.505000 0.785000 ;
        RECT 1.880000 0.785000 2.215000 1.685000 ;
        RECT 3.335000 0.785000 3.505000 1.115000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.895000 0.805000 ;
      RECT  0.180000  1.795000  0.895000 1.965000 ;
      RECT  0.180000  1.965000  0.350000 2.465000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.520000  2.135000  0.900000 2.635000 ;
      RECT  0.665000  0.805000  0.895000 1.795000 ;
      RECT  1.115000  0.345000  1.345000 2.465000 ;
      RECT  1.535000  0.275000  1.905000 0.445000 ;
      RECT  1.535000  0.445000  1.705000 1.860000 ;
      RECT  1.535000  1.860000  3.525000 2.075000 ;
      RECT  1.535000  2.075000  1.810000 2.445000 ;
      RECT  1.980000  2.245000  2.360000 2.635000 ;
      RECT  2.125000  0.085000  2.455000 0.445000 ;
      RECT  2.385000  0.955000  2.715000 1.125000 ;
      RECT  2.385000  1.125000  2.555000 1.860000 ;
      RECT  2.895000  2.245000  3.890000 2.415000 ;
      RECT  3.070000  0.275000  3.895000 0.445000 ;
      RECT  3.330000  1.355000  3.525000 1.860000 ;
      RECT  3.720000  1.825000  4.735000 1.995000 ;
      RECT  3.720000  1.995000  3.890000 2.245000 ;
      RECT  3.725000  0.445000  3.895000 0.695000 ;
      RECT  3.725000  0.695000  4.735000 0.865000 ;
      RECT  4.110000  2.165000  4.280000 2.635000 ;
      RECT  4.115000  0.085000  4.315000 0.525000 ;
      RECT  4.565000  0.365000  4.915000 0.535000 ;
      RECT  4.565000  0.535000  4.735000 0.695000 ;
      RECT  4.565000  0.865000  4.735000 1.825000 ;
      RECT  4.565000  1.995000  4.735000 2.065000 ;
      RECT  4.565000  2.065000  4.800000 2.440000 ;
      RECT  4.905000  0.705000  5.535000 1.035000 ;
      RECT  4.905000  1.035000  5.195000 1.905000 ;
      RECT  5.045000  2.190000  6.265000 2.360000 ;
      RECT  5.135000  0.365000  5.895000 0.535000 ;
      RECT  5.385000  1.655000  5.875000 2.010000 ;
      RECT  5.725000  0.535000  5.895000 1.245000 ;
      RECT  5.725000  1.245000  6.605000 1.485000 ;
      RECT  6.045000  1.485000  6.605000 1.575000 ;
      RECT  6.045000  1.575000  6.265000 2.190000 ;
      RECT  6.065000  0.765000  6.995000 1.065000 ;
      RECT  6.225000  0.085000  6.595000 0.585000 ;
      RECT  6.435000  1.835000  6.605000 2.635000 ;
      RECT  6.775000  0.365000  7.285000 0.535000 ;
      RECT  6.775000  0.535000  6.995000 0.765000 ;
      RECT  6.775000  1.065000  6.995000 2.135000 ;
      RECT  6.775000  2.135000  7.075000 2.465000 ;
      RECT  7.165000  0.705000  7.765000 1.035000 ;
      RECT  7.165000  1.245000  7.405000 1.965000 ;
      RECT  7.300000  2.165000  8.335000 2.335000 ;
      RECT  7.565000  0.365000  8.205000 0.535000 ;
      RECT  7.575000  1.035000  7.765000 1.575000 ;
      RECT  7.575000  1.575000  7.945000 1.905000 ;
      RECT  7.985000  0.535000  8.205000 0.995000 ;
      RECT  7.985000  0.995000  9.150000 1.325000 ;
      RECT  7.985000  1.325000  8.335000 1.405000 ;
      RECT  8.165000  1.405000  8.335000 2.165000 ;
      RECT  8.450000  0.085000  8.870000 0.615000 ;
      RECT  8.555000  1.575000  9.505000 1.905000 ;
      RECT  8.565000  2.135000  8.870000 2.635000 ;
      RECT  9.140000  0.300000  9.500000 0.825000 ;
      RECT  9.220000  1.905000  9.505000 2.455000 ;
      RECT  9.320000  0.825000  9.500000 1.075000 ;
      RECT  9.320000  1.075000 11.380000 1.325000 ;
      RECT  9.320000  1.325000  9.505000 1.575000 ;
      RECT  9.690000  0.085000  9.860000 0.695000 ;
      RECT  9.690000  1.625000  9.860000 2.635000 ;
      RECT 10.640000  0.085000 10.810000 0.565000 ;
      RECT 10.640000  1.845000 10.810000 2.635000 ;
      RECT 11.580000  0.085000 11.750000 0.565000 ;
      RECT 11.580000  1.845000 11.750000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.665000  1.740000  0.835000 1.910000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.155000  0.720000  1.325000 0.890000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.155000  0.720000  5.325000 0.890000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  1.740000  5.835000 1.910000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.225000  0.720000  7.395000 0.890000 ;
      RECT  7.225000  1.740000  7.395000 1.910000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.605000 1.710000 0.895000 1.800000 ;
      RECT 0.605000 1.800000 7.455000 1.940000 ;
      RECT 1.095000 0.690000 1.385000 0.780000 ;
      RECT 1.095000 0.780000 7.455000 0.920000 ;
      RECT 5.045000 0.690000 5.385000 0.780000 ;
      RECT 5.555000 1.710000 5.895000 1.800000 ;
      RECT 7.115000 0.690000 7.455000 0.780000 ;
      RECT 7.115000 1.710000 7.455000 1.800000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfxtp_4


MACRO sky130_fd_sc_hdll__sdfxtp_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  11.04000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.745000 1.355000 3.150000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.030000 0.305000 10.500000 0.820000 ;
        RECT 10.030000 1.545000 10.500000 2.395000 ;
        RECT 10.330000 0.820000 10.500000 1.545000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.035000 4.095000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.880000 0.615000 3.505000 0.785000 ;
        RECT 1.880000 0.785000 2.215000 1.685000 ;
        RECT 3.335000 0.785000 3.505000 1.115000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.895000 0.805000 ;
      RECT  0.180000  1.795000  0.895000 1.965000 ;
      RECT  0.180000  1.965000  0.350000 2.465000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.520000  2.135000  0.900000 2.635000 ;
      RECT  0.665000  0.805000  0.895000 1.795000 ;
      RECT  1.115000  0.345000  1.345000 2.465000 ;
      RECT  1.535000  0.275000  1.905000 0.445000 ;
      RECT  1.535000  0.445000  1.705000 1.860000 ;
      RECT  1.535000  1.860000  3.525000 2.075000 ;
      RECT  1.535000  2.075000  1.810000 2.445000 ;
      RECT  1.980000  2.245000  2.360000 2.635000 ;
      RECT  2.125000  0.085000  2.455000 0.445000 ;
      RECT  2.385000  0.955000  2.715000 1.125000 ;
      RECT  2.385000  1.125000  2.555000 1.860000 ;
      RECT  2.895000  2.245000  3.890000 2.415000 ;
      RECT  3.070000  0.275000  3.895000 0.445000 ;
      RECT  3.330000  1.355000  3.525000 1.860000 ;
      RECT  3.720000  1.825000  4.735000 1.995000 ;
      RECT  3.720000  1.995000  3.890000 2.245000 ;
      RECT  3.725000  0.445000  3.895000 0.695000 ;
      RECT  3.725000  0.695000  4.735000 0.865000 ;
      RECT  4.110000  2.165000  4.280000 2.635000 ;
      RECT  4.115000  0.085000  4.315000 0.525000 ;
      RECT  4.565000  0.365000  4.915000 0.535000 ;
      RECT  4.565000  0.535000  4.735000 0.695000 ;
      RECT  4.565000  0.865000  4.735000 1.825000 ;
      RECT  4.565000  1.995000  4.735000 2.065000 ;
      RECT  4.565000  2.065000  4.800000 2.440000 ;
      RECT  4.905000  0.705000  5.535000 1.035000 ;
      RECT  4.905000  1.035000  5.195000 1.905000 ;
      RECT  5.045000  2.190000  6.265000 2.360000 ;
      RECT  5.135000  0.365000  5.895000 0.535000 ;
      RECT  5.385000  1.655000  5.875000 2.010000 ;
      RECT  5.725000  0.535000  5.895000 1.245000 ;
      RECT  5.725000  1.245000  6.605000 1.485000 ;
      RECT  6.045000  1.485000  6.605000 1.575000 ;
      RECT  6.045000  1.575000  6.265000 2.190000 ;
      RECT  6.065000  0.765000  6.995000 1.065000 ;
      RECT  6.225000  0.085000  6.595000 0.585000 ;
      RECT  6.435000  1.835000  6.605000 2.635000 ;
      RECT  6.775000  0.365000  7.285000 0.535000 ;
      RECT  6.775000  0.535000  6.995000 0.765000 ;
      RECT  6.775000  1.065000  6.995000 2.135000 ;
      RECT  6.775000  2.135000  7.075000 2.465000 ;
      RECT  7.165000  0.705000  7.765000 1.035000 ;
      RECT  7.165000  1.245000  7.405000 1.965000 ;
      RECT  7.300000  2.165000  8.335000 2.335000 ;
      RECT  7.565000  0.365000  8.205000 0.535000 ;
      RECT  7.575000  1.035000  7.765000 1.575000 ;
      RECT  7.575000  1.575000  7.945000 1.905000 ;
      RECT  7.985000  0.535000  8.205000 0.995000 ;
      RECT  7.985000  0.995000  9.150000 1.325000 ;
      RECT  7.985000  1.325000  8.335000 1.405000 ;
      RECT  8.165000  1.405000  8.335000 2.165000 ;
      RECT  8.450000  0.085000  8.870000 0.615000 ;
      RECT  8.555000  1.575000  9.505000 1.905000 ;
      RECT  8.565000  2.135000  8.870000 2.635000 ;
      RECT  9.140000  0.300000  9.500000 0.825000 ;
      RECT  9.220000  1.905000  9.505000 2.455000 ;
      RECT  9.320000  0.825000  9.500000 0.995000 ;
      RECT  9.320000  0.995000 10.130000 1.325000 ;
      RECT  9.320000  1.325000  9.505000 1.575000 ;
      RECT  9.690000  0.085000  9.860000 0.695000 ;
      RECT  9.690000  1.625000  9.860000 2.635000 ;
      RECT 10.670000  0.085000 10.840000 0.565000 ;
      RECT 10.670000  1.845000 10.840000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.665000  1.740000  0.835000 1.910000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.155000  0.720000  1.325000 0.890000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.155000  0.720000  5.325000 0.890000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  1.740000  5.835000 1.910000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.225000  0.720000  7.395000 0.890000 ;
      RECT  7.225000  1.740000  7.395000 1.910000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.605000 1.710000 0.895000 1.800000 ;
      RECT 0.605000 1.800000 7.455000 1.940000 ;
      RECT 1.095000 0.690000 1.385000 0.780000 ;
      RECT 1.095000 0.780000 7.455000 0.920000 ;
      RECT 5.045000 0.690000 5.385000 0.780000 ;
      RECT 5.555000 1.710000 5.895000 1.800000 ;
      RECT 7.115000 0.690000 7.455000 0.780000 ;
      RECT 7.115000 1.710000 7.455000 1.800000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfxtp_2


MACRO sky130_fd_sc_hdll__sdfxtp_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.58000 BY  2.720000 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.745000 1.355000 3.150000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.471500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.930000 0.305000 10.470000 0.820000 ;
        RECT  9.930000 1.545000 10.470000 2.395000 ;
        RECT 10.230000 0.820000 10.470000 1.545000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.035000 4.095000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.880000 0.615000 3.505000 0.785000 ;
        RECT 1.880000 0.785000 2.215000 1.685000 ;
        RECT 3.335000 0.785000 3.505000 1.115000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.580000 0.085000 ;
      RECT 0.000000  2.635000 10.580000 2.805000 ;
      RECT 0.175000  0.345000  0.345000 0.635000 ;
      RECT 0.175000  0.635000  0.895000 0.805000 ;
      RECT 0.180000  1.795000  0.895000 1.965000 ;
      RECT 0.180000  1.965000  0.350000 2.465000 ;
      RECT 0.515000  0.085000  0.895000 0.465000 ;
      RECT 0.520000  2.135000  0.900000 2.635000 ;
      RECT 0.665000  0.805000  0.895000 1.795000 ;
      RECT 1.115000  0.345000  1.345000 2.465000 ;
      RECT 1.535000  0.275000  1.905000 0.445000 ;
      RECT 1.535000  0.445000  1.705000 1.860000 ;
      RECT 1.535000  1.860000  3.540000 2.075000 ;
      RECT 1.535000  2.075000  1.810000 2.445000 ;
      RECT 1.980000  2.245000  2.360000 2.635000 ;
      RECT 2.075000  0.085000  2.405000 0.445000 ;
      RECT 2.385000  0.955000  2.715000 1.125000 ;
      RECT 2.385000  1.125000  2.555000 1.860000 ;
      RECT 2.895000  2.245000  3.890000 2.415000 ;
      RECT 3.070000  0.275000  3.895000 0.445000 ;
      RECT 3.330000  1.355000  3.540000 1.860000 ;
      RECT 3.720000  1.825000  4.735000 1.995000 ;
      RECT 3.720000  1.995000  3.890000 2.245000 ;
      RECT 3.725000  0.445000  3.895000 0.695000 ;
      RECT 3.725000  0.695000  4.735000 0.865000 ;
      RECT 4.110000  2.165000  4.280000 2.635000 ;
      RECT 4.115000  0.085000  4.315000 0.525000 ;
      RECT 4.565000  0.365000  4.915000 0.535000 ;
      RECT 4.565000  0.535000  4.735000 0.695000 ;
      RECT 4.565000  0.865000  4.735000 1.825000 ;
      RECT 4.565000  1.995000  4.735000 2.065000 ;
      RECT 4.565000  2.065000  4.800000 2.440000 ;
      RECT 4.905000  0.705000  5.535000 1.035000 ;
      RECT 4.905000  1.035000  5.195000 1.905000 ;
      RECT 5.045000  2.190000  6.230000 2.360000 ;
      RECT 5.135000  0.365000  5.875000 0.535000 ;
      RECT 5.385000  1.655000  5.875000 2.010000 ;
      RECT 5.705000  0.535000  5.875000 1.315000 ;
      RECT 5.705000  1.315000  6.685000 1.485000 ;
      RECT 6.045000  0.765000  7.060000 1.095000 ;
      RECT 6.045000  1.485000  6.685000 1.575000 ;
      RECT 6.045000  1.575000  6.230000 2.190000 ;
      RECT 6.225000  0.085000  6.595000 0.585000 ;
      RECT 6.400000  1.835000  6.570000 2.635000 ;
      RECT 6.775000  0.365000  7.260000 0.535000 ;
      RECT 6.775000  0.535000  7.060000 0.765000 ;
      RECT 6.855000  1.095000  7.060000 2.465000 ;
      RECT 7.230000  1.245000  7.470000 1.965000 ;
      RECT 7.250000  0.705000  7.945000 1.035000 ;
      RECT 7.250000  2.165000  8.285000 2.335000 ;
      RECT 7.455000  0.365000  8.285000 0.535000 ;
      RECT 7.735000  1.035000  7.945000 1.905000 ;
      RECT 8.115000  0.535000  8.285000 0.995000 ;
      RECT 8.115000  0.995000  9.050000 1.325000 ;
      RECT 8.115000  1.325000  8.285000 2.165000 ;
      RECT 8.455000  0.085000  8.770000 0.615000 ;
      RECT 8.455000  1.575000  9.405000 1.905000 ;
      RECT 8.465000  2.135000  8.770000 2.635000 ;
      RECT 9.040000  0.300000  9.400000 0.825000 ;
      RECT 9.120000  1.905000  9.405000 2.455000 ;
      RECT 9.220000  0.825000  9.400000 0.995000 ;
      RECT 9.220000  0.995000 10.030000 1.325000 ;
      RECT 9.220000  1.325000  9.405000 1.575000 ;
      RECT 9.590000  0.085000  9.760000 0.695000 ;
      RECT 9.590000  1.625000  9.760000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.665000  1.740000  0.835000 1.910000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.155000  0.720000  1.325000 0.890000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.155000  0.720000  5.325000 0.890000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  1.740000  5.835000 1.910000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.240000  1.740000  7.410000 1.910000 ;
      RECT  7.310000  0.720000  7.480000 0.890000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 0.605000 1.710000 0.895000 1.800000 ;
      RECT 0.605000 1.800000 7.470000 1.940000 ;
      RECT 1.095000 0.690000 1.385000 0.780000 ;
      RECT 1.095000 0.780000 7.540000 0.920000 ;
      RECT 5.045000 0.690000 5.385000 0.780000 ;
      RECT 5.555000 1.710000 5.895000 1.800000 ;
      RECT 7.130000 1.710000 7.470000 1.800000 ;
      RECT 7.230000 0.690000 7.540000 0.780000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfxtp_1


END LIBRARY
